* NGSPICE file created from opamp133.ext - technology: sky130A

.subckt opamp133 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 CSoutput.t173 a_n8964_8799.t40 vdd.t300 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X1 a_n2472_13878.t27 a_n2650_13878.t43 a_n2650_13878.t44 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 a_n2472_13878.t7 a_n2650_13878.t60 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t299 a_n8964_8799.t41 CSoutput.t172 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 a_n8964_8799.t26 plus.t5 a_n3827_n3924.t39 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X5 CSoutput.t171 a_n8964_8799.t42 vdd.t298 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 gnd.t173 commonsourceibias.t64 CSoutput.t47 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 a_n3827_n3924.t17 diffpairibias.t20 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X8 a_n3827_n3924.t38 plus.t6 a_n8964_8799.t36 gnd.t300 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X9 CSoutput.t170 a_n8964_8799.t43 vdd.t297 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X10 commonsourceibias.t63 commonsourceibias.t62 gnd.t110 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 gnd.t293 gnd.t291 gnd.t292 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X12 vdd.t296 a_n8964_8799.t44 CSoutput.t169 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 vdd.t134 CSoutput.t184 output.t17 gnd.t158 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X14 a_n2650_8322.t27 a_n2650_13878.t61 a_n8964_8799.t21 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 gnd.t290 gnd.t288 gnd.t289 gnd.t202 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X16 CSoutput.t48 commonsourceibias.t65 gnd.t174 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 CSoutput.t168 a_n8964_8799.t45 vdd.t295 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 vdd.t294 a_n8964_8799.t46 CSoutput.t167 vdd.t280 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X19 CSoutput.t166 a_n8964_8799.t47 vdd.t293 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 gnd.t24 commonsourceibias.t60 commonsourceibias.t61 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t33 commonsourceibias.t66 gnd.t108 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 vdd.t292 a_n8964_8799.t48 CSoutput.t165 vdd.t280 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 vdd.t291 a_n8964_8799.t49 CSoutput.t164 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 gnd.t287 gnd.t285 gnd.t286 gnd.t202 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X25 commonsourceibias.t59 commonsourceibias.t58 gnd.t77 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 a_n2650_13878.t49 minus.t5 a_n3827_n3924.t16 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 a_n8964_8799.t12 plus.t7 a_n3827_n3924.t37 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 a_n8964_8799.t28 a_n2650_13878.t62 a_n2650_8322.t26 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 CSoutput.t22 commonsourceibias.t67 gnd.t75 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 a_n2650_13878.t0 minus.t6 a_n3827_n3924.t0 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X31 vdd.t290 a_n8964_8799.t50 CSoutput.t163 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 vdd.t289 a_n8964_8799.t51 CSoutput.t162 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 a_n8964_8799.t29 a_n2650_13878.t63 a_n2650_8322.t25 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X34 commonsourceibias.t57 commonsourceibias.t56 gnd.t79 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t284 gnd.t282 gnd.t283 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X36 CSoutput.t185 a_n2650_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X37 CSoutput.t161 a_n8964_8799.t52 vdd.t288 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X38 a_n3827_n3924.t36 plus.t8 a_n8964_8799.t6 gnd.t299 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X39 CSoutput.t46 commonsourceibias.t68 gnd.t172 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 a_n3827_n3924.t9 diffpairibias.t21 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X41 a_n3827_n3924.t4 minus.t7 a_n2650_13878.t4 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X42 CSoutput.t160 a_n8964_8799.t53 vdd.t287 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 gnd.t281 gnd.t278 gnd.t280 gnd.t279 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X44 gnd.t43 commonsourceibias.t69 CSoutput.t11 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 vdd.t284 a_n8964_8799.t54 CSoutput.t159 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 gnd.t111 commonsourceibias.t54 commonsourceibias.t55 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X47 output.t16 CSoutput.t186 vdd.t12 gnd.t157 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X48 CSoutput.t158 a_n8964_8799.t55 vdd.t286 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 commonsourceibias.t53 commonsourceibias.t52 gnd.t175 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 vdd.t285 a_n8964_8799.t56 CSoutput.t157 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X51 vdd.t96 vdd.t94 vdd.t95 vdd.t30 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X52 gnd.t74 commonsourceibias.t70 CSoutput.t21 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 a_n2472_13878.t26 a_n2650_13878.t27 a_n2650_13878.t28 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X54 a_n2650_13878.t10 a_n2650_13878.t9 a_n2472_13878.t25 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X55 CSoutput.t187 a_n2650_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X56 gnd.t171 commonsourceibias.t71 CSoutput.t45 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 CSoutput.t156 a_n8964_8799.t57 vdd.t283 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 output.t15 CSoutput.t188 vdd.t13 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X59 vdd.t93 vdd.t91 vdd.t92 vdd.t68 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X60 a_n3827_n3924.t35 plus.t9 a_n8964_8799.t32 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X61 vdd.t282 a_n8964_8799.t58 CSoutput.t155 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 vdd.t281 a_n8964_8799.t59 CSoutput.t154 vdd.t280 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 gnd.t176 commonsourceibias.t50 commonsourceibias.t51 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 plus.t2 gnd.t275 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X65 diffpairibias.t19 diffpairibias.t18 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X66 a_n3827_n3924.t34 plus.t10 a_n8964_8799.t39 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X67 gnd.t274 gnd.t272 gnd.t273 gnd.t248 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X68 commonsourceibias.t49 commonsourceibias.t48 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 a_n2650_13878.t42 a_n2650_13878.t41 a_n2472_13878.t24 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X70 CSoutput.t153 a_n8964_8799.t60 vdd.t279 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 vdd.t278 a_n8964_8799.t61 CSoutput.t152 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 a_n8964_8799.t24 a_n2650_13878.t64 a_n2650_8322.t24 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X73 CSoutput.t151 a_n8964_8799.t62 vdd.t277 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 commonsourceibias.t47 commonsourceibias.t46 gnd.t112 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 a_n2650_13878.t12 a_n2650_13878.t11 a_n2472_13878.t23 vdd.t117 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X76 vdd.t276 a_n8964_8799.t63 CSoutput.t150 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 vdd.t275 a_n8964_8799.t64 CSoutput.t149 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 a_n8964_8799.t25 a_n2650_13878.t65 a_n2650_8322.t23 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X79 gnd.t271 gnd.t269 gnd.t270 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X80 diffpairibias.t17 diffpairibias.t16 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X81 gnd.t177 commonsourceibias.t44 commonsourceibias.t45 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 CSoutput.t148 a_n8964_8799.t65 vdd.t274 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 CSoutput.t44 commonsourceibias.t72 gnd.t170 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 output.t19 outputibias.t8 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X85 a_n2650_8322.t22 a_n2650_13878.t66 a_n8964_8799.t16 vdd.t117 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X86 CSoutput.t147 a_n8964_8799.t66 vdd.t273 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 vdd.t16 CSoutput.t189 output.t14 gnd.t155 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X88 a_n3827_n3924.t11 minus.t8 a_n2650_13878.t7 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X89 vdd.t17 CSoutput.t190 output.t13 gnd.t154 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X90 gnd.t113 commonsourceibias.t42 commonsourceibias.t43 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 CSoutput.t32 commonsourceibias.t73 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 a_n3827_n3924.t33 plus.t11 a_n8964_8799.t20 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X93 CSoutput.t20 commonsourceibias.t74 gnd.t72 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 gnd.t268 gnd.t266 gnd.t267 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X95 a_n8964_8799.t33 plus.t12 a_n3827_n3924.t32 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X96 gnd.t265 gnd.t263 minus.t4 gnd.t264 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X97 CSoutput.t31 commonsourceibias.t75 gnd.t105 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X98 outputibias.t7 outputibias.t6 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X99 CSoutput.t19 commonsourceibias.t76 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 vdd.t90 vdd.t88 vdd.t89 vdd.t64 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X101 a_n3827_n3924.t8 diffpairibias.t22 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X102 vdd.t272 a_n8964_8799.t67 CSoutput.t146 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 vdd.t271 a_n8964_8799.t68 CSoutput.t145 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 a_n2650_13878.t14 a_n2650_13878.t13 a_n2472_13878.t22 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X105 vdd.t270 a_n8964_8799.t69 CSoutput.t144 vdd.t200 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X106 a_n3827_n3924.t31 plus.t13 a_n8964_8799.t19 gnd.t297 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X107 vdd.t269 a_n8964_8799.t70 CSoutput.t143 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 a_n8964_8799.t17 a_n2650_13878.t67 a_n2650_8322.t21 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X109 a_n2650_13878.t30 a_n2650_13878.t29 a_n2472_13878.t21 vdd.t0 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X110 gnd.t304 commonsourceibias.t40 commonsourceibias.t41 gnd.t303 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 gnd.t32 commonsourceibias.t38 commonsourceibias.t39 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 vdd.t268 a_n8964_8799.t71 CSoutput.t142 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 CSoutput.t141 a_n8964_8799.t72 vdd.t267 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 CSoutput.t140 a_n8964_8799.t73 vdd.t266 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 diffpairibias.t15 diffpairibias.t14 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X116 vdd.t87 vdd.t85 vdd.t86 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X117 CSoutput.t139 a_n8964_8799.t74 vdd.t265 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X118 gnd.t169 commonsourceibias.t77 CSoutput.t43 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 vdd.t84 vdd.t81 vdd.t83 vdd.t82 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 gnd.t42 commonsourceibias.t78 CSoutput.t10 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X121 gnd.t66 commonsourceibias.t79 CSoutput.t18 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 gnd.t184 commonsourceibias.t80 CSoutput.t51 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 CSoutput.t138 a_n8964_8799.t75 vdd.t264 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 output.t12 CSoutput.t191 vdd.t18 gnd.t153 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X125 vdd.t263 a_n8964_8799.t76 CSoutput.t137 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 vdd.t98 CSoutput.t192 output.t11 gnd.t152 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X127 vdd.t138 a_n2650_13878.t68 a_n2650_8322.t7 vdd.t137 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 a_n2650_13878.t46 a_n2650_13878.t45 a_n2472_13878.t20 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 gnd.t65 commonsourceibias.t81 CSoutput.t17 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X130 vdd.t80 vdd.t78 vdd.t79 vdd.t48 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X131 gnd.t262 gnd.t260 gnd.t261 gnd.t221 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X132 a_n2650_8322.t6 a_n2650_13878.t69 vdd.t140 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X133 a_n3827_n3924.t12 diffpairibias.t23 gnd.t98 gnd.t97 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X134 CSoutput.t136 a_n8964_8799.t77 vdd.t262 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X135 vdd.t108 a_n2650_13878.t70 a_n2472_13878.t6 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 vdd.t77 vdd.t75 vdd.t76 vdd.t64 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X137 gnd.t141 commonsourceibias.t82 CSoutput.t42 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 vdd.t74 vdd.t71 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 vdd.t261 a_n8964_8799.t78 CSoutput.t135 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X140 plus.t0 gnd.t257 gnd.t259 gnd.t258 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X141 vdd.t259 a_n8964_8799.t79 CSoutput.t134 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 gnd.t256 gnd.t254 minus.t3 gnd.t255 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X143 a_n8964_8799.t9 plus.t14 a_n3827_n3924.t30 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X144 a_n2650_13878.t54 minus.t9 a_n3827_n3924.t43 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X145 vdd.t70 vdd.t67 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X146 a_n2650_8322.t5 a_n2650_13878.t71 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X147 a_n8964_8799.t7 a_n2650_13878.t72 a_n2650_8322.t20 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X148 a_n8964_8799.t30 plus.t15 a_n3827_n3924.t29 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X149 CSoutput.t133 a_n8964_8799.t80 vdd.t258 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 diffpairibias.t13 diffpairibias.t12 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X151 vdd.t257 a_n8964_8799.t81 CSoutput.t132 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X152 a_n2650_13878.t24 a_n2650_13878.t23 a_n2472_13878.t19 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 vdd.t255 a_n8964_8799.t82 CSoutput.t131 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 a_n8964_8799.t8 a_n2650_13878.t73 a_n2650_8322.t19 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 CSoutput.t130 a_n8964_8799.t83 vdd.t254 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 CSoutput.t129 a_n8964_8799.t84 vdd.t252 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 CSoutput.t128 a_n8964_8799.t85 vdd.t251 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 CSoutput.t50 commonsourceibias.t83 gnd.t183 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 a_n2472_13878.t18 a_n2650_13878.t35 a_n2650_13878.t36 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 commonsourceibias.t37 commonsourceibias.t36 gnd.t124 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 CSoutput.t16 commonsourceibias.t84 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 CSoutput.t41 commonsourceibias.t85 gnd.t140 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X163 vdd.t99 CSoutput.t193 output.t10 gnd.t151 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X164 vdd.t66 vdd.t63 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X165 vdd.t62 vdd.t60 vdd.t61 vdd.t34 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X166 CSoutput.t49 commonsourceibias.t86 gnd.t182 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 gnd.t315 commonsourceibias.t87 CSoutput.t181 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 gnd.t253 gnd.t251 minus.t2 gnd.t252 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X169 CSoutput.t127 a_n8964_8799.t86 vdd.t250 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 gnd.t122 commonsourceibias.t34 commonsourceibias.t35 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 vdd.t303 a_n2650_13878.t74 a_n2650_8322.t4 vdd.t302 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X172 a_n2472_13878.t17 a_n2650_13878.t21 a_n2650_13878.t22 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X173 vdd.t249 a_n8964_8799.t87 CSoutput.t126 vdd.t236 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X174 vdd.t248 a_n8964_8799.t88 CSoutput.t125 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 a_n2650_13878.t57 minus.t10 a_n3827_n3924.t46 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X176 a_n3827_n3924.t28 plus.t16 a_n8964_8799.t3 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X177 vdd.t59 vdd.t57 vdd.t58 vdd.t48 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X178 a_n2650_13878.t16 a_n2650_13878.t15 a_n2472_13878.t16 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X179 commonsourceibias.t33 commonsourceibias.t32 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 gnd.t83 commonsourceibias.t30 commonsourceibias.t31 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 vdd.t247 a_n8964_8799.t89 CSoutput.t124 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 gnd.t84 commonsourceibias.t28 commonsourceibias.t29 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 a_n3827_n3924.t48 diffpairibias.t24 gnd.t322 gnd.t321 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X184 commonsourceibias.t27 commonsourceibias.t26 gnd.t114 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 a_n3827_n3924.t42 diffpairibias.t25 gnd.t307 gnd.t306 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 outputibias.t5 outputibias.t4 gnd.t327 gnd.t326 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X187 gnd.t30 commonsourceibias.t88 CSoutput.t6 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 a_n8964_8799.t37 plus.t17 a_n3827_n3924.t27 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X189 vdd.t246 a_n8964_8799.t90 CSoutput.t123 vdd.t236 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X190 vdd.t245 a_n8964_8799.t91 CSoutput.t122 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 gnd.t7 commonsourceibias.t89 CSoutput.t1 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 CSoutput.t121 a_n8964_8799.t92 vdd.t244 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X193 gnd.t53 commonsourceibias.t90 CSoutput.t15 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 gnd.t319 commonsourceibias.t91 CSoutput.t183 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X195 a_n8964_8799.t23 plus.t18 a_n3827_n3924.t26 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X196 gnd.t23 commonsourceibias.t92 CSoutput.t4 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X197 a_n2472_13878.t15 a_n2650_13878.t17 a_n2650_13878.t18 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X198 vdd.t56 vdd.t54 vdd.t55 vdd.t26 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X199 a_n2650_8322.t18 a_n2650_13878.t75 a_n8964_8799.t38 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X200 CSoutput.t120 a_n8964_8799.t93 vdd.t242 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X201 CSoutput.t119 a_n8964_8799.t94 vdd.t243 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 commonsourceibias.t25 commonsourceibias.t24 gnd.t178 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 CSoutput.t118 a_n8964_8799.t95 vdd.t241 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X204 outputibias.t3 outputibias.t2 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X205 gnd.t132 commonsourceibias.t93 CSoutput.t36 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 CSoutput.t24 commonsourceibias.t94 gnd.t90 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 diffpairibias.t11 diffpairibias.t10 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X208 a_n2472_13878.t5 a_n2650_13878.t76 vdd.t4 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 a_n2650_13878.t6 minus.t11 a_n3827_n3924.t6 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X210 gnd.t305 commonsourceibias.t95 CSoutput.t53 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 vdd.t6 a_n2650_13878.t77 a_n2472_13878.t4 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X212 gnd.t179 commonsourceibias.t22 commonsourceibias.t23 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 CSoutput.t117 a_n8964_8799.t96 vdd.t239 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X214 a_n3827_n3924.t25 plus.t19 a_n8964_8799.t14 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X215 vdd.t237 a_n8964_8799.t97 CSoutput.t116 vdd.t236 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X216 vdd.t235 a_n8964_8799.t98 CSoutput.t115 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 commonsourceibias.t21 commonsourceibias.t20 gnd.t127 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 vdd.t233 a_n8964_8799.t99 CSoutput.t114 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 CSoutput.t40 commonsourceibias.t96 gnd.t139 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 CSoutput.t113 a_n8964_8799.t100 vdd.t231 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 a_n2472_13878.t14 a_n2650_13878.t31 a_n2650_13878.t32 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X222 diffpairibias.t9 diffpairibias.t8 gnd.t324 gnd.t323 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X223 vdd.t230 a_n8964_8799.t101 CSoutput.t112 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 gnd.t126 commonsourceibias.t18 commonsourceibias.t19 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 CSoutput.t2 commonsourceibias.t97 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X226 a_n3827_n3924.t19 minus.t12 a_n2650_13878.t51 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X227 a_n2650_8322.t17 a_n2650_13878.t78 a_n8964_8799.t27 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X228 CSoutput.t111 a_n8964_8799.t102 vdd.t229 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 diffpairibias.t7 diffpairibias.t6 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X230 vdd.t228 a_n8964_8799.t103 CSoutput.t110 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 a_n2472_13878.t13 a_n2650_13878.t19 a_n2650_13878.t20 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X232 vdd.t129 a_n2650_13878.t79 a_n2650_8322.t3 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X233 vdd.t226 a_n8964_8799.t104 CSoutput.t109 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 a_n3827_n3924.t18 minus.t13 a_n2650_13878.t50 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X235 gnd.t250 gnd.t247 gnd.t249 gnd.t248 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X236 vdd.t100 CSoutput.t194 output.t9 gnd.t150 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X237 CSoutput.t195 a_n2650_8322.t31 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X238 CSoutput.t39 commonsourceibias.t98 gnd.t138 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 CSoutput.t5 commonsourceibias.t99 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 gnd.t5 commonsourceibias.t100 CSoutput.t0 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 gnd.t246 gnd.t244 plus.t3 gnd.t245 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X242 a_n3827_n3924.t44 minus.t14 a_n2650_13878.t55 gnd.t300 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X243 minus.t1 gnd.t237 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X244 CSoutput.t108 a_n8964_8799.t105 vdd.t224 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 gnd.t243 gnd.t240 gnd.t242 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X246 a_n2472_13878.t3 a_n2650_13878.t80 vdd.t102 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X247 outputibias.t1 outputibias.t0 gnd.t317 gnd.t316 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X248 vdd.t53 vdd.t51 vdd.t52 vdd.t34 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X249 CSoutput.t52 commonsourceibias.t101 gnd.t302 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 commonsourceibias.t17 commonsourceibias.t16 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X251 vdd.t223 a_n8964_8799.t106 CSoutput.t107 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 vdd.t221 a_n8964_8799.t107 CSoutput.t106 vdd.t200 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X253 CSoutput.t105 a_n8964_8799.t108 vdd.t220 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 CSoutput.t196 a_n2650_8322.t30 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X255 CSoutput.t104 a_n8964_8799.t109 vdd.t218 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 gnd.t236 gnd.t234 gnd.t235 gnd.t221 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X257 gnd.t233 gnd.t230 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X258 vdd.t217 a_n8964_8799.t110 CSoutput.t103 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X259 a_n3827_n3924.t7 diffpairibias.t26 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X260 vdd.t104 a_n2650_13878.t81 a_n2650_8322.t2 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X261 a_n2650_8322.t16 a_n2650_13878.t82 a_n8964_8799.t4 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X262 a_n8964_8799.t18 plus.t20 a_n3827_n3924.t24 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X263 gnd.t104 commonsourceibias.t102 CSoutput.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 a_n2650_13878.t1 minus.t15 a_n3827_n3924.t1 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X265 CSoutput.t102 a_n8964_8799.t111 vdd.t216 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 vdd.t50 vdd.t47 vdd.t49 vdd.t48 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X267 vdd.t215 a_n8964_8799.t112 CSoutput.t101 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 a_n3827_n3924.t13 minus.t16 a_n2650_13878.t8 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X269 vdd.t46 vdd.t44 vdd.t45 vdd.t22 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X270 vdd.t214 a_n8964_8799.t113 CSoutput.t100 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 vdd.t213 a_n8964_8799.t114 CSoutput.t99 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 output.t0 outputibias.t9 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X273 gnd.t318 commonsourceibias.t103 CSoutput.t182 gnd.t303 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 CSoutput.t3 commonsourceibias.t104 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 vdd.t43 vdd.t40 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X276 a_n3827_n3924.t45 minus.t17 a_n2650_13878.t56 gnd.t297 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X277 vdd.t212 a_n8964_8799.t115 CSoutput.t98 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X278 CSoutput.t97 a_n8964_8799.t116 vdd.t211 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 a_n3827_n3924.t47 minus.t18 a_n2650_13878.t58 gnd.t299 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X280 gnd.t131 commonsourceibias.t105 CSoutput.t35 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 a_n2472_13878.t12 a_n2650_13878.t33 a_n2650_13878.t34 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X282 CSoutput.t96 a_n8964_8799.t117 vdd.t209 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 CSoutput.t95 a_n8964_8799.t118 vdd.t208 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 CSoutput.t23 commonsourceibias.t106 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 a_n2650_8322.t15 a_n2650_13878.t83 a_n8964_8799.t5 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X286 vdd.t39 vdd.t37 vdd.t38 vdd.t22 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X287 diffpairibias.t5 diffpairibias.t4 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X288 commonsourceibias.t15 commonsourceibias.t14 gnd.t115 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X289 gnd.t103 commonsourceibias.t107 CSoutput.t29 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 gnd.t229 gnd.t227 gnd.t228 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X291 CSoutput.t38 commonsourceibias.t108 gnd.t137 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 gnd.t116 commonsourceibias.t12 commonsourceibias.t13 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 CSoutput.t94 a_n8964_8799.t119 vdd.t207 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 CSoutput.t93 a_n8964_8799.t120 vdd.t205 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 CSoutput.t92 a_n8964_8799.t121 vdd.t203 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 a_n3827_n3924.t15 diffpairibias.t27 gnd.t129 gnd.t128 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X297 vdd.t202 a_n8964_8799.t122 CSoutput.t91 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 vdd.t36 vdd.t33 vdd.t35 vdd.t34 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X299 CSoutput.t37 commonsourceibias.t109 gnd.t136 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 vdd.t201 a_n8964_8799.t123 CSoutput.t90 vdd.t200 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X301 gnd.t226 gnd.t224 plus.t1 gnd.t225 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X302 a_n2650_8322.t1 a_n2650_13878.t84 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X303 CSoutput.t89 a_n8964_8799.t124 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 CSoutput.t28 commonsourceibias.t110 gnd.t102 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X305 a_n3827_n3924.t5 minus.t19 a_n2650_13878.t5 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X306 vdd.t197 a_n8964_8799.t125 CSoutput.t88 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X307 CSoutput.t87 a_n8964_8799.t126 vdd.t196 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 vdd.t121 a_n2650_13878.t85 a_n2472_13878.t2 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X309 gnd.t134 commonsourceibias.t10 commonsourceibias.t11 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 vdd.t195 a_n8964_8799.t127 CSoutput.t86 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 CSoutput.t85 a_n8964_8799.t128 vdd.t193 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 output.t8 CSoutput.t197 vdd.t301 gnd.t149 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X313 CSoutput.t27 commonsourceibias.t111 gnd.t101 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 CSoutput.t84 a_n8964_8799.t129 vdd.t191 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 gnd.t100 commonsourceibias.t112 CSoutput.t26 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 vdd.t190 a_n8964_8799.t130 CSoutput.t83 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 vdd.t188 a_n8964_8799.t131 CSoutput.t82 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 vdd.t186 a_n8964_8799.t132 CSoutput.t81 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 CSoutput.t25 commonsourceibias.t113 gnd.t99 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 commonsourceibias.t9 commonsourceibias.t8 gnd.t325 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X321 a_n2650_8322.t14 a_n2650_13878.t86 a_n8964_8799.t1 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X322 CSoutput.t180 commonsourceibias.t114 gnd.t314 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 a_n8964_8799.t2 a_n2650_13878.t87 a_n2650_8322.t13 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X324 output.t7 CSoutput.t198 vdd.t115 gnd.t148 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X325 gnd.t320 commonsourceibias.t6 commonsourceibias.t7 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 a_n2472_13878.t1 a_n2650_13878.t88 vdd.t126 vdd.t125 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X327 gnd.t313 commonsourceibias.t115 CSoutput.t179 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 vdd.t32 vdd.t29 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X329 vdd.t185 a_n8964_8799.t133 CSoutput.t80 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 vdd.t28 vdd.t25 vdd.t27 vdd.t26 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X331 CSoutput.t79 a_n8964_8799.t134 vdd.t184 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 CSoutput.t78 a_n8964_8799.t135 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 CSoutput.t77 a_n8964_8799.t136 vdd.t180 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X334 gnd.t223 gnd.t220 gnd.t222 gnd.t221 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X335 gnd.t219 gnd.t217 plus.t4 gnd.t218 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X336 vdd.t24 vdd.t21 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X337 a_n3827_n3924.t23 plus.t21 a_n8964_8799.t15 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X338 minus.t0 gnd.t190 gnd.t192 gnd.t191 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X339 commonsourceibias.t5 commonsourceibias.t4 gnd.t67 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 a_n2650_13878.t53 minus.t20 a_n3827_n3924.t41 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X341 a_n8964_8799.t22 a_n2650_13878.t89 a_n2650_8322.t12 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X342 a_n2650_8322.t11 a_n2650_13878.t90 a_n8964_8799.t34 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X343 CSoutput.t199 a_n2650_8322.t29 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X344 gnd.t216 gnd.t213 gnd.t215 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X345 a_n2650_13878.t59 minus.t21 a_n3827_n3924.t49 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X346 vdd.t179 a_n8964_8799.t137 CSoutput.t76 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 CSoutput.t75 a_n8964_8799.t138 vdd.t177 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 CSoutput.t74 a_n8964_8799.t139 vdd.t175 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 gnd.t185 commonsourceibias.t2 commonsourceibias.t3 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 CSoutput.t73 a_n8964_8799.t140 vdd.t174 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 a_n2472_13878.t11 a_n2650_13878.t37 a_n2650_13878.t38 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X352 vdd.t173 a_n8964_8799.t141 CSoutput.t72 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 gnd.t312 commonsourceibias.t116 CSoutput.t178 gnd.t303 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 CSoutput.t174 commonsourceibias.t117 gnd.t308 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 output.t6 CSoutput.t200 vdd.t116 gnd.t147 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X356 gnd.t311 commonsourceibias.t118 CSoutput.t177 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 a_n3827_n3924.t40 minus.t22 a_n2650_13878.t52 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X358 a_n3827_n3924.t10 diffpairibias.t28 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X359 vdd.t172 a_n8964_8799.t142 CSoutput.t71 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X360 gnd.t212 gnd.t209 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X361 CSoutput.t70 a_n8964_8799.t143 vdd.t171 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X362 gnd.t208 gnd.t205 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X363 a_n2650_13878.t40 a_n2650_13878.t39 a_n2472_13878.t10 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X364 gnd.t204 gnd.t201 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X365 a_n8964_8799.t35 a_n2650_13878.t91 a_n2650_8322.t10 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X366 output.t18 outputibias.t10 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X367 vdd.t170 a_n8964_8799.t144 CSoutput.t69 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 gnd.t310 commonsourceibias.t119 CSoutput.t176 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 CSoutput.t68 a_n8964_8799.t145 vdd.t169 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X370 vdd.t112 CSoutput.t201 output.t5 gnd.t146 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X371 gnd.t200 gnd.t197 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X372 CSoutput.t34 commonsourceibias.t120 gnd.t125 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 CSoutput.t175 commonsourceibias.t121 gnd.t309 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 diffpairibias.t3 diffpairibias.t2 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X375 vdd.t167 a_n8964_8799.t146 CSoutput.t67 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t66 a_n8964_8799.t147 vdd.t165 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X377 output.t1 outputibias.t11 gnd.t119 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X378 CSoutput.t65 a_n8964_8799.t148 vdd.t164 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X379 a_n2650_8322.t9 a_n2650_13878.t92 a_n8964_8799.t31 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X380 a_n2650_13878.t3 minus.t23 a_n3827_n3924.t3 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X381 vdd.t162 a_n8964_8799.t149 CSoutput.t64 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 CSoutput.t63 a_n8964_8799.t150 vdd.t160 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X383 CSoutput.t62 a_n8964_8799.t151 vdd.t158 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 diffpairibias.t1 diffpairibias.t0 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X385 CSoutput.t14 commonsourceibias.t122 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X386 CSoutput.t202 a_n2650_8322.t28 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X387 vdd.t133 a_n2650_13878.t93 a_n2472_13878.t0 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X388 gnd.t40 commonsourceibias.t123 CSoutput.t9 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 CSoutput.t61 a_n8964_8799.t152 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X390 gnd.t196 gnd.t193 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X391 gnd.t189 gnd.t186 gnd.t188 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X392 vdd.t113 CSoutput.t203 output.t4 gnd.t145 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X393 vdd.t154 a_n8964_8799.t153 CSoutput.t60 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X394 vdd.t152 a_n8964_8799.t154 CSoutput.t59 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X395 CSoutput.t13 commonsourceibias.t124 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 CSoutput.t58 a_n8964_8799.t155 vdd.t150 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 output.t3 CSoutput.t204 vdd.t135 gnd.t144 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X398 gnd.t38 commonsourceibias.t125 CSoutput.t8 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 a_n8964_8799.t13 plus.t22 a_n3827_n3924.t22 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X400 a_n2650_13878.t2 minus.t24 a_n3827_n3924.t2 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X401 gnd.t47 commonsourceibias.t126 CSoutput.t12 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 a_n8964_8799.t10 plus.t23 a_n3827_n3924.t21 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X403 a_n2650_8322.t8 a_n2650_13878.t94 a_n8964_8799.t0 vdd.t0 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X404 vdd.t148 a_n8964_8799.t156 CSoutput.t57 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 vdd.t146 a_n8964_8799.t157 CSoutput.t56 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X406 CSoutput.t55 a_n8964_8799.t158 vdd.t144 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X407 output.t2 CSoutput.t205 vdd.t136 gnd.t143 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X408 gnd.t36 commonsourceibias.t127 CSoutput.t7 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 a_n2650_8322.t0 a_n2650_13878.t95 vdd.t2 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X410 a_n2472_13878.t9 a_n2650_13878.t25 a_n2650_13878.t26 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X411 commonsourceibias.t1 commonsourceibias.t0 gnd.t142 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X412 a_n3827_n3924.t20 plus.t24 a_n8964_8799.t11 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X413 a_n3827_n3924.t14 diffpairibias.t29 gnd.t121 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X414 CSoutput.t54 a_n8964_8799.t159 vdd.t142 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 a_n2650_13878.t48 a_n2650_13878.t47 a_n2472_13878.t8 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 a_n8964_8799.n226 a_n8964_8799.t136 485.149
R1 a_n8964_8799.n245 a_n8964_8799.t150 485.149
R2 a_n8964_8799.n265 a_n8964_8799.t92 485.149
R3 a_n8964_8799.n165 a_n8964_8799.t87 485.149
R4 a_n8964_8799.n184 a_n8964_8799.t97 485.149
R5 a_n8964_8799.n204 a_n8964_8799.t90 485.149
R6 a_n8964_8799.n56 a_n8964_8799.t107 485.135
R7 a_n8964_8799.n238 a_n8964_8799.t43 464.166
R8 a_n8964_8799.n220 a_n8964_8799.t113 464.166
R9 a_n8964_8799.n237 a_n8964_8799.t111 464.166
R10 a_n8964_8799.n236 a_n8964_8799.t49 464.166
R11 a_n8964_8799.n221 a_n8964_8799.t47 464.166
R12 a_n8964_8799.n235 a_n8964_8799.t133 464.166
R13 a_n8964_8799.n234 a_n8964_8799.t65 464.166
R14 a_n8964_8799.n222 a_n8964_8799.t51 464.166
R15 a_n8964_8799.n233 a_n8964_8799.t139 464.166
R16 a_n8964_8799.n232 a_n8964_8799.t91 464.166
R17 a_n8964_8799.n223 a_n8964_8799.t66 464.166
R18 a_n8964_8799.n231 a_n8964_8799.t157 464.166
R19 a_n8964_8799.n230 a_n8964_8799.t109 464.166
R20 a_n8964_8799.n224 a_n8964_8799.t68 464.166
R21 a_n8964_8799.n229 a_n8964_8799.t151 464.166
R22 a_n8964_8799.n228 a_n8964_8799.t112 464.166
R23 a_n8964_8799.n225 a_n8964_8799.t85 464.166
R24 a_n8964_8799.n227 a_n8964_8799.t48 464.166
R25 a_n8964_8799.n71 a_n8964_8799.t123 485.135
R26 a_n8964_8799.n257 a_n8964_8799.t55 464.166
R27 a_n8964_8799.n239 a_n8964_8799.t131 464.166
R28 a_n8964_8799.n256 a_n8964_8799.t129 464.166
R29 a_n8964_8799.n255 a_n8964_8799.t58 464.166
R30 a_n8964_8799.n240 a_n8964_8799.t57 464.166
R31 a_n8964_8799.n254 a_n8964_8799.t149 464.166
R32 a_n8964_8799.n253 a_n8964_8799.t74 464.166
R33 a_n8964_8799.n241 a_n8964_8799.t64 464.166
R34 a_n8964_8799.n252 a_n8964_8799.t152 464.166
R35 a_n8964_8799.n251 a_n8964_8799.t104 464.166
R36 a_n8964_8799.n242 a_n8964_8799.t77 464.166
R37 a_n8964_8799.n250 a_n8964_8799.t50 464.166
R38 a_n8964_8799.n249 a_n8964_8799.t124 464.166
R39 a_n8964_8799.n243 a_n8964_8799.t78 464.166
R40 a_n8964_8799.n248 a_n8964_8799.t42 464.166
R41 a_n8964_8799.n247 a_n8964_8799.t130 464.166
R42 a_n8964_8799.n244 a_n8964_8799.t93 464.166
R43 a_n8964_8799.n246 a_n8964_8799.t59 464.166
R44 a_n8964_8799.n86 a_n8964_8799.t69 485.135
R45 a_n8964_8799.n277 a_n8964_8799.t155 464.166
R46 a_n8964_8799.n259 a_n8964_8799.t122 464.166
R47 a_n8964_8799.n276 a_n8964_8799.t148 464.166
R48 a_n8964_8799.n275 a_n8964_8799.t103 464.166
R49 a_n8964_8799.n260 a_n8964_8799.t128 464.166
R50 a_n8964_8799.n274 a_n8964_8799.t63 464.166
R51 a_n8964_8799.n273 a_n8964_8799.t145 464.166
R52 a_n8964_8799.n261 a_n8964_8799.t81 464.166
R53 a_n8964_8799.n272 a_n8964_8799.t140 464.166
R54 a_n8964_8799.n271 a_n8964_8799.t67 464.166
R55 a_n8964_8799.n262 a_n8964_8799.t116 464.166
R56 a_n8964_8799.n270 a_n8964_8799.t54 464.166
R57 a_n8964_8799.n269 a_n8964_8799.t100 464.166
R58 a_n8964_8799.n263 a_n8964_8799.t76 464.166
R59 a_n8964_8799.n268 a_n8964_8799.t126 464.166
R60 a_n8964_8799.n267 a_n8964_8799.t61 464.166
R61 a_n8964_8799.n264 a_n8964_8799.t108 464.166
R62 a_n8964_8799.n266 a_n8964_8799.t46 464.166
R63 a_n8964_8799.n166 a_n8964_8799.t117 464.166
R64 a_n8964_8799.n167 a_n8964_8799.t44 464.166
R65 a_n8964_8799.n168 a_n8964_8799.t72 464.166
R66 a_n8964_8799.n169 a_n8964_8799.t110 464.166
R67 a_n8964_8799.n164 a_n8964_8799.t147 464.166
R68 a_n8964_8799.n170 a_n8964_8799.t70 464.166
R69 a_n8964_8799.n171 a_n8964_8799.t105 464.166
R70 a_n8964_8799.n172 a_n8964_8799.t142 464.166
R71 a_n8964_8799.n173 a_n8964_8799.t143 464.166
R72 a_n8964_8799.n163 a_n8964_8799.t89 464.166
R73 a_n8964_8799.n174 a_n8964_8799.t121 464.166
R74 a_n8964_8799.n162 a_n8964_8799.t141 464.166
R75 a_n8964_8799.n175 a_n8964_8799.t86 464.166
R76 a_n8964_8799.n176 a_n8964_8799.t88 464.166
R77 a_n8964_8799.n177 a_n8964_8799.t118 464.166
R78 a_n8964_8799.n178 a_n8964_8799.t71 464.166
R79 a_n8964_8799.n161 a_n8964_8799.t73 464.166
R80 a_n8964_8799.n179 a_n8964_8799.t114 464.166
R81 a_n8964_8799.n185 a_n8964_8799.t134 464.166
R82 a_n8964_8799.n186 a_n8964_8799.t56 464.166
R83 a_n8964_8799.n187 a_n8964_8799.t83 464.166
R84 a_n8964_8799.n188 a_n8964_8799.t125 464.166
R85 a_n8964_8799.n183 a_n8964_8799.t159 464.166
R86 a_n8964_8799.n189 a_n8964_8799.t79 464.166
R87 a_n8964_8799.n190 a_n8964_8799.t119 464.166
R88 a_n8964_8799.n191 a_n8964_8799.t156 464.166
R89 a_n8964_8799.n192 a_n8964_8799.t158 464.166
R90 a_n8964_8799.n182 a_n8964_8799.t101 464.166
R91 a_n8964_8799.n193 a_n8964_8799.t138 464.166
R92 a_n8964_8799.n181 a_n8964_8799.t154 464.166
R93 a_n8964_8799.n194 a_n8964_8799.t96 464.166
R94 a_n8964_8799.n195 a_n8964_8799.t98 464.166
R95 a_n8964_8799.n196 a_n8964_8799.t135 464.166
R96 a_n8964_8799.n197 a_n8964_8799.t82 464.166
R97 a_n8964_8799.n180 a_n8964_8799.t84 464.166
R98 a_n8964_8799.n198 a_n8964_8799.t132 464.166
R99 a_n8964_8799.n205 a_n8964_8799.t45 464.166
R100 a_n8964_8799.n206 a_n8964_8799.t106 464.166
R101 a_n8964_8799.n207 a_n8964_8799.t60 464.166
R102 a_n8964_8799.n208 a_n8964_8799.t127 464.166
R103 a_n8964_8799.n203 a_n8964_8799.t75 464.166
R104 a_n8964_8799.n209 a_n8964_8799.t99 464.166
R105 a_n8964_8799.n210 a_n8964_8799.t53 464.166
R106 a_n8964_8799.n211 a_n8964_8799.t115 464.166
R107 a_n8964_8799.n212 a_n8964_8799.t94 464.166
R108 a_n8964_8799.n202 a_n8964_8799.t137 464.166
R109 a_n8964_8799.n213 a_n8964_8799.t80 464.166
R110 a_n8964_8799.n201 a_n8964_8799.t144 464.166
R111 a_n8964_8799.n214 a_n8964_8799.t62 464.166
R112 a_n8964_8799.n215 a_n8964_8799.t41 464.166
R113 a_n8964_8799.n216 a_n8964_8799.t102 464.166
R114 a_n8964_8799.n217 a_n8964_8799.t146 464.166
R115 a_n8964_8799.n200 a_n8964_8799.t120 464.166
R116 a_n8964_8799.n218 a_n8964_8799.t153 464.166
R117 a_n8964_8799.n45 a_n8964_8799.n70 71.7212
R118 a_n8964_8799.n70 a_n8964_8799.n225 17.8606
R119 a_n8964_8799.n69 a_n8964_8799.n45 76.9909
R120 a_n8964_8799.n228 a_n8964_8799.n69 7.32118
R121 a_n8964_8799.n68 a_n8964_8799.n44 78.3454
R122 a_n8964_8799.n44 a_n8964_8799.n67 72.8951
R123 a_n8964_8799.n66 a_n8964_8799.n46 70.1674
R124 a_n8964_8799.n231 a_n8964_8799.n66 20.9683
R125 a_n8964_8799.n46 a_n8964_8799.n65 72.3034
R126 a_n8964_8799.n65 a_n8964_8799.n223 16.6962
R127 a_n8964_8799.n64 a_n8964_8799.n47 77.6622
R128 a_n8964_8799.n232 a_n8964_8799.n64 5.97853
R129 a_n8964_8799.n63 a_n8964_8799.n47 77.6622
R130 a_n8964_8799.n48 a_n8964_8799.n62 72.3034
R131 a_n8964_8799.n61 a_n8964_8799.n48 70.1674
R132 a_n8964_8799.n235 a_n8964_8799.n61 20.9683
R133 a_n8964_8799.n50 a_n8964_8799.n60 72.8951
R134 a_n8964_8799.n60 a_n8964_8799.n221 15.5127
R135 a_n8964_8799.n59 a_n8964_8799.n50 78.3454
R136 a_n8964_8799.n236 a_n8964_8799.n59 4.61226
R137 a_n8964_8799.n58 a_n8964_8799.n49 76.9909
R138 a_n8964_8799.n49 a_n8964_8799.n57 71.7212
R139 a_n8964_8799.n238 a_n8964_8799.n56 20.9683
R140 a_n8964_8799.n51 a_n8964_8799.n56 70.1674
R141 a_n8964_8799.n37 a_n8964_8799.n85 71.7212
R142 a_n8964_8799.n85 a_n8964_8799.n244 17.8606
R143 a_n8964_8799.n84 a_n8964_8799.n37 76.9909
R144 a_n8964_8799.n247 a_n8964_8799.n84 7.32118
R145 a_n8964_8799.n83 a_n8964_8799.n36 78.3454
R146 a_n8964_8799.n36 a_n8964_8799.n82 72.8951
R147 a_n8964_8799.n81 a_n8964_8799.n38 70.1674
R148 a_n8964_8799.n250 a_n8964_8799.n81 20.9683
R149 a_n8964_8799.n38 a_n8964_8799.n80 72.3034
R150 a_n8964_8799.n80 a_n8964_8799.n242 16.6962
R151 a_n8964_8799.n79 a_n8964_8799.n39 77.6622
R152 a_n8964_8799.n251 a_n8964_8799.n79 5.97853
R153 a_n8964_8799.n78 a_n8964_8799.n39 77.6622
R154 a_n8964_8799.n40 a_n8964_8799.n77 72.3034
R155 a_n8964_8799.n76 a_n8964_8799.n40 70.1674
R156 a_n8964_8799.n254 a_n8964_8799.n76 20.9683
R157 a_n8964_8799.n42 a_n8964_8799.n75 72.8951
R158 a_n8964_8799.n75 a_n8964_8799.n240 15.5127
R159 a_n8964_8799.n74 a_n8964_8799.n42 78.3454
R160 a_n8964_8799.n255 a_n8964_8799.n74 4.61226
R161 a_n8964_8799.n73 a_n8964_8799.n41 76.9909
R162 a_n8964_8799.n41 a_n8964_8799.n72 71.7212
R163 a_n8964_8799.n257 a_n8964_8799.n71 20.9683
R164 a_n8964_8799.n43 a_n8964_8799.n71 70.1674
R165 a_n8964_8799.n29 a_n8964_8799.n100 71.7212
R166 a_n8964_8799.n100 a_n8964_8799.n264 17.8606
R167 a_n8964_8799.n99 a_n8964_8799.n29 76.9909
R168 a_n8964_8799.n267 a_n8964_8799.n99 7.32118
R169 a_n8964_8799.n98 a_n8964_8799.n28 78.3454
R170 a_n8964_8799.n28 a_n8964_8799.n97 72.8951
R171 a_n8964_8799.n96 a_n8964_8799.n30 70.1674
R172 a_n8964_8799.n270 a_n8964_8799.n96 20.9683
R173 a_n8964_8799.n30 a_n8964_8799.n95 72.3034
R174 a_n8964_8799.n95 a_n8964_8799.n262 16.6962
R175 a_n8964_8799.n94 a_n8964_8799.n31 77.6622
R176 a_n8964_8799.n271 a_n8964_8799.n94 5.97853
R177 a_n8964_8799.n93 a_n8964_8799.n31 77.6622
R178 a_n8964_8799.n32 a_n8964_8799.n92 72.3034
R179 a_n8964_8799.n91 a_n8964_8799.n32 70.1674
R180 a_n8964_8799.n274 a_n8964_8799.n91 20.9683
R181 a_n8964_8799.n34 a_n8964_8799.n90 72.8951
R182 a_n8964_8799.n90 a_n8964_8799.n260 15.5127
R183 a_n8964_8799.n89 a_n8964_8799.n34 78.3454
R184 a_n8964_8799.n275 a_n8964_8799.n89 4.61226
R185 a_n8964_8799.n88 a_n8964_8799.n33 76.9909
R186 a_n8964_8799.n33 a_n8964_8799.n87 71.7212
R187 a_n8964_8799.n277 a_n8964_8799.n86 20.9683
R188 a_n8964_8799.n35 a_n8964_8799.n86 70.1674
R189 a_n8964_8799.n21 a_n8964_8799.n115 70.1674
R190 a_n8964_8799.n179 a_n8964_8799.n115 20.9683
R191 a_n8964_8799.n114 a_n8964_8799.n21 71.7212
R192 a_n8964_8799.n114 a_n8964_8799.n161 17.8606
R193 a_n8964_8799.n20 a_n8964_8799.n113 76.9909
R194 a_n8964_8799.n178 a_n8964_8799.n113 7.32118
R195 a_n8964_8799.n112 a_n8964_8799.n20 78.3454
R196 a_n8964_8799.n22 a_n8964_8799.n111 72.8951
R197 a_n8964_8799.n110 a_n8964_8799.n22 70.1674
R198 a_n8964_8799.n110 a_n8964_8799.n162 20.9683
R199 a_n8964_8799.n23 a_n8964_8799.n109 72.3034
R200 a_n8964_8799.n174 a_n8964_8799.n109 16.6962
R201 a_n8964_8799.n108 a_n8964_8799.n23 77.6622
R202 a_n8964_8799.n108 a_n8964_8799.n163 5.97853
R203 a_n8964_8799.n24 a_n8964_8799.n107 77.6622
R204 a_n8964_8799.n106 a_n8964_8799.n24 72.3034
R205 a_n8964_8799.n25 a_n8964_8799.n105 70.1674
R206 a_n8964_8799.n170 a_n8964_8799.n105 20.9683
R207 a_n8964_8799.n104 a_n8964_8799.n25 72.8951
R208 a_n8964_8799.n104 a_n8964_8799.n164 15.5127
R209 a_n8964_8799.n26 a_n8964_8799.n103 78.3454
R210 a_n8964_8799.n169 a_n8964_8799.n103 4.61226
R211 a_n8964_8799.n102 a_n8964_8799.n26 76.9909
R212 a_n8964_8799.n101 a_n8964_8799.n167 17.8606
R213 a_n8964_8799.n101 a_n8964_8799.n27 71.7212
R214 a_n8964_8799.n13 a_n8964_8799.n130 70.1674
R215 a_n8964_8799.n198 a_n8964_8799.n130 20.9683
R216 a_n8964_8799.n129 a_n8964_8799.n13 71.7212
R217 a_n8964_8799.n129 a_n8964_8799.n180 17.8606
R218 a_n8964_8799.n12 a_n8964_8799.n128 76.9909
R219 a_n8964_8799.n197 a_n8964_8799.n128 7.32118
R220 a_n8964_8799.n127 a_n8964_8799.n12 78.3454
R221 a_n8964_8799.n14 a_n8964_8799.n126 72.8951
R222 a_n8964_8799.n125 a_n8964_8799.n14 70.1674
R223 a_n8964_8799.n125 a_n8964_8799.n181 20.9683
R224 a_n8964_8799.n15 a_n8964_8799.n124 72.3034
R225 a_n8964_8799.n193 a_n8964_8799.n124 16.6962
R226 a_n8964_8799.n123 a_n8964_8799.n15 77.6622
R227 a_n8964_8799.n123 a_n8964_8799.n182 5.97853
R228 a_n8964_8799.n16 a_n8964_8799.n122 77.6622
R229 a_n8964_8799.n121 a_n8964_8799.n16 72.3034
R230 a_n8964_8799.n17 a_n8964_8799.n120 70.1674
R231 a_n8964_8799.n189 a_n8964_8799.n120 20.9683
R232 a_n8964_8799.n119 a_n8964_8799.n17 72.8951
R233 a_n8964_8799.n119 a_n8964_8799.n183 15.5127
R234 a_n8964_8799.n18 a_n8964_8799.n118 78.3454
R235 a_n8964_8799.n188 a_n8964_8799.n118 4.61226
R236 a_n8964_8799.n117 a_n8964_8799.n18 76.9909
R237 a_n8964_8799.n116 a_n8964_8799.n186 17.8606
R238 a_n8964_8799.n116 a_n8964_8799.n19 71.7212
R239 a_n8964_8799.n5 a_n8964_8799.n145 70.1674
R240 a_n8964_8799.n218 a_n8964_8799.n145 20.9683
R241 a_n8964_8799.n144 a_n8964_8799.n5 71.7212
R242 a_n8964_8799.n144 a_n8964_8799.n200 17.8606
R243 a_n8964_8799.n4 a_n8964_8799.n143 76.9909
R244 a_n8964_8799.n217 a_n8964_8799.n143 7.32118
R245 a_n8964_8799.n142 a_n8964_8799.n4 78.3454
R246 a_n8964_8799.n6 a_n8964_8799.n141 72.8951
R247 a_n8964_8799.n140 a_n8964_8799.n6 70.1674
R248 a_n8964_8799.n140 a_n8964_8799.n201 20.9683
R249 a_n8964_8799.n7 a_n8964_8799.n139 72.3034
R250 a_n8964_8799.n213 a_n8964_8799.n139 16.6962
R251 a_n8964_8799.n138 a_n8964_8799.n7 77.6622
R252 a_n8964_8799.n138 a_n8964_8799.n202 5.97853
R253 a_n8964_8799.n8 a_n8964_8799.n137 77.6622
R254 a_n8964_8799.n136 a_n8964_8799.n8 72.3034
R255 a_n8964_8799.n9 a_n8964_8799.n135 70.1674
R256 a_n8964_8799.n209 a_n8964_8799.n135 20.9683
R257 a_n8964_8799.n134 a_n8964_8799.n9 72.8951
R258 a_n8964_8799.n134 a_n8964_8799.n203 15.5127
R259 a_n8964_8799.n10 a_n8964_8799.n133 78.3454
R260 a_n8964_8799.n208 a_n8964_8799.n133 4.61226
R261 a_n8964_8799.n132 a_n8964_8799.n10 76.9909
R262 a_n8964_8799.n131 a_n8964_8799.n206 17.8606
R263 a_n8964_8799.n131 a_n8964_8799.n11 71.7212
R264 a_n8964_8799.n286 a_n8964_8799.n55 98.9632
R265 a_n8964_8799.n52 a_n8964_8799.n146 98.9631
R266 a_n8964_8799.n54 a_n8964_8799.n282 98.6055
R267 a_n8964_8799.n54 a_n8964_8799.n283 98.6055
R268 a_n8964_8799.n55 a_n8964_8799.n284 98.6055
R269 a_n8964_8799.n55 a_n8964_8799.n285 98.6055
R270 a_n8964_8799.n52 a_n8964_8799.n147 98.6055
R271 a_n8964_8799.n52 a_n8964_8799.n148 98.6055
R272 a_n8964_8799.n53 a_n8964_8799.n149 98.6055
R273 a_n8964_8799.n53 a_n8964_8799.n150 98.6055
R274 a_n8964_8799.n3 a_n8964_8799.n151 81.4626
R275 a_n8964_8799.n1 a_n8964_8799.n157 81.4626
R276 a_n8964_8799.n0 a_n8964_8799.n154 81.4626
R277 a_n8964_8799.n2 a_n8964_8799.n159 80.9324
R278 a_n8964_8799.n2 a_n8964_8799.n160 80.9324
R279 a_n8964_8799.n3 a_n8964_8799.n153 80.9324
R280 a_n8964_8799.n3 a_n8964_8799.n152 80.9324
R281 a_n8964_8799.n1 a_n8964_8799.n158 80.9324
R282 a_n8964_8799.n1 a_n8964_8799.n156 80.9324
R283 a_n8964_8799.n0 a_n8964_8799.n155 80.9324
R284 a_n8964_8799.n45 a_n8964_8799.n226 70.4033
R285 a_n8964_8799.n37 a_n8964_8799.n245 70.4033
R286 a_n8964_8799.n29 a_n8964_8799.n265 70.4033
R287 a_n8964_8799.n165 a_n8964_8799.n27 70.4033
R288 a_n8964_8799.n184 a_n8964_8799.n19 70.4033
R289 a_n8964_8799.n204 a_n8964_8799.n11 70.4033
R290 a_n8964_8799.n237 a_n8964_8799.n236 48.2005
R291 a_n8964_8799.n61 a_n8964_8799.n234 20.9683
R292 a_n8964_8799.n233 a_n8964_8799.n232 48.2005
R293 a_n8964_8799.n66 a_n8964_8799.n230 20.9683
R294 a_n8964_8799.n229 a_n8964_8799.n228 48.2005
R295 a_n8964_8799.n256 a_n8964_8799.n255 48.2005
R296 a_n8964_8799.n76 a_n8964_8799.n253 20.9683
R297 a_n8964_8799.n252 a_n8964_8799.n251 48.2005
R298 a_n8964_8799.n81 a_n8964_8799.n249 20.9683
R299 a_n8964_8799.n248 a_n8964_8799.n247 48.2005
R300 a_n8964_8799.n276 a_n8964_8799.n275 48.2005
R301 a_n8964_8799.n91 a_n8964_8799.n273 20.9683
R302 a_n8964_8799.n272 a_n8964_8799.n271 48.2005
R303 a_n8964_8799.n96 a_n8964_8799.n269 20.9683
R304 a_n8964_8799.n268 a_n8964_8799.n267 48.2005
R305 a_n8964_8799.n169 a_n8964_8799.n168 48.2005
R306 a_n8964_8799.n171 a_n8964_8799.n105 20.9683
R307 a_n8964_8799.n173 a_n8964_8799.n163 48.2005
R308 a_n8964_8799.n175 a_n8964_8799.n110 20.9683
R309 a_n8964_8799.n178 a_n8964_8799.n177 48.2005
R310 a_n8964_8799.t40 a_n8964_8799.n115 485.135
R311 a_n8964_8799.n188 a_n8964_8799.n187 48.2005
R312 a_n8964_8799.n190 a_n8964_8799.n120 20.9683
R313 a_n8964_8799.n192 a_n8964_8799.n182 48.2005
R314 a_n8964_8799.n194 a_n8964_8799.n125 20.9683
R315 a_n8964_8799.n197 a_n8964_8799.n196 48.2005
R316 a_n8964_8799.t52 a_n8964_8799.n130 485.135
R317 a_n8964_8799.n208 a_n8964_8799.n207 48.2005
R318 a_n8964_8799.n210 a_n8964_8799.n135 20.9683
R319 a_n8964_8799.n212 a_n8964_8799.n202 48.2005
R320 a_n8964_8799.n214 a_n8964_8799.n140 20.9683
R321 a_n8964_8799.n217 a_n8964_8799.n216 48.2005
R322 a_n8964_8799.t95 a_n8964_8799.n145 485.135
R323 a_n8964_8799.n57 a_n8964_8799.n220 17.8606
R324 a_n8964_8799.n227 a_n8964_8799.n70 25.894
R325 a_n8964_8799.n72 a_n8964_8799.n239 17.8606
R326 a_n8964_8799.n246 a_n8964_8799.n85 25.894
R327 a_n8964_8799.n87 a_n8964_8799.n259 17.8606
R328 a_n8964_8799.n266 a_n8964_8799.n100 25.894
R329 a_n8964_8799.n179 a_n8964_8799.n114 25.894
R330 a_n8964_8799.n198 a_n8964_8799.n129 25.894
R331 a_n8964_8799.n218 a_n8964_8799.n144 25.894
R332 a_n8964_8799.n68 a_n8964_8799.n224 43.3183
R333 a_n8964_8799.n83 a_n8964_8799.n243 43.3183
R334 a_n8964_8799.n98 a_n8964_8799.n263 43.3183
R335 a_n8964_8799.n176 a_n8964_8799.n112 43.3183
R336 a_n8964_8799.n195 a_n8964_8799.n127 43.3183
R337 a_n8964_8799.n215 a_n8964_8799.n142 43.3183
R338 a_n8964_8799.n62 a_n8964_8799.n222 16.6962
R339 a_n8964_8799.n231 a_n8964_8799.n65 27.6507
R340 a_n8964_8799.n77 a_n8964_8799.n241 16.6962
R341 a_n8964_8799.n250 a_n8964_8799.n80 27.6507
R342 a_n8964_8799.n92 a_n8964_8799.n261 16.6962
R343 a_n8964_8799.n270 a_n8964_8799.n95 27.6507
R344 a_n8964_8799.n172 a_n8964_8799.n106 16.6962
R345 a_n8964_8799.n162 a_n8964_8799.n109 27.6507
R346 a_n8964_8799.n191 a_n8964_8799.n121 16.6962
R347 a_n8964_8799.n181 a_n8964_8799.n124 27.6507
R348 a_n8964_8799.n211 a_n8964_8799.n136 16.6962
R349 a_n8964_8799.n201 a_n8964_8799.n139 27.6507
R350 a_n8964_8799.n63 a_n8964_8799.n222 41.7634
R351 a_n8964_8799.n78 a_n8964_8799.n241 41.7634
R352 a_n8964_8799.n93 a_n8964_8799.n261 41.7634
R353 a_n8964_8799.n107 a_n8964_8799.n172 41.7634
R354 a_n8964_8799.n122 a_n8964_8799.n191 41.7634
R355 a_n8964_8799.n137 a_n8964_8799.n211 41.7634
R356 a_n8964_8799.n235 a_n8964_8799.n60 29.3885
R357 a_n8964_8799.n67 a_n8964_8799.n224 15.5127
R358 a_n8964_8799.n254 a_n8964_8799.n75 29.3885
R359 a_n8964_8799.n82 a_n8964_8799.n243 15.5127
R360 a_n8964_8799.n274 a_n8964_8799.n90 29.3885
R361 a_n8964_8799.n97 a_n8964_8799.n263 15.5127
R362 a_n8964_8799.n170 a_n8964_8799.n104 29.3885
R363 a_n8964_8799.n176 a_n8964_8799.n111 15.5127
R364 a_n8964_8799.n189 a_n8964_8799.n119 29.3885
R365 a_n8964_8799.n195 a_n8964_8799.n126 15.5127
R366 a_n8964_8799.n209 a_n8964_8799.n134 29.3885
R367 a_n8964_8799.n215 a_n8964_8799.n141 15.5127
R368 a_n8964_8799.n2 a_n8964_8799.n1 33.5285
R369 a_n8964_8799.n281 a_n8964_8799.n53 33.0756
R370 a_n8964_8799.n58 a_n8964_8799.n220 40.1848
R371 a_n8964_8799.n73 a_n8964_8799.n239 40.1848
R372 a_n8964_8799.n88 a_n8964_8799.n259 40.1848
R373 a_n8964_8799.n167 a_n8964_8799.n102 40.1848
R374 a_n8964_8799.n186 a_n8964_8799.n117 40.1848
R375 a_n8964_8799.n206 a_n8964_8799.n132 40.1848
R376 a_n8964_8799.n227 a_n8964_8799.n226 20.9576
R377 a_n8964_8799.n246 a_n8964_8799.n245 20.9576
R378 a_n8964_8799.n266 a_n8964_8799.n265 20.9576
R379 a_n8964_8799.n166 a_n8964_8799.n165 20.9576
R380 a_n8964_8799.n185 a_n8964_8799.n184 20.9576
R381 a_n8964_8799.n205 a_n8964_8799.n204 20.9576
R382 a_n8964_8799.n54 a_n8964_8799.n281 19.6671
R383 a_n8964_8799.n58 a_n8964_8799.n237 7.32118
R384 a_n8964_8799.n69 a_n8964_8799.n225 40.1848
R385 a_n8964_8799.n73 a_n8964_8799.n256 7.32118
R386 a_n8964_8799.n84 a_n8964_8799.n244 40.1848
R387 a_n8964_8799.n88 a_n8964_8799.n276 7.32118
R388 a_n8964_8799.n99 a_n8964_8799.n264 40.1848
R389 a_n8964_8799.n168 a_n8964_8799.n102 7.32118
R390 a_n8964_8799.n161 a_n8964_8799.n113 40.1848
R391 a_n8964_8799.n187 a_n8964_8799.n117 7.32118
R392 a_n8964_8799.n180 a_n8964_8799.n128 40.1848
R393 a_n8964_8799.n207 a_n8964_8799.n132 7.32118
R394 a_n8964_8799.n200 a_n8964_8799.n143 40.1848
R395 a_n8964_8799.n230 a_n8964_8799.n67 29.3885
R396 a_n8964_8799.n249 a_n8964_8799.n82 29.3885
R397 a_n8964_8799.n269 a_n8964_8799.n97 29.3885
R398 a_n8964_8799.n111 a_n8964_8799.n175 29.3885
R399 a_n8964_8799.n126 a_n8964_8799.n194 29.3885
R400 a_n8964_8799.n141 a_n8964_8799.n214 29.3885
R401 a_n8964_8799.n63 a_n8964_8799.n233 5.97853
R402 a_n8964_8799.n64 a_n8964_8799.n223 41.7634
R403 a_n8964_8799.n78 a_n8964_8799.n252 5.97853
R404 a_n8964_8799.n79 a_n8964_8799.n242 41.7634
R405 a_n8964_8799.n93 a_n8964_8799.n272 5.97853
R406 a_n8964_8799.n94 a_n8964_8799.n262 41.7634
R407 a_n8964_8799.n173 a_n8964_8799.n107 5.97853
R408 a_n8964_8799.n174 a_n8964_8799.n108 41.7634
R409 a_n8964_8799.n192 a_n8964_8799.n122 5.97853
R410 a_n8964_8799.n193 a_n8964_8799.n123 41.7634
R411 a_n8964_8799.n212 a_n8964_8799.n137 5.97853
R412 a_n8964_8799.n213 a_n8964_8799.n138 41.7634
R413 a_n8964_8799.n280 a_n8964_8799.n3 12.3339
R414 a_n8964_8799.n281 a_n8964_8799.n280 11.4887
R415 a_n8964_8799.n234 a_n8964_8799.n62 27.6507
R416 a_n8964_8799.n253 a_n8964_8799.n77 27.6507
R417 a_n8964_8799.n273 a_n8964_8799.n92 27.6507
R418 a_n8964_8799.n171 a_n8964_8799.n106 27.6507
R419 a_n8964_8799.n190 a_n8964_8799.n121 27.6507
R420 a_n8964_8799.n210 a_n8964_8799.n136 27.6507
R421 a_n8964_8799.n59 a_n8964_8799.n221 43.3183
R422 a_n8964_8799.n68 a_n8964_8799.n229 4.61226
R423 a_n8964_8799.n74 a_n8964_8799.n240 43.3183
R424 a_n8964_8799.n83 a_n8964_8799.n248 4.61226
R425 a_n8964_8799.n89 a_n8964_8799.n260 43.3183
R426 a_n8964_8799.n98 a_n8964_8799.n268 4.61226
R427 a_n8964_8799.n164 a_n8964_8799.n103 43.3183
R428 a_n8964_8799.n177 a_n8964_8799.n112 4.61226
R429 a_n8964_8799.n183 a_n8964_8799.n118 43.3183
R430 a_n8964_8799.n196 a_n8964_8799.n127 4.61226
R431 a_n8964_8799.n203 a_n8964_8799.n133 43.3183
R432 a_n8964_8799.n216 a_n8964_8799.n142 4.61226
R433 a_n8964_8799.n258 a_n8964_8799.n51 9.04406
R434 a_n8964_8799.n199 a_n8964_8799.n21 9.04406
R435 a_n8964_8799.n238 a_n8964_8799.n57 25.894
R436 a_n8964_8799.n257 a_n8964_8799.n72 25.894
R437 a_n8964_8799.n277 a_n8964_8799.n87 25.894
R438 a_n8964_8799.n101 a_n8964_8799.n166 25.894
R439 a_n8964_8799.n116 a_n8964_8799.n185 25.894
R440 a_n8964_8799.n131 a_n8964_8799.n205 25.894
R441 a_n8964_8799.n279 a_n8964_8799.n219 7.10923
R442 a_n8964_8799.n279 a_n8964_8799.n278 6.68968
R443 a_n8964_8799.n258 a_n8964_8799.n43 4.93611
R444 a_n8964_8799.n278 a_n8964_8799.n35 4.93611
R445 a_n8964_8799.n199 a_n8964_8799.n13 4.93611
R446 a_n8964_8799.n219 a_n8964_8799.n5 4.93611
R447 a_n8964_8799.n278 a_n8964_8799.n258 4.10845
R448 a_n8964_8799.n219 a_n8964_8799.n199 4.10845
R449 a_n8964_8799.n282 a_n8964_8799.t38 3.61217
R450 a_n8964_8799.n282 a_n8964_8799.t25 3.61217
R451 a_n8964_8799.n283 a_n8964_8799.t31 3.61217
R452 a_n8964_8799.n283 a_n8964_8799.t28 3.61217
R453 a_n8964_8799.n284 a_n8964_8799.t5 3.61217
R454 a_n8964_8799.n284 a_n8964_8799.t35 3.61217
R455 a_n8964_8799.n285 a_n8964_8799.t27 3.61217
R456 a_n8964_8799.n285 a_n8964_8799.t17 3.61217
R457 a_n8964_8799.n146 a_n8964_8799.t4 3.61217
R458 a_n8964_8799.n146 a_n8964_8799.t29 3.61217
R459 a_n8964_8799.n147 a_n8964_8799.t21 3.61217
R460 a_n8964_8799.n147 a_n8964_8799.t7 3.61217
R461 a_n8964_8799.n148 a_n8964_8799.t1 3.61217
R462 a_n8964_8799.n148 a_n8964_8799.t2 3.61217
R463 a_n8964_8799.n149 a_n8964_8799.t34 3.61217
R464 a_n8964_8799.n149 a_n8964_8799.t24 3.61217
R465 a_n8964_8799.n150 a_n8964_8799.t16 3.61217
R466 a_n8964_8799.n150 a_n8964_8799.t22 3.61217
R467 a_n8964_8799.t0 a_n8964_8799.n286 3.61217
R468 a_n8964_8799.n286 a_n8964_8799.t8 3.61217
R469 a_n8964_8799.n280 a_n8964_8799.n279 3.4105
R470 a_n8964_8799.n159 a_n8964_8799.t39 2.82907
R471 a_n8964_8799.n159 a_n8964_8799.t10 2.82907
R472 a_n8964_8799.n160 a_n8964_8799.t19 2.82907
R473 a_n8964_8799.n160 a_n8964_8799.t30 2.82907
R474 a_n8964_8799.n153 a_n8964_8799.t3 2.82907
R475 a_n8964_8799.n153 a_n8964_8799.t37 2.82907
R476 a_n8964_8799.n152 a_n8964_8799.t15 2.82907
R477 a_n8964_8799.n152 a_n8964_8799.t18 2.82907
R478 a_n8964_8799.n151 a_n8964_8799.t20 2.82907
R479 a_n8964_8799.n151 a_n8964_8799.t26 2.82907
R480 a_n8964_8799.n157 a_n8964_8799.t32 2.82907
R481 a_n8964_8799.n157 a_n8964_8799.t9 2.82907
R482 a_n8964_8799.n158 a_n8964_8799.t11 2.82907
R483 a_n8964_8799.n158 a_n8964_8799.t13 2.82907
R484 a_n8964_8799.n156 a_n8964_8799.t14 2.82907
R485 a_n8964_8799.n156 a_n8964_8799.t23 2.82907
R486 a_n8964_8799.n155 a_n8964_8799.t6 2.82907
R487 a_n8964_8799.n155 a_n8964_8799.t12 2.82907
R488 a_n8964_8799.n154 a_n8964_8799.t36 2.82907
R489 a_n8964_8799.n154 a_n8964_8799.t33 2.82907
R490 a_n8964_8799.n3 a_n8964_8799.n2 1.59102
R491 a_n8964_8799.n45 a_n8964_8799.n44 1.13686
R492 a_n8964_8799.n37 a_n8964_8799.n36 1.13686
R493 a_n8964_8799.n29 a_n8964_8799.n28 1.13686
R494 a_n8964_8799.n21 a_n8964_8799.n20 1.13686
R495 a_n8964_8799.n13 a_n8964_8799.n12 1.13686
R496 a_n8964_8799.n5 a_n8964_8799.n4 1.13686
R497 a_n8964_8799.n55 a_n8964_8799.n54 1.07378
R498 a_n8964_8799.n53 a_n8964_8799.n52 1.07378
R499 a_n8964_8799.n1 a_n8964_8799.n0 1.06084
R500 a_n8964_8799.n50 a_n8964_8799.n49 0.758076
R501 a_n8964_8799.n50 a_n8964_8799.n48 0.758076
R502 a_n8964_8799.n48 a_n8964_8799.n47 0.758076
R503 a_n8964_8799.n47 a_n8964_8799.n46 0.758076
R504 a_n8964_8799.n44 a_n8964_8799.n46 0.758076
R505 a_n8964_8799.n42 a_n8964_8799.n41 0.758076
R506 a_n8964_8799.n42 a_n8964_8799.n40 0.758076
R507 a_n8964_8799.n40 a_n8964_8799.n39 0.758076
R508 a_n8964_8799.n39 a_n8964_8799.n38 0.758076
R509 a_n8964_8799.n36 a_n8964_8799.n38 0.758076
R510 a_n8964_8799.n34 a_n8964_8799.n33 0.758076
R511 a_n8964_8799.n34 a_n8964_8799.n32 0.758076
R512 a_n8964_8799.n32 a_n8964_8799.n31 0.758076
R513 a_n8964_8799.n31 a_n8964_8799.n30 0.758076
R514 a_n8964_8799.n28 a_n8964_8799.n30 0.758076
R515 a_n8964_8799.n25 a_n8964_8799.n26 0.758076
R516 a_n8964_8799.n24 a_n8964_8799.n25 0.758076
R517 a_n8964_8799.n23 a_n8964_8799.n24 0.758076
R518 a_n8964_8799.n22 a_n8964_8799.n23 0.758076
R519 a_n8964_8799.n20 a_n8964_8799.n22 0.758076
R520 a_n8964_8799.n17 a_n8964_8799.n18 0.758076
R521 a_n8964_8799.n16 a_n8964_8799.n17 0.758076
R522 a_n8964_8799.n15 a_n8964_8799.n16 0.758076
R523 a_n8964_8799.n14 a_n8964_8799.n15 0.758076
R524 a_n8964_8799.n12 a_n8964_8799.n14 0.758076
R525 a_n8964_8799.n9 a_n8964_8799.n10 0.758076
R526 a_n8964_8799.n8 a_n8964_8799.n9 0.758076
R527 a_n8964_8799.n7 a_n8964_8799.n8 0.758076
R528 a_n8964_8799.n6 a_n8964_8799.n7 0.758076
R529 a_n8964_8799.n4 a_n8964_8799.n6 0.758076
R530 a_n8964_8799.n10 a_n8964_8799.n11 0.568682
R531 a_n8964_8799.n18 a_n8964_8799.n19 0.568682
R532 a_n8964_8799.n26 a_n8964_8799.n27 0.568682
R533 a_n8964_8799.n33 a_n8964_8799.n35 0.568682
R534 a_n8964_8799.n41 a_n8964_8799.n43 0.568682
R535 a_n8964_8799.n49 a_n8964_8799.n51 0.568682
R536 vdd.n327 vdd.n291 756.745
R537 vdd.n268 vdd.n232 756.745
R538 vdd.n225 vdd.n189 756.745
R539 vdd.n166 vdd.n130 756.745
R540 vdd.n124 vdd.n88 756.745
R541 vdd.n65 vdd.n29 756.745
R542 vdd.n1826 vdd.n1790 756.745
R543 vdd.n1885 vdd.n1849 756.745
R544 vdd.n1724 vdd.n1688 756.745
R545 vdd.n1783 vdd.n1747 756.745
R546 vdd.n1623 vdd.n1587 756.745
R547 vdd.n1682 vdd.n1646 756.745
R548 vdd.n1136 vdd.t29 640.208
R549 vdd.n997 vdd.t67 640.208
R550 vdd.n1130 vdd.t94 640.208
R551 vdd.n988 vdd.t91 640.208
R552 vdd.n885 vdd.t40 640.208
R553 vdd.n2761 vdd.t85 640.208
R554 vdd.n832 vdd.t54 640.208
R555 vdd.n2830 vdd.t71 640.208
R556 vdd.n799 vdd.t25 640.208
R557 vdd.n1058 vdd.t81 640.208
R558 vdd.n1397 vdd.t63 592.009
R559 vdd.n1435 vdd.t75 592.009
R560 vdd.n1331 vdd.t88 592.009
R561 vdd.n2200 vdd.t47 592.009
R562 vdd.n2050 vdd.t57 592.009
R563 vdd.n2010 vdd.t78 592.009
R564 vdd.n426 vdd.t60 592.009
R565 vdd.n440 vdd.t33 592.009
R566 vdd.n452 vdd.t51 592.009
R567 vdd.n768 vdd.t21 592.009
R568 vdd.n3366 vdd.t37 592.009
R569 vdd.n688 vdd.t44 592.009
R570 vdd.n328 vdd.n327 585
R571 vdd.n326 vdd.n293 585
R572 vdd.n325 vdd.n324 585
R573 vdd.n296 vdd.n294 585
R574 vdd.n319 vdd.n318 585
R575 vdd.n317 vdd.n316 585
R576 vdd.n300 vdd.n299 585
R577 vdd.n311 vdd.n310 585
R578 vdd.n309 vdd.n308 585
R579 vdd.n304 vdd.n303 585
R580 vdd.n269 vdd.n268 585
R581 vdd.n267 vdd.n234 585
R582 vdd.n266 vdd.n265 585
R583 vdd.n237 vdd.n235 585
R584 vdd.n260 vdd.n259 585
R585 vdd.n258 vdd.n257 585
R586 vdd.n241 vdd.n240 585
R587 vdd.n252 vdd.n251 585
R588 vdd.n250 vdd.n249 585
R589 vdd.n245 vdd.n244 585
R590 vdd.n226 vdd.n225 585
R591 vdd.n224 vdd.n191 585
R592 vdd.n223 vdd.n222 585
R593 vdd.n194 vdd.n192 585
R594 vdd.n217 vdd.n216 585
R595 vdd.n215 vdd.n214 585
R596 vdd.n198 vdd.n197 585
R597 vdd.n209 vdd.n208 585
R598 vdd.n207 vdd.n206 585
R599 vdd.n202 vdd.n201 585
R600 vdd.n167 vdd.n166 585
R601 vdd.n165 vdd.n132 585
R602 vdd.n164 vdd.n163 585
R603 vdd.n135 vdd.n133 585
R604 vdd.n158 vdd.n157 585
R605 vdd.n156 vdd.n155 585
R606 vdd.n139 vdd.n138 585
R607 vdd.n150 vdd.n149 585
R608 vdd.n148 vdd.n147 585
R609 vdd.n143 vdd.n142 585
R610 vdd.n125 vdd.n124 585
R611 vdd.n123 vdd.n90 585
R612 vdd.n122 vdd.n121 585
R613 vdd.n93 vdd.n91 585
R614 vdd.n116 vdd.n115 585
R615 vdd.n114 vdd.n113 585
R616 vdd.n97 vdd.n96 585
R617 vdd.n108 vdd.n107 585
R618 vdd.n106 vdd.n105 585
R619 vdd.n101 vdd.n100 585
R620 vdd.n66 vdd.n65 585
R621 vdd.n64 vdd.n31 585
R622 vdd.n63 vdd.n62 585
R623 vdd.n34 vdd.n32 585
R624 vdd.n57 vdd.n56 585
R625 vdd.n55 vdd.n54 585
R626 vdd.n38 vdd.n37 585
R627 vdd.n49 vdd.n48 585
R628 vdd.n47 vdd.n46 585
R629 vdd.n42 vdd.n41 585
R630 vdd.n1827 vdd.n1826 585
R631 vdd.n1825 vdd.n1792 585
R632 vdd.n1824 vdd.n1823 585
R633 vdd.n1795 vdd.n1793 585
R634 vdd.n1818 vdd.n1817 585
R635 vdd.n1816 vdd.n1815 585
R636 vdd.n1799 vdd.n1798 585
R637 vdd.n1810 vdd.n1809 585
R638 vdd.n1808 vdd.n1807 585
R639 vdd.n1803 vdd.n1802 585
R640 vdd.n1886 vdd.n1885 585
R641 vdd.n1884 vdd.n1851 585
R642 vdd.n1883 vdd.n1882 585
R643 vdd.n1854 vdd.n1852 585
R644 vdd.n1877 vdd.n1876 585
R645 vdd.n1875 vdd.n1874 585
R646 vdd.n1858 vdd.n1857 585
R647 vdd.n1869 vdd.n1868 585
R648 vdd.n1867 vdd.n1866 585
R649 vdd.n1862 vdd.n1861 585
R650 vdd.n1725 vdd.n1724 585
R651 vdd.n1723 vdd.n1690 585
R652 vdd.n1722 vdd.n1721 585
R653 vdd.n1693 vdd.n1691 585
R654 vdd.n1716 vdd.n1715 585
R655 vdd.n1714 vdd.n1713 585
R656 vdd.n1697 vdd.n1696 585
R657 vdd.n1708 vdd.n1707 585
R658 vdd.n1706 vdd.n1705 585
R659 vdd.n1701 vdd.n1700 585
R660 vdd.n1784 vdd.n1783 585
R661 vdd.n1782 vdd.n1749 585
R662 vdd.n1781 vdd.n1780 585
R663 vdd.n1752 vdd.n1750 585
R664 vdd.n1775 vdd.n1774 585
R665 vdd.n1773 vdd.n1772 585
R666 vdd.n1756 vdd.n1755 585
R667 vdd.n1767 vdd.n1766 585
R668 vdd.n1765 vdd.n1764 585
R669 vdd.n1760 vdd.n1759 585
R670 vdd.n1624 vdd.n1623 585
R671 vdd.n1622 vdd.n1589 585
R672 vdd.n1621 vdd.n1620 585
R673 vdd.n1592 vdd.n1590 585
R674 vdd.n1615 vdd.n1614 585
R675 vdd.n1613 vdd.n1612 585
R676 vdd.n1596 vdd.n1595 585
R677 vdd.n1607 vdd.n1606 585
R678 vdd.n1605 vdd.n1604 585
R679 vdd.n1600 vdd.n1599 585
R680 vdd.n1683 vdd.n1682 585
R681 vdd.n1681 vdd.n1648 585
R682 vdd.n1680 vdd.n1679 585
R683 vdd.n1651 vdd.n1649 585
R684 vdd.n1674 vdd.n1673 585
R685 vdd.n1672 vdd.n1671 585
R686 vdd.n1655 vdd.n1654 585
R687 vdd.n1666 vdd.n1665 585
R688 vdd.n1664 vdd.n1663 585
R689 vdd.n1659 vdd.n1658 585
R690 vdd.n3538 vdd.n392 509.269
R691 vdd.n3534 vdd.n393 509.269
R692 vdd.n3406 vdd.n685 509.269
R693 vdd.n3403 vdd.n684 509.269
R694 vdd.n2195 vdd.n1155 509.269
R695 vdd.n2198 vdd.n2197 509.269
R696 vdd.n1304 vdd.n1268 509.269
R697 vdd.n1500 vdd.n1269 509.269
R698 vdd.n305 vdd.t180 329.043
R699 vdd.n246 vdd.t221 329.043
R700 vdd.n203 vdd.t160 329.043
R701 vdd.n144 vdd.t201 329.043
R702 vdd.n102 vdd.t244 329.043
R703 vdd.n43 vdd.t270 329.043
R704 vdd.n1804 vdd.t300 329.043
R705 vdd.n1863 vdd.t249 329.043
R706 vdd.n1702 vdd.t288 329.043
R707 vdd.n1761 vdd.t237 329.043
R708 vdd.n1601 vdd.t241 329.043
R709 vdd.n1660 vdd.t246 329.043
R710 vdd.n1397 vdd.t66 319.788
R711 vdd.n1435 vdd.t77 319.788
R712 vdd.n1331 vdd.t90 319.788
R713 vdd.n2200 vdd.t49 319.788
R714 vdd.n2050 vdd.t58 319.788
R715 vdd.n2010 vdd.t79 319.788
R716 vdd.n426 vdd.t61 319.788
R717 vdd.n440 vdd.t35 319.788
R718 vdd.n452 vdd.t52 319.788
R719 vdd.n768 vdd.t24 319.788
R720 vdd.n3366 vdd.t39 319.788
R721 vdd.n688 vdd.t46 319.788
R722 vdd.n1398 vdd.t65 303.69
R723 vdd.n1436 vdd.t76 303.69
R724 vdd.n1332 vdd.t89 303.69
R725 vdd.n2201 vdd.t50 303.69
R726 vdd.n2051 vdd.t59 303.69
R727 vdd.n2011 vdd.t80 303.69
R728 vdd.n427 vdd.t62 303.69
R729 vdd.n441 vdd.t36 303.69
R730 vdd.n453 vdd.t53 303.69
R731 vdd.n769 vdd.t23 303.69
R732 vdd.n3367 vdd.t38 303.69
R733 vdd.n689 vdd.t45 303.69
R734 vdd.n3016 vdd.n947 285.366
R735 vdd.n3240 vdd.n809 285.366
R736 vdd.n3177 vdd.n806 285.366
R737 vdd.n2895 vdd.n944 285.366
R738 vdd.n2725 vdd.n985 285.366
R739 vdd.n2656 vdd.n2655 285.366
R740 vdd.n2396 vdd.n1111 285.366
R741 vdd.n2466 vdd.n1113 285.366
R742 vdd.n3156 vdd.n807 285.366
R743 vdd.n3243 vdd.n3242 285.366
R744 vdd.n3009 vdd.n945 285.366
R745 vdd.n3018 vdd.n943 285.366
R746 vdd.n2653 vdd.n995 285.366
R747 vdd.n993 vdd.n967 285.366
R748 vdd.n2282 vdd.n1112 285.366
R749 vdd.n2468 vdd.n1109 285.366
R750 vdd.n1153 vdd.n1110 216.982
R751 vdd.n3405 vdd.n692 216.982
R752 vdd.n3158 vdd.n807 185
R753 vdd.n3241 vdd.n807 185
R754 vdd.n3160 vdd.n3159 185
R755 vdd.n3159 vdd.n805 185
R756 vdd.n3161 vdd.n839 185
R757 vdd.n3171 vdd.n839 185
R758 vdd.n3162 vdd.n848 185
R759 vdd.n848 vdd.n846 185
R760 vdd.n3164 vdd.n3163 185
R761 vdd.n3165 vdd.n3164 185
R762 vdd.n3117 vdd.n847 185
R763 vdd.n847 vdd.n843 185
R764 vdd.n3116 vdd.n3115 185
R765 vdd.n3115 vdd.n3114 185
R766 vdd.n850 vdd.n849 185
R767 vdd.n851 vdd.n850 185
R768 vdd.n3107 vdd.n3106 185
R769 vdd.n3108 vdd.n3107 185
R770 vdd.n3105 vdd.n859 185
R771 vdd.n864 vdd.n859 185
R772 vdd.n3104 vdd.n3103 185
R773 vdd.n3103 vdd.n3102 185
R774 vdd.n861 vdd.n860 185
R775 vdd.n870 vdd.n861 185
R776 vdd.n3095 vdd.n3094 185
R777 vdd.n3096 vdd.n3095 185
R778 vdd.n3093 vdd.n871 185
R779 vdd.n877 vdd.n871 185
R780 vdd.n3092 vdd.n3091 185
R781 vdd.n3091 vdd.n3090 185
R782 vdd.n873 vdd.n872 185
R783 vdd.n874 vdd.n873 185
R784 vdd.n3083 vdd.n3082 185
R785 vdd.n3084 vdd.n3083 185
R786 vdd.n3081 vdd.n884 185
R787 vdd.n884 vdd.n881 185
R788 vdd.n3079 vdd.n3078 185
R789 vdd.n3078 vdd.n3077 185
R790 vdd.n887 vdd.n886 185
R791 vdd.n888 vdd.n887 185
R792 vdd.n3070 vdd.n3069 185
R793 vdd.n3071 vdd.n3070 185
R794 vdd.n3068 vdd.n896 185
R795 vdd.n901 vdd.n896 185
R796 vdd.n3067 vdd.n3066 185
R797 vdd.n3066 vdd.n3065 185
R798 vdd.n898 vdd.n897 185
R799 vdd.n2977 vdd.n898 185
R800 vdd.n3058 vdd.n3057 185
R801 vdd.n3059 vdd.n3058 185
R802 vdd.n3056 vdd.n908 185
R803 vdd.n908 vdd.n905 185
R804 vdd.n3055 vdd.n3054 185
R805 vdd.n3054 vdd.n3053 185
R806 vdd.n910 vdd.n909 185
R807 vdd.n911 vdd.n910 185
R808 vdd.n3046 vdd.n3045 185
R809 vdd.n3047 vdd.n3046 185
R810 vdd.n3044 vdd.n919 185
R811 vdd.n2989 vdd.n919 185
R812 vdd.n3043 vdd.n3042 185
R813 vdd.n3042 vdd.n3041 185
R814 vdd.n921 vdd.n920 185
R815 vdd.n930 vdd.n921 185
R816 vdd.n3034 vdd.n3033 185
R817 vdd.n3035 vdd.n3034 185
R818 vdd.n3032 vdd.n931 185
R819 vdd.n931 vdd.n927 185
R820 vdd.n3031 vdd.n3030 185
R821 vdd.n3030 vdd.n3029 185
R822 vdd.n933 vdd.n932 185
R823 vdd.n3001 vdd.n933 185
R824 vdd.n3022 vdd.n3021 185
R825 vdd.n3023 vdd.n3022 185
R826 vdd.n3020 vdd.n941 185
R827 vdd.n946 vdd.n941 185
R828 vdd.n3019 vdd.n3018 185
R829 vdd.n3018 vdd.n3017 185
R830 vdd.n943 vdd.n942 185
R831 vdd.n2765 vdd.n2764 185
R832 vdd.n2767 vdd.n2766 185
R833 vdd.n2769 vdd.n2768 185
R834 vdd.n2771 vdd.n2770 185
R835 vdd.n2773 vdd.n2772 185
R836 vdd.n2775 vdd.n2774 185
R837 vdd.n2777 vdd.n2776 185
R838 vdd.n2779 vdd.n2778 185
R839 vdd.n2781 vdd.n2780 185
R840 vdd.n2783 vdd.n2782 185
R841 vdd.n2785 vdd.n2784 185
R842 vdd.n2787 vdd.n2786 185
R843 vdd.n2789 vdd.n2788 185
R844 vdd.n2791 vdd.n2790 185
R845 vdd.n2793 vdd.n2792 185
R846 vdd.n2795 vdd.n2794 185
R847 vdd.n2797 vdd.n2796 185
R848 vdd.n2799 vdd.n2798 185
R849 vdd.n2801 vdd.n2800 185
R850 vdd.n2803 vdd.n2802 185
R851 vdd.n2805 vdd.n2804 185
R852 vdd.n2807 vdd.n2806 185
R853 vdd.n2809 vdd.n2808 185
R854 vdd.n2811 vdd.n2810 185
R855 vdd.n2813 vdd.n2812 185
R856 vdd.n2815 vdd.n2814 185
R857 vdd.n2817 vdd.n2816 185
R858 vdd.n2819 vdd.n2818 185
R859 vdd.n2821 vdd.n2820 185
R860 vdd.n2823 vdd.n2822 185
R861 vdd.n2825 vdd.n2824 185
R862 vdd.n2827 vdd.n2826 185
R863 vdd.n2828 vdd.n2760 185
R864 vdd.n3009 vdd.n3008 185
R865 vdd.n3010 vdd.n3009 185
R866 vdd.n3244 vdd.n3243 185
R867 vdd.n3245 vdd.n798 185
R868 vdd.n3247 vdd.n3246 185
R869 vdd.n3249 vdd.n796 185
R870 vdd.n3251 vdd.n3250 185
R871 vdd.n3252 vdd.n795 185
R872 vdd.n3254 vdd.n3253 185
R873 vdd.n3256 vdd.n793 185
R874 vdd.n3258 vdd.n3257 185
R875 vdd.n3259 vdd.n792 185
R876 vdd.n3261 vdd.n3260 185
R877 vdd.n3263 vdd.n790 185
R878 vdd.n3265 vdd.n3264 185
R879 vdd.n3266 vdd.n789 185
R880 vdd.n3268 vdd.n3267 185
R881 vdd.n3270 vdd.n788 185
R882 vdd.n3271 vdd.n786 185
R883 vdd.n3274 vdd.n3273 185
R884 vdd.n787 vdd.n785 185
R885 vdd.n3130 vdd.n3129 185
R886 vdd.n3132 vdd.n3131 185
R887 vdd.n3134 vdd.n3126 185
R888 vdd.n3136 vdd.n3135 185
R889 vdd.n3137 vdd.n3125 185
R890 vdd.n3139 vdd.n3138 185
R891 vdd.n3141 vdd.n3123 185
R892 vdd.n3143 vdd.n3142 185
R893 vdd.n3144 vdd.n3122 185
R894 vdd.n3146 vdd.n3145 185
R895 vdd.n3148 vdd.n3120 185
R896 vdd.n3150 vdd.n3149 185
R897 vdd.n3151 vdd.n3119 185
R898 vdd.n3153 vdd.n3152 185
R899 vdd.n3155 vdd.n3118 185
R900 vdd.n3157 vdd.n3156 185
R901 vdd.n3156 vdd.n692 185
R902 vdd.n3242 vdd.n802 185
R903 vdd.n3242 vdd.n3241 185
R904 vdd.n2908 vdd.n804 185
R905 vdd.n805 vdd.n804 185
R906 vdd.n2909 vdd.n838 185
R907 vdd.n3171 vdd.n838 185
R908 vdd.n2911 vdd.n2910 185
R909 vdd.n2910 vdd.n846 185
R910 vdd.n2912 vdd.n845 185
R911 vdd.n3165 vdd.n845 185
R912 vdd.n2914 vdd.n2913 185
R913 vdd.n2913 vdd.n843 185
R914 vdd.n2915 vdd.n853 185
R915 vdd.n3114 vdd.n853 185
R916 vdd.n2917 vdd.n2916 185
R917 vdd.n2916 vdd.n851 185
R918 vdd.n2918 vdd.n858 185
R919 vdd.n3108 vdd.n858 185
R920 vdd.n2920 vdd.n2919 185
R921 vdd.n2919 vdd.n864 185
R922 vdd.n2921 vdd.n863 185
R923 vdd.n3102 vdd.n863 185
R924 vdd.n2923 vdd.n2922 185
R925 vdd.n2922 vdd.n870 185
R926 vdd.n2924 vdd.n869 185
R927 vdd.n3096 vdd.n869 185
R928 vdd.n2926 vdd.n2925 185
R929 vdd.n2925 vdd.n877 185
R930 vdd.n2927 vdd.n876 185
R931 vdd.n3090 vdd.n876 185
R932 vdd.n2929 vdd.n2928 185
R933 vdd.n2928 vdd.n874 185
R934 vdd.n2930 vdd.n883 185
R935 vdd.n3084 vdd.n883 185
R936 vdd.n2932 vdd.n2931 185
R937 vdd.n2931 vdd.n881 185
R938 vdd.n2933 vdd.n890 185
R939 vdd.n3077 vdd.n890 185
R940 vdd.n2935 vdd.n2934 185
R941 vdd.n2934 vdd.n888 185
R942 vdd.n2936 vdd.n895 185
R943 vdd.n3071 vdd.n895 185
R944 vdd.n2938 vdd.n2937 185
R945 vdd.n2937 vdd.n901 185
R946 vdd.n2939 vdd.n900 185
R947 vdd.n3065 vdd.n900 185
R948 vdd.n2979 vdd.n2978 185
R949 vdd.n2978 vdd.n2977 185
R950 vdd.n2980 vdd.n907 185
R951 vdd.n3059 vdd.n907 185
R952 vdd.n2982 vdd.n2981 185
R953 vdd.n2981 vdd.n905 185
R954 vdd.n2983 vdd.n913 185
R955 vdd.n3053 vdd.n913 185
R956 vdd.n2985 vdd.n2984 185
R957 vdd.n2984 vdd.n911 185
R958 vdd.n2986 vdd.n918 185
R959 vdd.n3047 vdd.n918 185
R960 vdd.n2988 vdd.n2987 185
R961 vdd.n2989 vdd.n2988 185
R962 vdd.n2907 vdd.n923 185
R963 vdd.n3041 vdd.n923 185
R964 vdd.n2906 vdd.n2905 185
R965 vdd.n2905 vdd.n930 185
R966 vdd.n2904 vdd.n929 185
R967 vdd.n3035 vdd.n929 185
R968 vdd.n2903 vdd.n2902 185
R969 vdd.n2902 vdd.n927 185
R970 vdd.n2829 vdd.n935 185
R971 vdd.n3029 vdd.n935 185
R972 vdd.n3003 vdd.n3002 185
R973 vdd.n3002 vdd.n3001 185
R974 vdd.n3004 vdd.n940 185
R975 vdd.n3023 vdd.n940 185
R976 vdd.n3006 vdd.n3005 185
R977 vdd.n3005 vdd.n946 185
R978 vdd.n3007 vdd.n945 185
R979 vdd.n3017 vdd.n945 185
R980 vdd.n2195 vdd.n2194 185
R981 vdd.n2196 vdd.n2195 185
R982 vdd.n1156 vdd.n1154 185
R983 vdd.n1974 vdd.n1154 185
R984 vdd.n1977 vdd.n1976 185
R985 vdd.n1976 vdd.n1975 185
R986 vdd.n1159 vdd.n1158 185
R987 vdd.n1160 vdd.n1159 185
R988 vdd.n1963 vdd.n1962 185
R989 vdd.n1964 vdd.n1963 185
R990 vdd.n1168 vdd.n1167 185
R991 vdd.n1955 vdd.n1167 185
R992 vdd.n1958 vdd.n1957 185
R993 vdd.n1957 vdd.n1956 185
R994 vdd.n1171 vdd.n1170 185
R995 vdd.n1178 vdd.n1171 185
R996 vdd.n1946 vdd.n1945 185
R997 vdd.n1947 vdd.n1946 185
R998 vdd.n1180 vdd.n1179 185
R999 vdd.n1179 vdd.n1177 185
R1000 vdd.n1941 vdd.n1940 185
R1001 vdd.n1940 vdd.n1939 185
R1002 vdd.n1183 vdd.n1182 185
R1003 vdd.n1184 vdd.n1183 185
R1004 vdd.n1930 vdd.n1929 185
R1005 vdd.n1931 vdd.n1930 185
R1006 vdd.n1191 vdd.n1190 185
R1007 vdd.n1922 vdd.n1190 185
R1008 vdd.n1925 vdd.n1924 185
R1009 vdd.n1924 vdd.n1923 185
R1010 vdd.n1194 vdd.n1193 185
R1011 vdd.n1200 vdd.n1194 185
R1012 vdd.n1913 vdd.n1912 185
R1013 vdd.n1914 vdd.n1913 185
R1014 vdd.n1202 vdd.n1201 185
R1015 vdd.n1905 vdd.n1201 185
R1016 vdd.n1908 vdd.n1907 185
R1017 vdd.n1907 vdd.n1906 185
R1018 vdd.n1205 vdd.n1204 185
R1019 vdd.n1206 vdd.n1205 185
R1020 vdd.n1896 vdd.n1895 185
R1021 vdd.n1897 vdd.n1896 185
R1022 vdd.n1214 vdd.n1213 185
R1023 vdd.n1213 vdd.n1212 185
R1024 vdd.n1584 vdd.n1583 185
R1025 vdd.n1583 vdd.n1582 185
R1026 vdd.n1217 vdd.n1216 185
R1027 vdd.n1223 vdd.n1217 185
R1028 vdd.n1573 vdd.n1572 185
R1029 vdd.n1574 vdd.n1573 185
R1030 vdd.n1225 vdd.n1224 185
R1031 vdd.n1565 vdd.n1224 185
R1032 vdd.n1568 vdd.n1567 185
R1033 vdd.n1567 vdd.n1566 185
R1034 vdd.n1228 vdd.n1227 185
R1035 vdd.n1235 vdd.n1228 185
R1036 vdd.n1556 vdd.n1555 185
R1037 vdd.n1557 vdd.n1556 185
R1038 vdd.n1237 vdd.n1236 185
R1039 vdd.n1236 vdd.n1234 185
R1040 vdd.n1551 vdd.n1550 185
R1041 vdd.n1550 vdd.n1549 185
R1042 vdd.n1240 vdd.n1239 185
R1043 vdd.n1241 vdd.n1240 185
R1044 vdd.n1540 vdd.n1539 185
R1045 vdd.n1541 vdd.n1540 185
R1046 vdd.n1248 vdd.n1247 185
R1047 vdd.n1532 vdd.n1247 185
R1048 vdd.n1535 vdd.n1534 185
R1049 vdd.n1534 vdd.n1533 185
R1050 vdd.n1251 vdd.n1250 185
R1051 vdd.n1257 vdd.n1251 185
R1052 vdd.n1523 vdd.n1522 185
R1053 vdd.n1524 vdd.n1523 185
R1054 vdd.n1259 vdd.n1258 185
R1055 vdd.n1515 vdd.n1258 185
R1056 vdd.n1518 vdd.n1517 185
R1057 vdd.n1517 vdd.n1516 185
R1058 vdd.n1262 vdd.n1261 185
R1059 vdd.n1263 vdd.n1262 185
R1060 vdd.n1506 vdd.n1505 185
R1061 vdd.n1507 vdd.n1506 185
R1062 vdd.n1270 vdd.n1269 185
R1063 vdd.n1305 vdd.n1269 185
R1064 vdd.n1501 vdd.n1500 185
R1065 vdd.n1273 vdd.n1272 185
R1066 vdd.n1497 vdd.n1496 185
R1067 vdd.n1498 vdd.n1497 185
R1068 vdd.n1307 vdd.n1306 185
R1069 vdd.n1492 vdd.n1309 185
R1070 vdd.n1491 vdd.n1310 185
R1071 vdd.n1490 vdd.n1311 185
R1072 vdd.n1313 vdd.n1312 185
R1073 vdd.n1486 vdd.n1315 185
R1074 vdd.n1485 vdd.n1316 185
R1075 vdd.n1484 vdd.n1317 185
R1076 vdd.n1319 vdd.n1318 185
R1077 vdd.n1480 vdd.n1321 185
R1078 vdd.n1479 vdd.n1322 185
R1079 vdd.n1478 vdd.n1323 185
R1080 vdd.n1325 vdd.n1324 185
R1081 vdd.n1474 vdd.n1327 185
R1082 vdd.n1473 vdd.n1328 185
R1083 vdd.n1472 vdd.n1329 185
R1084 vdd.n1333 vdd.n1330 185
R1085 vdd.n1468 vdd.n1335 185
R1086 vdd.n1467 vdd.n1336 185
R1087 vdd.n1466 vdd.n1337 185
R1088 vdd.n1339 vdd.n1338 185
R1089 vdd.n1462 vdd.n1341 185
R1090 vdd.n1461 vdd.n1342 185
R1091 vdd.n1460 vdd.n1343 185
R1092 vdd.n1345 vdd.n1344 185
R1093 vdd.n1456 vdd.n1347 185
R1094 vdd.n1455 vdd.n1348 185
R1095 vdd.n1454 vdd.n1349 185
R1096 vdd.n1351 vdd.n1350 185
R1097 vdd.n1450 vdd.n1353 185
R1098 vdd.n1449 vdd.n1354 185
R1099 vdd.n1448 vdd.n1355 185
R1100 vdd.n1357 vdd.n1356 185
R1101 vdd.n1444 vdd.n1359 185
R1102 vdd.n1443 vdd.n1360 185
R1103 vdd.n1442 vdd.n1361 185
R1104 vdd.n1363 vdd.n1362 185
R1105 vdd.n1438 vdd.n1365 185
R1106 vdd.n1437 vdd.n1434 185
R1107 vdd.n1433 vdd.n1366 185
R1108 vdd.n1368 vdd.n1367 185
R1109 vdd.n1429 vdd.n1370 185
R1110 vdd.n1428 vdd.n1371 185
R1111 vdd.n1427 vdd.n1372 185
R1112 vdd.n1374 vdd.n1373 185
R1113 vdd.n1423 vdd.n1376 185
R1114 vdd.n1422 vdd.n1377 185
R1115 vdd.n1421 vdd.n1378 185
R1116 vdd.n1380 vdd.n1379 185
R1117 vdd.n1417 vdd.n1382 185
R1118 vdd.n1416 vdd.n1383 185
R1119 vdd.n1415 vdd.n1384 185
R1120 vdd.n1386 vdd.n1385 185
R1121 vdd.n1411 vdd.n1388 185
R1122 vdd.n1410 vdd.n1389 185
R1123 vdd.n1409 vdd.n1390 185
R1124 vdd.n1392 vdd.n1391 185
R1125 vdd.n1405 vdd.n1394 185
R1126 vdd.n1404 vdd.n1395 185
R1127 vdd.n1403 vdd.n1396 185
R1128 vdd.n1400 vdd.n1304 185
R1129 vdd.n1498 vdd.n1304 185
R1130 vdd.n2199 vdd.n2198 185
R1131 vdd.n2203 vdd.n1149 185
R1132 vdd.n2079 vdd.n1148 185
R1133 vdd.n2082 vdd.n2081 185
R1134 vdd.n2084 vdd.n2083 185
R1135 vdd.n2087 vdd.n2086 185
R1136 vdd.n2089 vdd.n2088 185
R1137 vdd.n2091 vdd.n2077 185
R1138 vdd.n2093 vdd.n2092 185
R1139 vdd.n2094 vdd.n2071 185
R1140 vdd.n2096 vdd.n2095 185
R1141 vdd.n2098 vdd.n2069 185
R1142 vdd.n2100 vdd.n2099 185
R1143 vdd.n2101 vdd.n2064 185
R1144 vdd.n2103 vdd.n2102 185
R1145 vdd.n2105 vdd.n2062 185
R1146 vdd.n2107 vdd.n2106 185
R1147 vdd.n2108 vdd.n2058 185
R1148 vdd.n2110 vdd.n2109 185
R1149 vdd.n2112 vdd.n2055 185
R1150 vdd.n2114 vdd.n2113 185
R1151 vdd.n2056 vdd.n2049 185
R1152 vdd.n2118 vdd.n2053 185
R1153 vdd.n2119 vdd.n2045 185
R1154 vdd.n2121 vdd.n2120 185
R1155 vdd.n2123 vdd.n2043 185
R1156 vdd.n2125 vdd.n2124 185
R1157 vdd.n2126 vdd.n2038 185
R1158 vdd.n2128 vdd.n2127 185
R1159 vdd.n2130 vdd.n2036 185
R1160 vdd.n2132 vdd.n2131 185
R1161 vdd.n2133 vdd.n2031 185
R1162 vdd.n2135 vdd.n2134 185
R1163 vdd.n2137 vdd.n2029 185
R1164 vdd.n2139 vdd.n2138 185
R1165 vdd.n2140 vdd.n2024 185
R1166 vdd.n2142 vdd.n2141 185
R1167 vdd.n2144 vdd.n2022 185
R1168 vdd.n2146 vdd.n2145 185
R1169 vdd.n2147 vdd.n2018 185
R1170 vdd.n2149 vdd.n2148 185
R1171 vdd.n2151 vdd.n2015 185
R1172 vdd.n2153 vdd.n2152 185
R1173 vdd.n2016 vdd.n2009 185
R1174 vdd.n2157 vdd.n2013 185
R1175 vdd.n2158 vdd.n2005 185
R1176 vdd.n2160 vdd.n2159 185
R1177 vdd.n2162 vdd.n2003 185
R1178 vdd.n2164 vdd.n2163 185
R1179 vdd.n2165 vdd.n1998 185
R1180 vdd.n2167 vdd.n2166 185
R1181 vdd.n2169 vdd.n1996 185
R1182 vdd.n2171 vdd.n2170 185
R1183 vdd.n2172 vdd.n1991 185
R1184 vdd.n2174 vdd.n2173 185
R1185 vdd.n2176 vdd.n1990 185
R1186 vdd.n2177 vdd.n1987 185
R1187 vdd.n2180 vdd.n2179 185
R1188 vdd.n1989 vdd.n1985 185
R1189 vdd.n2184 vdd.n1983 185
R1190 vdd.n2186 vdd.n2185 185
R1191 vdd.n2188 vdd.n1981 185
R1192 vdd.n2190 vdd.n2189 185
R1193 vdd.n2191 vdd.n1155 185
R1194 vdd.n2197 vdd.n1152 185
R1195 vdd.n2197 vdd.n2196 185
R1196 vdd.n1163 vdd.n1151 185
R1197 vdd.n1974 vdd.n1151 185
R1198 vdd.n1973 vdd.n1972 185
R1199 vdd.n1975 vdd.n1973 185
R1200 vdd.n1162 vdd.n1161 185
R1201 vdd.n1161 vdd.n1160 185
R1202 vdd.n1966 vdd.n1965 185
R1203 vdd.n1965 vdd.n1964 185
R1204 vdd.n1166 vdd.n1165 185
R1205 vdd.n1955 vdd.n1166 185
R1206 vdd.n1954 vdd.n1953 185
R1207 vdd.n1956 vdd.n1954 185
R1208 vdd.n1173 vdd.n1172 185
R1209 vdd.n1178 vdd.n1172 185
R1210 vdd.n1949 vdd.n1948 185
R1211 vdd.n1948 vdd.n1947 185
R1212 vdd.n1176 vdd.n1175 185
R1213 vdd.n1177 vdd.n1176 185
R1214 vdd.n1938 vdd.n1937 185
R1215 vdd.n1939 vdd.n1938 185
R1216 vdd.n1186 vdd.n1185 185
R1217 vdd.n1185 vdd.n1184 185
R1218 vdd.n1933 vdd.n1932 185
R1219 vdd.n1932 vdd.n1931 185
R1220 vdd.n1189 vdd.n1188 185
R1221 vdd.n1922 vdd.n1189 185
R1222 vdd.n1921 vdd.n1920 185
R1223 vdd.n1923 vdd.n1921 185
R1224 vdd.n1196 vdd.n1195 185
R1225 vdd.n1200 vdd.n1195 185
R1226 vdd.n1916 vdd.n1915 185
R1227 vdd.n1915 vdd.n1914 185
R1228 vdd.n1199 vdd.n1198 185
R1229 vdd.n1905 vdd.n1199 185
R1230 vdd.n1904 vdd.n1903 185
R1231 vdd.n1906 vdd.n1904 185
R1232 vdd.n1208 vdd.n1207 185
R1233 vdd.n1207 vdd.n1206 185
R1234 vdd.n1899 vdd.n1898 185
R1235 vdd.n1898 vdd.n1897 185
R1236 vdd.n1211 vdd.n1210 185
R1237 vdd.n1212 vdd.n1211 185
R1238 vdd.n1581 vdd.n1580 185
R1239 vdd.n1582 vdd.n1581 185
R1240 vdd.n1219 vdd.n1218 185
R1241 vdd.n1223 vdd.n1218 185
R1242 vdd.n1576 vdd.n1575 185
R1243 vdd.n1575 vdd.n1574 185
R1244 vdd.n1222 vdd.n1221 185
R1245 vdd.n1565 vdd.n1222 185
R1246 vdd.n1564 vdd.n1563 185
R1247 vdd.n1566 vdd.n1564 185
R1248 vdd.n1230 vdd.n1229 185
R1249 vdd.n1235 vdd.n1229 185
R1250 vdd.n1559 vdd.n1558 185
R1251 vdd.n1558 vdd.n1557 185
R1252 vdd.n1233 vdd.n1232 185
R1253 vdd.n1234 vdd.n1233 185
R1254 vdd.n1548 vdd.n1547 185
R1255 vdd.n1549 vdd.n1548 185
R1256 vdd.n1243 vdd.n1242 185
R1257 vdd.n1242 vdd.n1241 185
R1258 vdd.n1543 vdd.n1542 185
R1259 vdd.n1542 vdd.n1541 185
R1260 vdd.n1246 vdd.n1245 185
R1261 vdd.n1532 vdd.n1246 185
R1262 vdd.n1531 vdd.n1530 185
R1263 vdd.n1533 vdd.n1531 185
R1264 vdd.n1253 vdd.n1252 185
R1265 vdd.n1257 vdd.n1252 185
R1266 vdd.n1526 vdd.n1525 185
R1267 vdd.n1525 vdd.n1524 185
R1268 vdd.n1256 vdd.n1255 185
R1269 vdd.n1515 vdd.n1256 185
R1270 vdd.n1514 vdd.n1513 185
R1271 vdd.n1516 vdd.n1514 185
R1272 vdd.n1265 vdd.n1264 185
R1273 vdd.n1264 vdd.n1263 185
R1274 vdd.n1509 vdd.n1508 185
R1275 vdd.n1508 vdd.n1507 185
R1276 vdd.n1268 vdd.n1267 185
R1277 vdd.n1305 vdd.n1268 185
R1278 vdd.n987 vdd.n985 185
R1279 vdd.n2654 vdd.n985 185
R1280 vdd.n2576 vdd.n1005 185
R1281 vdd.n1005 vdd.n992 185
R1282 vdd.n2578 vdd.n2577 185
R1283 vdd.n2579 vdd.n2578 185
R1284 vdd.n2575 vdd.n1004 185
R1285 vdd.n2334 vdd.n1004 185
R1286 vdd.n2574 vdd.n2573 185
R1287 vdd.n2573 vdd.n2572 185
R1288 vdd.n1007 vdd.n1006 185
R1289 vdd.n1008 vdd.n1007 185
R1290 vdd.n2563 vdd.n2562 185
R1291 vdd.n2564 vdd.n2563 185
R1292 vdd.n2561 vdd.n1018 185
R1293 vdd.n1018 vdd.n1015 185
R1294 vdd.n2560 vdd.n2559 185
R1295 vdd.n2559 vdd.n2558 185
R1296 vdd.n1020 vdd.n1019 185
R1297 vdd.n2346 vdd.n1020 185
R1298 vdd.n2551 vdd.n2550 185
R1299 vdd.n2552 vdd.n2551 185
R1300 vdd.n2549 vdd.n1028 185
R1301 vdd.n1033 vdd.n1028 185
R1302 vdd.n2548 vdd.n2547 185
R1303 vdd.n2547 vdd.n2546 185
R1304 vdd.n1030 vdd.n1029 185
R1305 vdd.n1039 vdd.n1030 185
R1306 vdd.n2539 vdd.n2538 185
R1307 vdd.n2540 vdd.n2539 185
R1308 vdd.n2537 vdd.n1040 185
R1309 vdd.n2358 vdd.n1040 185
R1310 vdd.n2536 vdd.n2535 185
R1311 vdd.n2535 vdd.n2534 185
R1312 vdd.n1042 vdd.n1041 185
R1313 vdd.n1043 vdd.n1042 185
R1314 vdd.n2527 vdd.n2526 185
R1315 vdd.n2528 vdd.n2527 185
R1316 vdd.n2525 vdd.n1052 185
R1317 vdd.n1052 vdd.n1049 185
R1318 vdd.n2524 vdd.n2523 185
R1319 vdd.n2523 vdd.n2522 185
R1320 vdd.n1054 vdd.n1053 185
R1321 vdd.n1063 vdd.n1054 185
R1322 vdd.n2514 vdd.n2513 185
R1323 vdd.n2515 vdd.n2514 185
R1324 vdd.n2512 vdd.n1064 185
R1325 vdd.n1070 vdd.n1064 185
R1326 vdd.n2511 vdd.n2510 185
R1327 vdd.n2510 vdd.n2509 185
R1328 vdd.n1066 vdd.n1065 185
R1329 vdd.n1067 vdd.n1066 185
R1330 vdd.n2502 vdd.n2501 185
R1331 vdd.n2503 vdd.n2502 185
R1332 vdd.n2500 vdd.n1077 185
R1333 vdd.n1077 vdd.n1074 185
R1334 vdd.n2499 vdd.n2498 185
R1335 vdd.n2498 vdd.n2497 185
R1336 vdd.n1079 vdd.n1078 185
R1337 vdd.n1080 vdd.n1079 185
R1338 vdd.n2490 vdd.n2489 185
R1339 vdd.n2491 vdd.n2490 185
R1340 vdd.n2488 vdd.n1089 185
R1341 vdd.n1089 vdd.n1086 185
R1342 vdd.n2487 vdd.n2486 185
R1343 vdd.n2486 vdd.n2485 185
R1344 vdd.n1091 vdd.n1090 185
R1345 vdd.n1092 vdd.n1091 185
R1346 vdd.n2478 vdd.n2477 185
R1347 vdd.n2479 vdd.n2478 185
R1348 vdd.n2476 vdd.n1101 185
R1349 vdd.n1101 vdd.n1098 185
R1350 vdd.n2475 vdd.n2474 185
R1351 vdd.n2474 vdd.n2473 185
R1352 vdd.n1103 vdd.n1102 185
R1353 vdd.n1104 vdd.n1103 185
R1354 vdd.n2466 vdd.n2465 185
R1355 vdd.n2467 vdd.n2466 185
R1356 vdd.n2464 vdd.n1113 185
R1357 vdd.n2463 vdd.n2462 185
R1358 vdd.n2460 vdd.n1114 185
R1359 vdd.n2460 vdd.n1110 185
R1360 vdd.n2459 vdd.n2458 185
R1361 vdd.n2457 vdd.n2456 185
R1362 vdd.n2455 vdd.n1116 185
R1363 vdd.n2453 vdd.n2452 185
R1364 vdd.n2451 vdd.n1117 185
R1365 vdd.n2450 vdd.n2449 185
R1366 vdd.n2447 vdd.n1118 185
R1367 vdd.n2445 vdd.n2444 185
R1368 vdd.n2443 vdd.n1119 185
R1369 vdd.n2442 vdd.n2441 185
R1370 vdd.n2439 vdd.n1120 185
R1371 vdd.n2437 vdd.n2436 185
R1372 vdd.n2435 vdd.n1121 185
R1373 vdd.n2434 vdd.n2433 185
R1374 vdd.n2431 vdd.n1122 185
R1375 vdd.n2429 vdd.n2428 185
R1376 vdd.n2427 vdd.n1123 185
R1377 vdd.n2426 vdd.n2425 185
R1378 vdd.n2423 vdd.n1124 185
R1379 vdd.n2421 vdd.n2420 185
R1380 vdd.n2419 vdd.n1125 185
R1381 vdd.n2418 vdd.n2417 185
R1382 vdd.n2415 vdd.n1126 185
R1383 vdd.n2413 vdd.n2412 185
R1384 vdd.n2411 vdd.n1127 185
R1385 vdd.n2410 vdd.n2409 185
R1386 vdd.n2407 vdd.n1128 185
R1387 vdd.n2405 vdd.n2404 185
R1388 vdd.n2403 vdd.n1129 185
R1389 vdd.n2401 vdd.n2400 185
R1390 vdd.n2398 vdd.n1132 185
R1391 vdd.n2396 vdd.n2395 185
R1392 vdd.n2657 vdd.n2656 185
R1393 vdd.n2659 vdd.n2658 185
R1394 vdd.n2661 vdd.n2660 185
R1395 vdd.n2664 vdd.n2663 185
R1396 vdd.n2666 vdd.n2665 185
R1397 vdd.n2668 vdd.n2667 185
R1398 vdd.n2670 vdd.n2669 185
R1399 vdd.n2672 vdd.n2671 185
R1400 vdd.n2674 vdd.n2673 185
R1401 vdd.n2676 vdd.n2675 185
R1402 vdd.n2678 vdd.n2677 185
R1403 vdd.n2680 vdd.n2679 185
R1404 vdd.n2682 vdd.n2681 185
R1405 vdd.n2684 vdd.n2683 185
R1406 vdd.n2686 vdd.n2685 185
R1407 vdd.n2688 vdd.n2687 185
R1408 vdd.n2690 vdd.n2689 185
R1409 vdd.n2692 vdd.n2691 185
R1410 vdd.n2694 vdd.n2693 185
R1411 vdd.n2696 vdd.n2695 185
R1412 vdd.n2698 vdd.n2697 185
R1413 vdd.n2700 vdd.n2699 185
R1414 vdd.n2702 vdd.n2701 185
R1415 vdd.n2704 vdd.n2703 185
R1416 vdd.n2706 vdd.n2705 185
R1417 vdd.n2708 vdd.n2707 185
R1418 vdd.n2710 vdd.n2709 185
R1419 vdd.n2712 vdd.n2711 185
R1420 vdd.n2714 vdd.n2713 185
R1421 vdd.n2716 vdd.n2715 185
R1422 vdd.n2718 vdd.n2717 185
R1423 vdd.n2720 vdd.n2719 185
R1424 vdd.n2722 vdd.n2721 185
R1425 vdd.n2723 vdd.n986 185
R1426 vdd.n2725 vdd.n2724 185
R1427 vdd.n2726 vdd.n2725 185
R1428 vdd.n2655 vdd.n990 185
R1429 vdd.n2655 vdd.n2654 185
R1430 vdd.n2332 vdd.n991 185
R1431 vdd.n992 vdd.n991 185
R1432 vdd.n2333 vdd.n1002 185
R1433 vdd.n2579 vdd.n1002 185
R1434 vdd.n2336 vdd.n2335 185
R1435 vdd.n2335 vdd.n2334 185
R1436 vdd.n2337 vdd.n1009 185
R1437 vdd.n2572 vdd.n1009 185
R1438 vdd.n2339 vdd.n2338 185
R1439 vdd.n2338 vdd.n1008 185
R1440 vdd.n2340 vdd.n1016 185
R1441 vdd.n2564 vdd.n1016 185
R1442 vdd.n2342 vdd.n2341 185
R1443 vdd.n2341 vdd.n1015 185
R1444 vdd.n2343 vdd.n1021 185
R1445 vdd.n2558 vdd.n1021 185
R1446 vdd.n2345 vdd.n2344 185
R1447 vdd.n2346 vdd.n2345 185
R1448 vdd.n2331 vdd.n1026 185
R1449 vdd.n2552 vdd.n1026 185
R1450 vdd.n2330 vdd.n2329 185
R1451 vdd.n2329 vdd.n1033 185
R1452 vdd.n2328 vdd.n1031 185
R1453 vdd.n2546 vdd.n1031 185
R1454 vdd.n2327 vdd.n2326 185
R1455 vdd.n2326 vdd.n1039 185
R1456 vdd.n1133 vdd.n1037 185
R1457 vdd.n2540 vdd.n1037 185
R1458 vdd.n2360 vdd.n2359 185
R1459 vdd.n2359 vdd.n2358 185
R1460 vdd.n2361 vdd.n1044 185
R1461 vdd.n2534 vdd.n1044 185
R1462 vdd.n2363 vdd.n2362 185
R1463 vdd.n2362 vdd.n1043 185
R1464 vdd.n2364 vdd.n1050 185
R1465 vdd.n2528 vdd.n1050 185
R1466 vdd.n2366 vdd.n2365 185
R1467 vdd.n2365 vdd.n1049 185
R1468 vdd.n2367 vdd.n1055 185
R1469 vdd.n2522 vdd.n1055 185
R1470 vdd.n2369 vdd.n2368 185
R1471 vdd.n2368 vdd.n1063 185
R1472 vdd.n2370 vdd.n1061 185
R1473 vdd.n2515 vdd.n1061 185
R1474 vdd.n2372 vdd.n2371 185
R1475 vdd.n2371 vdd.n1070 185
R1476 vdd.n2373 vdd.n1068 185
R1477 vdd.n2509 vdd.n1068 185
R1478 vdd.n2375 vdd.n2374 185
R1479 vdd.n2374 vdd.n1067 185
R1480 vdd.n2376 vdd.n1075 185
R1481 vdd.n2503 vdd.n1075 185
R1482 vdd.n2378 vdd.n2377 185
R1483 vdd.n2377 vdd.n1074 185
R1484 vdd.n2379 vdd.n1081 185
R1485 vdd.n2497 vdd.n1081 185
R1486 vdd.n2381 vdd.n2380 185
R1487 vdd.n2380 vdd.n1080 185
R1488 vdd.n2382 vdd.n1087 185
R1489 vdd.n2491 vdd.n1087 185
R1490 vdd.n2384 vdd.n2383 185
R1491 vdd.n2383 vdd.n1086 185
R1492 vdd.n2385 vdd.n1093 185
R1493 vdd.n2485 vdd.n1093 185
R1494 vdd.n2387 vdd.n2386 185
R1495 vdd.n2386 vdd.n1092 185
R1496 vdd.n2388 vdd.n1099 185
R1497 vdd.n2479 vdd.n1099 185
R1498 vdd.n2390 vdd.n2389 185
R1499 vdd.n2389 vdd.n1098 185
R1500 vdd.n2391 vdd.n1105 185
R1501 vdd.n2473 vdd.n1105 185
R1502 vdd.n2393 vdd.n2392 185
R1503 vdd.n2392 vdd.n1104 185
R1504 vdd.n2394 vdd.n1111 185
R1505 vdd.n2467 vdd.n1111 185
R1506 vdd.n3539 vdd.n3538 185
R1507 vdd.n3538 vdd.n3537 185
R1508 vdd.n3540 vdd.n387 185
R1509 vdd.n387 vdd.n386 185
R1510 vdd.n3542 vdd.n3541 185
R1511 vdd.n3543 vdd.n3542 185
R1512 vdd.n382 vdd.n381 185
R1513 vdd.n3544 vdd.n382 185
R1514 vdd.n3547 vdd.n3546 185
R1515 vdd.n3546 vdd.n3545 185
R1516 vdd.n3548 vdd.n376 185
R1517 vdd.n376 vdd.n375 185
R1518 vdd.n3550 vdd.n3549 185
R1519 vdd.n3551 vdd.n3550 185
R1520 vdd.n371 vdd.n370 185
R1521 vdd.n3552 vdd.n371 185
R1522 vdd.n3555 vdd.n3554 185
R1523 vdd.n3554 vdd.n3553 185
R1524 vdd.n3556 vdd.n365 185
R1525 vdd.n3513 vdd.n365 185
R1526 vdd.n3558 vdd.n3557 185
R1527 vdd.n3559 vdd.n3558 185
R1528 vdd.n360 vdd.n359 185
R1529 vdd.n3560 vdd.n360 185
R1530 vdd.n3563 vdd.n3562 185
R1531 vdd.n3562 vdd.n3561 185
R1532 vdd.n3564 vdd.n354 185
R1533 vdd.n361 vdd.n354 185
R1534 vdd.n3566 vdd.n3565 185
R1535 vdd.n3567 vdd.n3566 185
R1536 vdd.n350 vdd.n349 185
R1537 vdd.n3568 vdd.n350 185
R1538 vdd.n3571 vdd.n3570 185
R1539 vdd.n3570 vdd.n3569 185
R1540 vdd.n3572 vdd.n345 185
R1541 vdd.n345 vdd.n344 185
R1542 vdd.n3574 vdd.n3573 185
R1543 vdd.n3575 vdd.n3574 185
R1544 vdd.n339 vdd.n337 185
R1545 vdd.n3576 vdd.n339 185
R1546 vdd.n3579 vdd.n3578 185
R1547 vdd.n3578 vdd.n3577 185
R1548 vdd.n338 vdd.n336 185
R1549 vdd.n340 vdd.n338 185
R1550 vdd.n3489 vdd.n3488 185
R1551 vdd.n3490 vdd.n3489 185
R1552 vdd.n635 vdd.n634 185
R1553 vdd.n634 vdd.n633 185
R1554 vdd.n3484 vdd.n3483 185
R1555 vdd.n3483 vdd.n3482 185
R1556 vdd.n638 vdd.n637 185
R1557 vdd.n644 vdd.n638 185
R1558 vdd.n3470 vdd.n3469 185
R1559 vdd.n3471 vdd.n3470 185
R1560 vdd.n646 vdd.n645 185
R1561 vdd.n3462 vdd.n645 185
R1562 vdd.n3465 vdd.n3464 185
R1563 vdd.n3464 vdd.n3463 185
R1564 vdd.n649 vdd.n648 185
R1565 vdd.n656 vdd.n649 185
R1566 vdd.n3453 vdd.n3452 185
R1567 vdd.n3454 vdd.n3453 185
R1568 vdd.n658 vdd.n657 185
R1569 vdd.n657 vdd.n655 185
R1570 vdd.n3448 vdd.n3447 185
R1571 vdd.n3447 vdd.n3446 185
R1572 vdd.n661 vdd.n660 185
R1573 vdd.n662 vdd.n661 185
R1574 vdd.n3437 vdd.n3436 185
R1575 vdd.n3438 vdd.n3437 185
R1576 vdd.n669 vdd.n668 185
R1577 vdd.n3429 vdd.n668 185
R1578 vdd.n3432 vdd.n3431 185
R1579 vdd.n3431 vdd.n3430 185
R1580 vdd.n672 vdd.n671 185
R1581 vdd.n679 vdd.n672 185
R1582 vdd.n3420 vdd.n3419 185
R1583 vdd.n3421 vdd.n3420 185
R1584 vdd.n681 vdd.n680 185
R1585 vdd.n680 vdd.n678 185
R1586 vdd.n3415 vdd.n3414 185
R1587 vdd.n3414 vdd.n3413 185
R1588 vdd.n684 vdd.n683 185
R1589 vdd.n723 vdd.n684 185
R1590 vdd.n3403 vdd.n3402 185
R1591 vdd.n3401 vdd.n725 185
R1592 vdd.n3400 vdd.n724 185
R1593 vdd.n3405 vdd.n724 185
R1594 vdd.n729 vdd.n728 185
R1595 vdd.n733 vdd.n732 185
R1596 vdd.n3396 vdd.n734 185
R1597 vdd.n3395 vdd.n3394 185
R1598 vdd.n3393 vdd.n3392 185
R1599 vdd.n3391 vdd.n3390 185
R1600 vdd.n3389 vdd.n3388 185
R1601 vdd.n3387 vdd.n3386 185
R1602 vdd.n3385 vdd.n3384 185
R1603 vdd.n3383 vdd.n3382 185
R1604 vdd.n3381 vdd.n3380 185
R1605 vdd.n3379 vdd.n3378 185
R1606 vdd.n3377 vdd.n3376 185
R1607 vdd.n3375 vdd.n3374 185
R1608 vdd.n3373 vdd.n3372 185
R1609 vdd.n3371 vdd.n3370 185
R1610 vdd.n3369 vdd.n3368 185
R1611 vdd.n3360 vdd.n747 185
R1612 vdd.n3362 vdd.n3361 185
R1613 vdd.n3359 vdd.n3358 185
R1614 vdd.n3357 vdd.n3356 185
R1615 vdd.n3355 vdd.n3354 185
R1616 vdd.n3353 vdd.n3352 185
R1617 vdd.n3351 vdd.n3350 185
R1618 vdd.n3349 vdd.n3348 185
R1619 vdd.n3347 vdd.n3346 185
R1620 vdd.n3345 vdd.n3344 185
R1621 vdd.n3343 vdd.n3342 185
R1622 vdd.n3341 vdd.n3340 185
R1623 vdd.n3339 vdd.n3338 185
R1624 vdd.n3337 vdd.n3336 185
R1625 vdd.n3335 vdd.n3334 185
R1626 vdd.n3333 vdd.n3332 185
R1627 vdd.n3331 vdd.n3330 185
R1628 vdd.n3329 vdd.n3328 185
R1629 vdd.n3327 vdd.n3326 185
R1630 vdd.n3325 vdd.n3324 185
R1631 vdd.n3323 vdd.n3322 185
R1632 vdd.n3321 vdd.n3320 185
R1633 vdd.n3314 vdd.n767 185
R1634 vdd.n3316 vdd.n3315 185
R1635 vdd.n3313 vdd.n3312 185
R1636 vdd.n3311 vdd.n3310 185
R1637 vdd.n3309 vdd.n3308 185
R1638 vdd.n3307 vdd.n3306 185
R1639 vdd.n3305 vdd.n3304 185
R1640 vdd.n3303 vdd.n3302 185
R1641 vdd.n3301 vdd.n3300 185
R1642 vdd.n3299 vdd.n3298 185
R1643 vdd.n3297 vdd.n3296 185
R1644 vdd.n3295 vdd.n3294 185
R1645 vdd.n3293 vdd.n3292 185
R1646 vdd.n3291 vdd.n3290 185
R1647 vdd.n3289 vdd.n3288 185
R1648 vdd.n3287 vdd.n3286 185
R1649 vdd.n3285 vdd.n3284 185
R1650 vdd.n3283 vdd.n3282 185
R1651 vdd.n3281 vdd.n3280 185
R1652 vdd.n3279 vdd.n3278 185
R1653 vdd.n3277 vdd.n691 185
R1654 vdd.n3407 vdd.n3406 185
R1655 vdd.n3406 vdd.n3405 185
R1656 vdd.n3534 vdd.n3533 185
R1657 vdd.n618 vdd.n425 185
R1658 vdd.n617 vdd.n616 185
R1659 vdd.n615 vdd.n614 185
R1660 vdd.n613 vdd.n430 185
R1661 vdd.n609 vdd.n608 185
R1662 vdd.n607 vdd.n606 185
R1663 vdd.n605 vdd.n604 185
R1664 vdd.n603 vdd.n432 185
R1665 vdd.n599 vdd.n598 185
R1666 vdd.n597 vdd.n596 185
R1667 vdd.n595 vdd.n594 185
R1668 vdd.n593 vdd.n434 185
R1669 vdd.n589 vdd.n588 185
R1670 vdd.n587 vdd.n586 185
R1671 vdd.n585 vdd.n584 185
R1672 vdd.n583 vdd.n436 185
R1673 vdd.n579 vdd.n578 185
R1674 vdd.n577 vdd.n576 185
R1675 vdd.n575 vdd.n574 185
R1676 vdd.n573 vdd.n438 185
R1677 vdd.n569 vdd.n568 185
R1678 vdd.n567 vdd.n566 185
R1679 vdd.n565 vdd.n564 185
R1680 vdd.n563 vdd.n442 185
R1681 vdd.n559 vdd.n558 185
R1682 vdd.n557 vdd.n556 185
R1683 vdd.n555 vdd.n554 185
R1684 vdd.n553 vdd.n444 185
R1685 vdd.n549 vdd.n548 185
R1686 vdd.n547 vdd.n546 185
R1687 vdd.n545 vdd.n544 185
R1688 vdd.n543 vdd.n446 185
R1689 vdd.n539 vdd.n538 185
R1690 vdd.n537 vdd.n536 185
R1691 vdd.n535 vdd.n534 185
R1692 vdd.n533 vdd.n448 185
R1693 vdd.n529 vdd.n528 185
R1694 vdd.n527 vdd.n526 185
R1695 vdd.n525 vdd.n524 185
R1696 vdd.n523 vdd.n450 185
R1697 vdd.n519 vdd.n518 185
R1698 vdd.n517 vdd.n516 185
R1699 vdd.n515 vdd.n514 185
R1700 vdd.n513 vdd.n454 185
R1701 vdd.n509 vdd.n508 185
R1702 vdd.n507 vdd.n506 185
R1703 vdd.n505 vdd.n504 185
R1704 vdd.n503 vdd.n456 185
R1705 vdd.n499 vdd.n498 185
R1706 vdd.n497 vdd.n496 185
R1707 vdd.n495 vdd.n494 185
R1708 vdd.n493 vdd.n458 185
R1709 vdd.n489 vdd.n488 185
R1710 vdd.n487 vdd.n486 185
R1711 vdd.n485 vdd.n484 185
R1712 vdd.n483 vdd.n460 185
R1713 vdd.n479 vdd.n478 185
R1714 vdd.n477 vdd.n476 185
R1715 vdd.n475 vdd.n474 185
R1716 vdd.n473 vdd.n462 185
R1717 vdd.n469 vdd.n468 185
R1718 vdd.n467 vdd.n466 185
R1719 vdd.n465 vdd.n392 185
R1720 vdd.n3530 vdd.n393 185
R1721 vdd.n3537 vdd.n393 185
R1722 vdd.n3529 vdd.n3528 185
R1723 vdd.n3528 vdd.n386 185
R1724 vdd.n3527 vdd.n385 185
R1725 vdd.n3543 vdd.n385 185
R1726 vdd.n621 vdd.n384 185
R1727 vdd.n3544 vdd.n384 185
R1728 vdd.n3523 vdd.n383 185
R1729 vdd.n3545 vdd.n383 185
R1730 vdd.n3522 vdd.n3521 185
R1731 vdd.n3521 vdd.n375 185
R1732 vdd.n3520 vdd.n374 185
R1733 vdd.n3551 vdd.n374 185
R1734 vdd.n623 vdd.n373 185
R1735 vdd.n3552 vdd.n373 185
R1736 vdd.n3516 vdd.n372 185
R1737 vdd.n3553 vdd.n372 185
R1738 vdd.n3515 vdd.n3514 185
R1739 vdd.n3514 vdd.n3513 185
R1740 vdd.n3512 vdd.n364 185
R1741 vdd.n3559 vdd.n364 185
R1742 vdd.n625 vdd.n363 185
R1743 vdd.n3560 vdd.n363 185
R1744 vdd.n3508 vdd.n362 185
R1745 vdd.n3561 vdd.n362 185
R1746 vdd.n3507 vdd.n3506 185
R1747 vdd.n3506 vdd.n361 185
R1748 vdd.n3505 vdd.n353 185
R1749 vdd.n3567 vdd.n353 185
R1750 vdd.n627 vdd.n352 185
R1751 vdd.n3568 vdd.n352 185
R1752 vdd.n3501 vdd.n351 185
R1753 vdd.n3569 vdd.n351 185
R1754 vdd.n3500 vdd.n3499 185
R1755 vdd.n3499 vdd.n344 185
R1756 vdd.n3498 vdd.n343 185
R1757 vdd.n3575 vdd.n343 185
R1758 vdd.n629 vdd.n342 185
R1759 vdd.n3576 vdd.n342 185
R1760 vdd.n3494 vdd.n341 185
R1761 vdd.n3577 vdd.n341 185
R1762 vdd.n3493 vdd.n3492 185
R1763 vdd.n3492 vdd.n340 185
R1764 vdd.n3491 vdd.n631 185
R1765 vdd.n3491 vdd.n3490 185
R1766 vdd.n3479 vdd.n632 185
R1767 vdd.n633 vdd.n632 185
R1768 vdd.n3481 vdd.n3480 185
R1769 vdd.n3482 vdd.n3481 185
R1770 vdd.n640 vdd.n639 185
R1771 vdd.n644 vdd.n639 185
R1772 vdd.n3473 vdd.n3472 185
R1773 vdd.n3472 vdd.n3471 185
R1774 vdd.n643 vdd.n642 185
R1775 vdd.n3462 vdd.n643 185
R1776 vdd.n3461 vdd.n3460 185
R1777 vdd.n3463 vdd.n3461 185
R1778 vdd.n651 vdd.n650 185
R1779 vdd.n656 vdd.n650 185
R1780 vdd.n3456 vdd.n3455 185
R1781 vdd.n3455 vdd.n3454 185
R1782 vdd.n654 vdd.n653 185
R1783 vdd.n655 vdd.n654 185
R1784 vdd.n3445 vdd.n3444 185
R1785 vdd.n3446 vdd.n3445 185
R1786 vdd.n664 vdd.n663 185
R1787 vdd.n663 vdd.n662 185
R1788 vdd.n3440 vdd.n3439 185
R1789 vdd.n3439 vdd.n3438 185
R1790 vdd.n667 vdd.n666 185
R1791 vdd.n3429 vdd.n667 185
R1792 vdd.n3428 vdd.n3427 185
R1793 vdd.n3430 vdd.n3428 185
R1794 vdd.n674 vdd.n673 185
R1795 vdd.n679 vdd.n673 185
R1796 vdd.n3423 vdd.n3422 185
R1797 vdd.n3422 vdd.n3421 185
R1798 vdd.n677 vdd.n676 185
R1799 vdd.n678 vdd.n677 185
R1800 vdd.n3412 vdd.n3411 185
R1801 vdd.n3413 vdd.n3412 185
R1802 vdd.n686 vdd.n685 185
R1803 vdd.n723 vdd.n685 185
R1804 vdd.n3014 vdd.n947 185
R1805 vdd.n3013 vdd.n3012 185
R1806 vdd.n949 vdd.n948 185
R1807 vdd.n3010 vdd.n949 185
R1808 vdd.n2833 vdd.n2832 185
R1809 vdd.n2835 vdd.n2834 185
R1810 vdd.n2837 vdd.n2836 185
R1811 vdd.n2839 vdd.n2838 185
R1812 vdd.n2841 vdd.n2840 185
R1813 vdd.n2843 vdd.n2842 185
R1814 vdd.n2845 vdd.n2844 185
R1815 vdd.n2847 vdd.n2846 185
R1816 vdd.n2849 vdd.n2848 185
R1817 vdd.n2851 vdd.n2850 185
R1818 vdd.n2853 vdd.n2852 185
R1819 vdd.n2855 vdd.n2854 185
R1820 vdd.n2857 vdd.n2856 185
R1821 vdd.n2859 vdd.n2858 185
R1822 vdd.n2861 vdd.n2860 185
R1823 vdd.n2863 vdd.n2862 185
R1824 vdd.n2865 vdd.n2864 185
R1825 vdd.n2867 vdd.n2866 185
R1826 vdd.n2869 vdd.n2868 185
R1827 vdd.n2871 vdd.n2870 185
R1828 vdd.n2873 vdd.n2872 185
R1829 vdd.n2875 vdd.n2874 185
R1830 vdd.n2877 vdd.n2876 185
R1831 vdd.n2879 vdd.n2878 185
R1832 vdd.n2881 vdd.n2880 185
R1833 vdd.n2883 vdd.n2882 185
R1834 vdd.n2885 vdd.n2884 185
R1835 vdd.n2887 vdd.n2886 185
R1836 vdd.n2889 vdd.n2888 185
R1837 vdd.n2892 vdd.n2891 185
R1838 vdd.n2894 vdd.n2893 185
R1839 vdd.n2896 vdd.n2895 185
R1840 vdd.n3177 vdd.n3176 185
R1841 vdd.n3179 vdd.n834 185
R1842 vdd.n3181 vdd.n3180 185
R1843 vdd.n3183 vdd.n831 185
R1844 vdd.n3185 vdd.n3184 185
R1845 vdd.n3187 vdd.n829 185
R1846 vdd.n3189 vdd.n3188 185
R1847 vdd.n3190 vdd.n828 185
R1848 vdd.n3192 vdd.n3191 185
R1849 vdd.n3194 vdd.n826 185
R1850 vdd.n3196 vdd.n3195 185
R1851 vdd.n3197 vdd.n825 185
R1852 vdd.n3199 vdd.n3198 185
R1853 vdd.n3201 vdd.n823 185
R1854 vdd.n3203 vdd.n3202 185
R1855 vdd.n3204 vdd.n822 185
R1856 vdd.n3206 vdd.n3205 185
R1857 vdd.n3208 vdd.n731 185
R1858 vdd.n3210 vdd.n3209 185
R1859 vdd.n3212 vdd.n820 185
R1860 vdd.n3214 vdd.n3213 185
R1861 vdd.n3215 vdd.n819 185
R1862 vdd.n3217 vdd.n3216 185
R1863 vdd.n3219 vdd.n817 185
R1864 vdd.n3221 vdd.n3220 185
R1865 vdd.n3222 vdd.n816 185
R1866 vdd.n3224 vdd.n3223 185
R1867 vdd.n3226 vdd.n814 185
R1868 vdd.n3228 vdd.n3227 185
R1869 vdd.n3229 vdd.n813 185
R1870 vdd.n3231 vdd.n3230 185
R1871 vdd.n3233 vdd.n812 185
R1872 vdd.n3234 vdd.n811 185
R1873 vdd.n3237 vdd.n3236 185
R1874 vdd.n3238 vdd.n809 185
R1875 vdd.n809 vdd.n692 185
R1876 vdd.n3175 vdd.n806 185
R1877 vdd.n3241 vdd.n806 185
R1878 vdd.n3174 vdd.n3173 185
R1879 vdd.n3173 vdd.n805 185
R1880 vdd.n3172 vdd.n836 185
R1881 vdd.n3172 vdd.n3171 185
R1882 vdd.n2946 vdd.n837 185
R1883 vdd.n846 vdd.n837 185
R1884 vdd.n2947 vdd.n844 185
R1885 vdd.n3165 vdd.n844 185
R1886 vdd.n2949 vdd.n2948 185
R1887 vdd.n2948 vdd.n843 185
R1888 vdd.n2950 vdd.n852 185
R1889 vdd.n3114 vdd.n852 185
R1890 vdd.n2952 vdd.n2951 185
R1891 vdd.n2951 vdd.n851 185
R1892 vdd.n2953 vdd.n857 185
R1893 vdd.n3108 vdd.n857 185
R1894 vdd.n2955 vdd.n2954 185
R1895 vdd.n2954 vdd.n864 185
R1896 vdd.n2956 vdd.n862 185
R1897 vdd.n3102 vdd.n862 185
R1898 vdd.n2958 vdd.n2957 185
R1899 vdd.n2957 vdd.n870 185
R1900 vdd.n2959 vdd.n868 185
R1901 vdd.n3096 vdd.n868 185
R1902 vdd.n2961 vdd.n2960 185
R1903 vdd.n2960 vdd.n877 185
R1904 vdd.n2962 vdd.n875 185
R1905 vdd.n3090 vdd.n875 185
R1906 vdd.n2964 vdd.n2963 185
R1907 vdd.n2963 vdd.n874 185
R1908 vdd.n2965 vdd.n882 185
R1909 vdd.n3084 vdd.n882 185
R1910 vdd.n2967 vdd.n2966 185
R1911 vdd.n2966 vdd.n881 185
R1912 vdd.n2968 vdd.n889 185
R1913 vdd.n3077 vdd.n889 185
R1914 vdd.n2970 vdd.n2969 185
R1915 vdd.n2969 vdd.n888 185
R1916 vdd.n2971 vdd.n894 185
R1917 vdd.n3071 vdd.n894 185
R1918 vdd.n2973 vdd.n2972 185
R1919 vdd.n2972 vdd.n901 185
R1920 vdd.n2974 vdd.n899 185
R1921 vdd.n3065 vdd.n899 185
R1922 vdd.n2976 vdd.n2975 185
R1923 vdd.n2977 vdd.n2976 185
R1924 vdd.n2945 vdd.n906 185
R1925 vdd.n3059 vdd.n906 185
R1926 vdd.n2944 vdd.n2943 185
R1927 vdd.n2943 vdd.n905 185
R1928 vdd.n2942 vdd.n912 185
R1929 vdd.n3053 vdd.n912 185
R1930 vdd.n2941 vdd.n2940 185
R1931 vdd.n2940 vdd.n911 185
R1932 vdd.n2901 vdd.n917 185
R1933 vdd.n3047 vdd.n917 185
R1934 vdd.n2991 vdd.n2990 185
R1935 vdd.n2990 vdd.n2989 185
R1936 vdd.n2992 vdd.n922 185
R1937 vdd.n3041 vdd.n922 185
R1938 vdd.n2994 vdd.n2993 185
R1939 vdd.n2993 vdd.n930 185
R1940 vdd.n2995 vdd.n928 185
R1941 vdd.n3035 vdd.n928 185
R1942 vdd.n2997 vdd.n2996 185
R1943 vdd.n2996 vdd.n927 185
R1944 vdd.n2998 vdd.n934 185
R1945 vdd.n3029 vdd.n934 185
R1946 vdd.n3000 vdd.n2999 185
R1947 vdd.n3001 vdd.n3000 185
R1948 vdd.n2900 vdd.n939 185
R1949 vdd.n3023 vdd.n939 185
R1950 vdd.n2899 vdd.n2898 185
R1951 vdd.n2898 vdd.n946 185
R1952 vdd.n2897 vdd.n944 185
R1953 vdd.n3017 vdd.n944 185
R1954 vdd.n3016 vdd.n3015 185
R1955 vdd.n3017 vdd.n3016 185
R1956 vdd.n938 vdd.n937 185
R1957 vdd.n946 vdd.n938 185
R1958 vdd.n3025 vdd.n3024 185
R1959 vdd.n3024 vdd.n3023 185
R1960 vdd.n3026 vdd.n936 185
R1961 vdd.n3001 vdd.n936 185
R1962 vdd.n3028 vdd.n3027 185
R1963 vdd.n3029 vdd.n3028 185
R1964 vdd.n926 vdd.n925 185
R1965 vdd.n927 vdd.n926 185
R1966 vdd.n3037 vdd.n3036 185
R1967 vdd.n3036 vdd.n3035 185
R1968 vdd.n3038 vdd.n924 185
R1969 vdd.n930 vdd.n924 185
R1970 vdd.n3040 vdd.n3039 185
R1971 vdd.n3041 vdd.n3040 185
R1972 vdd.n916 vdd.n915 185
R1973 vdd.n2989 vdd.n916 185
R1974 vdd.n3049 vdd.n3048 185
R1975 vdd.n3048 vdd.n3047 185
R1976 vdd.n3050 vdd.n914 185
R1977 vdd.n914 vdd.n911 185
R1978 vdd.n3052 vdd.n3051 185
R1979 vdd.n3053 vdd.n3052 185
R1980 vdd.n904 vdd.n903 185
R1981 vdd.n905 vdd.n904 185
R1982 vdd.n3061 vdd.n3060 185
R1983 vdd.n3060 vdd.n3059 185
R1984 vdd.n3062 vdd.n902 185
R1985 vdd.n2977 vdd.n902 185
R1986 vdd.n3064 vdd.n3063 185
R1987 vdd.n3065 vdd.n3064 185
R1988 vdd.n893 vdd.n892 185
R1989 vdd.n901 vdd.n893 185
R1990 vdd.n3073 vdd.n3072 185
R1991 vdd.n3072 vdd.n3071 185
R1992 vdd.n3074 vdd.n891 185
R1993 vdd.n891 vdd.n888 185
R1994 vdd.n3076 vdd.n3075 185
R1995 vdd.n3077 vdd.n3076 185
R1996 vdd.n880 vdd.n879 185
R1997 vdd.n881 vdd.n880 185
R1998 vdd.n3086 vdd.n3085 185
R1999 vdd.n3085 vdd.n3084 185
R2000 vdd.n3087 vdd.n878 185
R2001 vdd.n878 vdd.n874 185
R2002 vdd.n3089 vdd.n3088 185
R2003 vdd.n3090 vdd.n3089 185
R2004 vdd.n867 vdd.n866 185
R2005 vdd.n877 vdd.n867 185
R2006 vdd.n3098 vdd.n3097 185
R2007 vdd.n3097 vdd.n3096 185
R2008 vdd.n3099 vdd.n865 185
R2009 vdd.n870 vdd.n865 185
R2010 vdd.n3101 vdd.n3100 185
R2011 vdd.n3102 vdd.n3101 185
R2012 vdd.n856 vdd.n855 185
R2013 vdd.n864 vdd.n856 185
R2014 vdd.n3110 vdd.n3109 185
R2015 vdd.n3109 vdd.n3108 185
R2016 vdd.n3111 vdd.n854 185
R2017 vdd.n854 vdd.n851 185
R2018 vdd.n3113 vdd.n3112 185
R2019 vdd.n3114 vdd.n3113 185
R2020 vdd.n842 vdd.n841 185
R2021 vdd.n843 vdd.n842 185
R2022 vdd.n3167 vdd.n3166 185
R2023 vdd.n3166 vdd.n3165 185
R2024 vdd.n3168 vdd.n840 185
R2025 vdd.n846 vdd.n840 185
R2026 vdd.n3170 vdd.n3169 185
R2027 vdd.n3171 vdd.n3170 185
R2028 vdd.n810 vdd.n808 185
R2029 vdd.n808 vdd.n805 185
R2030 vdd.n3240 vdd.n3239 185
R2031 vdd.n3241 vdd.n3240 185
R2032 vdd.n2653 vdd.n2652 185
R2033 vdd.n2654 vdd.n2653 185
R2034 vdd.n996 vdd.n994 185
R2035 vdd.n994 vdd.n992 185
R2036 vdd.n2568 vdd.n1003 185
R2037 vdd.n2579 vdd.n1003 185
R2038 vdd.n2569 vdd.n1012 185
R2039 vdd.n2334 vdd.n1012 185
R2040 vdd.n2571 vdd.n2570 185
R2041 vdd.n2572 vdd.n2571 185
R2042 vdd.n2567 vdd.n1011 185
R2043 vdd.n1011 vdd.n1008 185
R2044 vdd.n2566 vdd.n2565 185
R2045 vdd.n2565 vdd.n2564 185
R2046 vdd.n1014 vdd.n1013 185
R2047 vdd.n1015 vdd.n1014 185
R2048 vdd.n2557 vdd.n2556 185
R2049 vdd.n2558 vdd.n2557 185
R2050 vdd.n2555 vdd.n1023 185
R2051 vdd.n2346 vdd.n1023 185
R2052 vdd.n2554 vdd.n2553 185
R2053 vdd.n2553 vdd.n2552 185
R2054 vdd.n1025 vdd.n1024 185
R2055 vdd.n1033 vdd.n1025 185
R2056 vdd.n2545 vdd.n2544 185
R2057 vdd.n2546 vdd.n2545 185
R2058 vdd.n2543 vdd.n1034 185
R2059 vdd.n1039 vdd.n1034 185
R2060 vdd.n2542 vdd.n2541 185
R2061 vdd.n2541 vdd.n2540 185
R2062 vdd.n1036 vdd.n1035 185
R2063 vdd.n2358 vdd.n1036 185
R2064 vdd.n2533 vdd.n2532 185
R2065 vdd.n2534 vdd.n2533 185
R2066 vdd.n2531 vdd.n1046 185
R2067 vdd.n1046 vdd.n1043 185
R2068 vdd.n2530 vdd.n2529 185
R2069 vdd.n2529 vdd.n2528 185
R2070 vdd.n1048 vdd.n1047 185
R2071 vdd.n1049 vdd.n1048 185
R2072 vdd.n2521 vdd.n2520 185
R2073 vdd.n2522 vdd.n2521 185
R2074 vdd.n2518 vdd.n1057 185
R2075 vdd.n1063 vdd.n1057 185
R2076 vdd.n2517 vdd.n2516 185
R2077 vdd.n2516 vdd.n2515 185
R2078 vdd.n1060 vdd.n1059 185
R2079 vdd.n1070 vdd.n1060 185
R2080 vdd.n2508 vdd.n2507 185
R2081 vdd.n2509 vdd.n2508 185
R2082 vdd.n2506 vdd.n1071 185
R2083 vdd.n1071 vdd.n1067 185
R2084 vdd.n2505 vdd.n2504 185
R2085 vdd.n2504 vdd.n2503 185
R2086 vdd.n1073 vdd.n1072 185
R2087 vdd.n1074 vdd.n1073 185
R2088 vdd.n2496 vdd.n2495 185
R2089 vdd.n2497 vdd.n2496 185
R2090 vdd.n2494 vdd.n1083 185
R2091 vdd.n1083 vdd.n1080 185
R2092 vdd.n2493 vdd.n2492 185
R2093 vdd.n2492 vdd.n2491 185
R2094 vdd.n1085 vdd.n1084 185
R2095 vdd.n1086 vdd.n1085 185
R2096 vdd.n2484 vdd.n2483 185
R2097 vdd.n2485 vdd.n2484 185
R2098 vdd.n2482 vdd.n1095 185
R2099 vdd.n1095 vdd.n1092 185
R2100 vdd.n2481 vdd.n2480 185
R2101 vdd.n2480 vdd.n2479 185
R2102 vdd.n1097 vdd.n1096 185
R2103 vdd.n1098 vdd.n1097 185
R2104 vdd.n2472 vdd.n2471 185
R2105 vdd.n2473 vdd.n2472 185
R2106 vdd.n2470 vdd.n1107 185
R2107 vdd.n1107 vdd.n1104 185
R2108 vdd.n2469 vdd.n2468 185
R2109 vdd.n2468 vdd.n2467 185
R2110 vdd.n2584 vdd.n967 185
R2111 vdd.n2726 vdd.n967 185
R2112 vdd.n2586 vdd.n2585 185
R2113 vdd.n2588 vdd.n2587 185
R2114 vdd.n2590 vdd.n2589 185
R2115 vdd.n2592 vdd.n2591 185
R2116 vdd.n2594 vdd.n2593 185
R2117 vdd.n2596 vdd.n2595 185
R2118 vdd.n2598 vdd.n2597 185
R2119 vdd.n2600 vdd.n2599 185
R2120 vdd.n2602 vdd.n2601 185
R2121 vdd.n2604 vdd.n2603 185
R2122 vdd.n2606 vdd.n2605 185
R2123 vdd.n2608 vdd.n2607 185
R2124 vdd.n2610 vdd.n2609 185
R2125 vdd.n2612 vdd.n2611 185
R2126 vdd.n2614 vdd.n2613 185
R2127 vdd.n2616 vdd.n2615 185
R2128 vdd.n2618 vdd.n2617 185
R2129 vdd.n2620 vdd.n2619 185
R2130 vdd.n2622 vdd.n2621 185
R2131 vdd.n2624 vdd.n2623 185
R2132 vdd.n2626 vdd.n2625 185
R2133 vdd.n2628 vdd.n2627 185
R2134 vdd.n2630 vdd.n2629 185
R2135 vdd.n2632 vdd.n2631 185
R2136 vdd.n2634 vdd.n2633 185
R2137 vdd.n2636 vdd.n2635 185
R2138 vdd.n2638 vdd.n2637 185
R2139 vdd.n2640 vdd.n2639 185
R2140 vdd.n2642 vdd.n2641 185
R2141 vdd.n2644 vdd.n2643 185
R2142 vdd.n2646 vdd.n2645 185
R2143 vdd.n2648 vdd.n2647 185
R2144 vdd.n2650 vdd.n2649 185
R2145 vdd.n2651 vdd.n995 185
R2146 vdd.n2583 vdd.n993 185
R2147 vdd.n2654 vdd.n993 185
R2148 vdd.n2582 vdd.n2581 185
R2149 vdd.n2581 vdd.n992 185
R2150 vdd.n2580 vdd.n1000 185
R2151 vdd.n2580 vdd.n2579 185
R2152 vdd.n2318 vdd.n1001 185
R2153 vdd.n2334 vdd.n1001 185
R2154 vdd.n2319 vdd.n1010 185
R2155 vdd.n2572 vdd.n1010 185
R2156 vdd.n2321 vdd.n2320 185
R2157 vdd.n2320 vdd.n1008 185
R2158 vdd.n2322 vdd.n1017 185
R2159 vdd.n2564 vdd.n1017 185
R2160 vdd.n2324 vdd.n2323 185
R2161 vdd.n2323 vdd.n1015 185
R2162 vdd.n2325 vdd.n1022 185
R2163 vdd.n2558 vdd.n1022 185
R2164 vdd.n2348 vdd.n2347 185
R2165 vdd.n2347 vdd.n2346 185
R2166 vdd.n2349 vdd.n1027 185
R2167 vdd.n2552 vdd.n1027 185
R2168 vdd.n2351 vdd.n2350 185
R2169 vdd.n2350 vdd.n1033 185
R2170 vdd.n2352 vdd.n1032 185
R2171 vdd.n2546 vdd.n1032 185
R2172 vdd.n2354 vdd.n2353 185
R2173 vdd.n2353 vdd.n1039 185
R2174 vdd.n2355 vdd.n1038 185
R2175 vdd.n2540 vdd.n1038 185
R2176 vdd.n2357 vdd.n2356 185
R2177 vdd.n2358 vdd.n2357 185
R2178 vdd.n2317 vdd.n1045 185
R2179 vdd.n2534 vdd.n1045 185
R2180 vdd.n2316 vdd.n2315 185
R2181 vdd.n2315 vdd.n1043 185
R2182 vdd.n2314 vdd.n1051 185
R2183 vdd.n2528 vdd.n1051 185
R2184 vdd.n2313 vdd.n2312 185
R2185 vdd.n2312 vdd.n1049 185
R2186 vdd.n2311 vdd.n1056 185
R2187 vdd.n2522 vdd.n1056 185
R2188 vdd.n2310 vdd.n2309 185
R2189 vdd.n2309 vdd.n1063 185
R2190 vdd.n2308 vdd.n1062 185
R2191 vdd.n2515 vdd.n1062 185
R2192 vdd.n2307 vdd.n2306 185
R2193 vdd.n2306 vdd.n1070 185
R2194 vdd.n2305 vdd.n1069 185
R2195 vdd.n2509 vdd.n1069 185
R2196 vdd.n2304 vdd.n2303 185
R2197 vdd.n2303 vdd.n1067 185
R2198 vdd.n2302 vdd.n1076 185
R2199 vdd.n2503 vdd.n1076 185
R2200 vdd.n2301 vdd.n2300 185
R2201 vdd.n2300 vdd.n1074 185
R2202 vdd.n2299 vdd.n1082 185
R2203 vdd.n2497 vdd.n1082 185
R2204 vdd.n2298 vdd.n2297 185
R2205 vdd.n2297 vdd.n1080 185
R2206 vdd.n2296 vdd.n1088 185
R2207 vdd.n2491 vdd.n1088 185
R2208 vdd.n2295 vdd.n2294 185
R2209 vdd.n2294 vdd.n1086 185
R2210 vdd.n2293 vdd.n1094 185
R2211 vdd.n2485 vdd.n1094 185
R2212 vdd.n2292 vdd.n2291 185
R2213 vdd.n2291 vdd.n1092 185
R2214 vdd.n2290 vdd.n1100 185
R2215 vdd.n2479 vdd.n1100 185
R2216 vdd.n2289 vdd.n2288 185
R2217 vdd.n2288 vdd.n1098 185
R2218 vdd.n2287 vdd.n1106 185
R2219 vdd.n2473 vdd.n1106 185
R2220 vdd.n2286 vdd.n2285 185
R2221 vdd.n2285 vdd.n1104 185
R2222 vdd.n2284 vdd.n1112 185
R2223 vdd.n2467 vdd.n1112 185
R2224 vdd.n1109 vdd.n1108 185
R2225 vdd.n2216 vdd.n2214 185
R2226 vdd.n2219 vdd.n2218 185
R2227 vdd.n2220 vdd.n2213 185
R2228 vdd.n2222 vdd.n2221 185
R2229 vdd.n2224 vdd.n2212 185
R2230 vdd.n2227 vdd.n2226 185
R2231 vdd.n2228 vdd.n2211 185
R2232 vdd.n2230 vdd.n2229 185
R2233 vdd.n2232 vdd.n2210 185
R2234 vdd.n2235 vdd.n2234 185
R2235 vdd.n2236 vdd.n2209 185
R2236 vdd.n2238 vdd.n2237 185
R2237 vdd.n2240 vdd.n2208 185
R2238 vdd.n2243 vdd.n2242 185
R2239 vdd.n2244 vdd.n2207 185
R2240 vdd.n2246 vdd.n2245 185
R2241 vdd.n2248 vdd.n2206 185
R2242 vdd.n2251 vdd.n2250 185
R2243 vdd.n2252 vdd.n1143 185
R2244 vdd.n2254 vdd.n2253 185
R2245 vdd.n2256 vdd.n1142 185
R2246 vdd.n2259 vdd.n2258 185
R2247 vdd.n2260 vdd.n1141 185
R2248 vdd.n2262 vdd.n2261 185
R2249 vdd.n2264 vdd.n1140 185
R2250 vdd.n2267 vdd.n2266 185
R2251 vdd.n2268 vdd.n1139 185
R2252 vdd.n2270 vdd.n2269 185
R2253 vdd.n2272 vdd.n1138 185
R2254 vdd.n2275 vdd.n2274 185
R2255 vdd.n2276 vdd.n1135 185
R2256 vdd.n2279 vdd.n2278 185
R2257 vdd.n2281 vdd.n1134 185
R2258 vdd.n2283 vdd.n2282 185
R2259 vdd.n2282 vdd.n1110 185
R2260 vdd.n327 vdd.n326 171.744
R2261 vdd.n326 vdd.n325 171.744
R2262 vdd.n325 vdd.n294 171.744
R2263 vdd.n318 vdd.n294 171.744
R2264 vdd.n318 vdd.n317 171.744
R2265 vdd.n317 vdd.n299 171.744
R2266 vdd.n310 vdd.n299 171.744
R2267 vdd.n310 vdd.n309 171.744
R2268 vdd.n309 vdd.n303 171.744
R2269 vdd.n268 vdd.n267 171.744
R2270 vdd.n267 vdd.n266 171.744
R2271 vdd.n266 vdd.n235 171.744
R2272 vdd.n259 vdd.n235 171.744
R2273 vdd.n259 vdd.n258 171.744
R2274 vdd.n258 vdd.n240 171.744
R2275 vdd.n251 vdd.n240 171.744
R2276 vdd.n251 vdd.n250 171.744
R2277 vdd.n250 vdd.n244 171.744
R2278 vdd.n225 vdd.n224 171.744
R2279 vdd.n224 vdd.n223 171.744
R2280 vdd.n223 vdd.n192 171.744
R2281 vdd.n216 vdd.n192 171.744
R2282 vdd.n216 vdd.n215 171.744
R2283 vdd.n215 vdd.n197 171.744
R2284 vdd.n208 vdd.n197 171.744
R2285 vdd.n208 vdd.n207 171.744
R2286 vdd.n207 vdd.n201 171.744
R2287 vdd.n166 vdd.n165 171.744
R2288 vdd.n165 vdd.n164 171.744
R2289 vdd.n164 vdd.n133 171.744
R2290 vdd.n157 vdd.n133 171.744
R2291 vdd.n157 vdd.n156 171.744
R2292 vdd.n156 vdd.n138 171.744
R2293 vdd.n149 vdd.n138 171.744
R2294 vdd.n149 vdd.n148 171.744
R2295 vdd.n148 vdd.n142 171.744
R2296 vdd.n124 vdd.n123 171.744
R2297 vdd.n123 vdd.n122 171.744
R2298 vdd.n122 vdd.n91 171.744
R2299 vdd.n115 vdd.n91 171.744
R2300 vdd.n115 vdd.n114 171.744
R2301 vdd.n114 vdd.n96 171.744
R2302 vdd.n107 vdd.n96 171.744
R2303 vdd.n107 vdd.n106 171.744
R2304 vdd.n106 vdd.n100 171.744
R2305 vdd.n65 vdd.n64 171.744
R2306 vdd.n64 vdd.n63 171.744
R2307 vdd.n63 vdd.n32 171.744
R2308 vdd.n56 vdd.n32 171.744
R2309 vdd.n56 vdd.n55 171.744
R2310 vdd.n55 vdd.n37 171.744
R2311 vdd.n48 vdd.n37 171.744
R2312 vdd.n48 vdd.n47 171.744
R2313 vdd.n47 vdd.n41 171.744
R2314 vdd.n1826 vdd.n1825 171.744
R2315 vdd.n1825 vdd.n1824 171.744
R2316 vdd.n1824 vdd.n1793 171.744
R2317 vdd.n1817 vdd.n1793 171.744
R2318 vdd.n1817 vdd.n1816 171.744
R2319 vdd.n1816 vdd.n1798 171.744
R2320 vdd.n1809 vdd.n1798 171.744
R2321 vdd.n1809 vdd.n1808 171.744
R2322 vdd.n1808 vdd.n1802 171.744
R2323 vdd.n1885 vdd.n1884 171.744
R2324 vdd.n1884 vdd.n1883 171.744
R2325 vdd.n1883 vdd.n1852 171.744
R2326 vdd.n1876 vdd.n1852 171.744
R2327 vdd.n1876 vdd.n1875 171.744
R2328 vdd.n1875 vdd.n1857 171.744
R2329 vdd.n1868 vdd.n1857 171.744
R2330 vdd.n1868 vdd.n1867 171.744
R2331 vdd.n1867 vdd.n1861 171.744
R2332 vdd.n1724 vdd.n1723 171.744
R2333 vdd.n1723 vdd.n1722 171.744
R2334 vdd.n1722 vdd.n1691 171.744
R2335 vdd.n1715 vdd.n1691 171.744
R2336 vdd.n1715 vdd.n1714 171.744
R2337 vdd.n1714 vdd.n1696 171.744
R2338 vdd.n1707 vdd.n1696 171.744
R2339 vdd.n1707 vdd.n1706 171.744
R2340 vdd.n1706 vdd.n1700 171.744
R2341 vdd.n1783 vdd.n1782 171.744
R2342 vdd.n1782 vdd.n1781 171.744
R2343 vdd.n1781 vdd.n1750 171.744
R2344 vdd.n1774 vdd.n1750 171.744
R2345 vdd.n1774 vdd.n1773 171.744
R2346 vdd.n1773 vdd.n1755 171.744
R2347 vdd.n1766 vdd.n1755 171.744
R2348 vdd.n1766 vdd.n1765 171.744
R2349 vdd.n1765 vdd.n1759 171.744
R2350 vdd.n1623 vdd.n1622 171.744
R2351 vdd.n1622 vdd.n1621 171.744
R2352 vdd.n1621 vdd.n1590 171.744
R2353 vdd.n1614 vdd.n1590 171.744
R2354 vdd.n1614 vdd.n1613 171.744
R2355 vdd.n1613 vdd.n1595 171.744
R2356 vdd.n1606 vdd.n1595 171.744
R2357 vdd.n1606 vdd.n1605 171.744
R2358 vdd.n1605 vdd.n1599 171.744
R2359 vdd.n1682 vdd.n1681 171.744
R2360 vdd.n1681 vdd.n1680 171.744
R2361 vdd.n1680 vdd.n1649 171.744
R2362 vdd.n1673 vdd.n1649 171.744
R2363 vdd.n1673 vdd.n1672 171.744
R2364 vdd.n1672 vdd.n1654 171.744
R2365 vdd.n1665 vdd.n1654 171.744
R2366 vdd.n1665 vdd.n1664 171.744
R2367 vdd.n1664 vdd.n1658 171.744
R2368 vdd.n468 vdd.n467 146.341
R2369 vdd.n474 vdd.n473 146.341
R2370 vdd.n478 vdd.n477 146.341
R2371 vdd.n484 vdd.n483 146.341
R2372 vdd.n488 vdd.n487 146.341
R2373 vdd.n494 vdd.n493 146.341
R2374 vdd.n498 vdd.n497 146.341
R2375 vdd.n504 vdd.n503 146.341
R2376 vdd.n508 vdd.n507 146.341
R2377 vdd.n514 vdd.n513 146.341
R2378 vdd.n518 vdd.n517 146.341
R2379 vdd.n524 vdd.n523 146.341
R2380 vdd.n528 vdd.n527 146.341
R2381 vdd.n534 vdd.n533 146.341
R2382 vdd.n538 vdd.n537 146.341
R2383 vdd.n544 vdd.n543 146.341
R2384 vdd.n548 vdd.n547 146.341
R2385 vdd.n554 vdd.n553 146.341
R2386 vdd.n558 vdd.n557 146.341
R2387 vdd.n564 vdd.n563 146.341
R2388 vdd.n568 vdd.n567 146.341
R2389 vdd.n574 vdd.n573 146.341
R2390 vdd.n578 vdd.n577 146.341
R2391 vdd.n584 vdd.n583 146.341
R2392 vdd.n588 vdd.n587 146.341
R2393 vdd.n594 vdd.n593 146.341
R2394 vdd.n598 vdd.n597 146.341
R2395 vdd.n604 vdd.n603 146.341
R2396 vdd.n608 vdd.n607 146.341
R2397 vdd.n614 vdd.n613 146.341
R2398 vdd.n616 vdd.n425 146.341
R2399 vdd.n3412 vdd.n685 146.341
R2400 vdd.n3412 vdd.n677 146.341
R2401 vdd.n3422 vdd.n677 146.341
R2402 vdd.n3422 vdd.n673 146.341
R2403 vdd.n3428 vdd.n673 146.341
R2404 vdd.n3428 vdd.n667 146.341
R2405 vdd.n3439 vdd.n667 146.341
R2406 vdd.n3439 vdd.n663 146.341
R2407 vdd.n3445 vdd.n663 146.341
R2408 vdd.n3445 vdd.n654 146.341
R2409 vdd.n3455 vdd.n654 146.341
R2410 vdd.n3455 vdd.n650 146.341
R2411 vdd.n3461 vdd.n650 146.341
R2412 vdd.n3461 vdd.n643 146.341
R2413 vdd.n3472 vdd.n643 146.341
R2414 vdd.n3472 vdd.n639 146.341
R2415 vdd.n3481 vdd.n639 146.341
R2416 vdd.n3481 vdd.n632 146.341
R2417 vdd.n3491 vdd.n632 146.341
R2418 vdd.n3492 vdd.n3491 146.341
R2419 vdd.n3492 vdd.n341 146.341
R2420 vdd.n342 vdd.n341 146.341
R2421 vdd.n343 vdd.n342 146.341
R2422 vdd.n3499 vdd.n343 146.341
R2423 vdd.n3499 vdd.n351 146.341
R2424 vdd.n352 vdd.n351 146.341
R2425 vdd.n353 vdd.n352 146.341
R2426 vdd.n3506 vdd.n353 146.341
R2427 vdd.n3506 vdd.n362 146.341
R2428 vdd.n363 vdd.n362 146.341
R2429 vdd.n364 vdd.n363 146.341
R2430 vdd.n3514 vdd.n364 146.341
R2431 vdd.n3514 vdd.n372 146.341
R2432 vdd.n373 vdd.n372 146.341
R2433 vdd.n374 vdd.n373 146.341
R2434 vdd.n3521 vdd.n374 146.341
R2435 vdd.n3521 vdd.n383 146.341
R2436 vdd.n384 vdd.n383 146.341
R2437 vdd.n385 vdd.n384 146.341
R2438 vdd.n3528 vdd.n385 146.341
R2439 vdd.n3528 vdd.n393 146.341
R2440 vdd.n725 vdd.n724 146.341
R2441 vdd.n728 vdd.n724 146.341
R2442 vdd.n734 vdd.n733 146.341
R2443 vdd.n3394 vdd.n3393 146.341
R2444 vdd.n3390 vdd.n3389 146.341
R2445 vdd.n3386 vdd.n3385 146.341
R2446 vdd.n3382 vdd.n3381 146.341
R2447 vdd.n3378 vdd.n3377 146.341
R2448 vdd.n3374 vdd.n3373 146.341
R2449 vdd.n3370 vdd.n3369 146.341
R2450 vdd.n3361 vdd.n3360 146.341
R2451 vdd.n3358 vdd.n3357 146.341
R2452 vdd.n3354 vdd.n3353 146.341
R2453 vdd.n3350 vdd.n3349 146.341
R2454 vdd.n3346 vdd.n3345 146.341
R2455 vdd.n3342 vdd.n3341 146.341
R2456 vdd.n3338 vdd.n3337 146.341
R2457 vdd.n3334 vdd.n3333 146.341
R2458 vdd.n3330 vdd.n3329 146.341
R2459 vdd.n3326 vdd.n3325 146.341
R2460 vdd.n3322 vdd.n3321 146.341
R2461 vdd.n3315 vdd.n3314 146.341
R2462 vdd.n3312 vdd.n3311 146.341
R2463 vdd.n3308 vdd.n3307 146.341
R2464 vdd.n3304 vdd.n3303 146.341
R2465 vdd.n3300 vdd.n3299 146.341
R2466 vdd.n3296 vdd.n3295 146.341
R2467 vdd.n3292 vdd.n3291 146.341
R2468 vdd.n3288 vdd.n3287 146.341
R2469 vdd.n3284 vdd.n3283 146.341
R2470 vdd.n3280 vdd.n3279 146.341
R2471 vdd.n3406 vdd.n691 146.341
R2472 vdd.n3414 vdd.n684 146.341
R2473 vdd.n3414 vdd.n680 146.341
R2474 vdd.n3420 vdd.n680 146.341
R2475 vdd.n3420 vdd.n672 146.341
R2476 vdd.n3431 vdd.n672 146.341
R2477 vdd.n3431 vdd.n668 146.341
R2478 vdd.n3437 vdd.n668 146.341
R2479 vdd.n3437 vdd.n661 146.341
R2480 vdd.n3447 vdd.n661 146.341
R2481 vdd.n3447 vdd.n657 146.341
R2482 vdd.n3453 vdd.n657 146.341
R2483 vdd.n3453 vdd.n649 146.341
R2484 vdd.n3464 vdd.n649 146.341
R2485 vdd.n3464 vdd.n645 146.341
R2486 vdd.n3470 vdd.n645 146.341
R2487 vdd.n3470 vdd.n638 146.341
R2488 vdd.n3483 vdd.n638 146.341
R2489 vdd.n3483 vdd.n634 146.341
R2490 vdd.n3489 vdd.n634 146.341
R2491 vdd.n3489 vdd.n338 146.341
R2492 vdd.n3578 vdd.n338 146.341
R2493 vdd.n3578 vdd.n339 146.341
R2494 vdd.n3574 vdd.n339 146.341
R2495 vdd.n3574 vdd.n345 146.341
R2496 vdd.n3570 vdd.n345 146.341
R2497 vdd.n3570 vdd.n350 146.341
R2498 vdd.n3566 vdd.n350 146.341
R2499 vdd.n3566 vdd.n354 146.341
R2500 vdd.n3562 vdd.n354 146.341
R2501 vdd.n3562 vdd.n360 146.341
R2502 vdd.n3558 vdd.n360 146.341
R2503 vdd.n3558 vdd.n365 146.341
R2504 vdd.n3554 vdd.n365 146.341
R2505 vdd.n3554 vdd.n371 146.341
R2506 vdd.n3550 vdd.n371 146.341
R2507 vdd.n3550 vdd.n376 146.341
R2508 vdd.n3546 vdd.n376 146.341
R2509 vdd.n3546 vdd.n382 146.341
R2510 vdd.n3542 vdd.n382 146.341
R2511 vdd.n3542 vdd.n387 146.341
R2512 vdd.n3538 vdd.n387 146.341
R2513 vdd.n2189 vdd.n2188 146.341
R2514 vdd.n2186 vdd.n1983 146.341
R2515 vdd.n2179 vdd.n1989 146.341
R2516 vdd.n2177 vdd.n2176 146.341
R2517 vdd.n2174 vdd.n1991 146.341
R2518 vdd.n2170 vdd.n2169 146.341
R2519 vdd.n2167 vdd.n1998 146.341
R2520 vdd.n2163 vdd.n2162 146.341
R2521 vdd.n2160 vdd.n2005 146.341
R2522 vdd.n2016 vdd.n2013 146.341
R2523 vdd.n2152 vdd.n2151 146.341
R2524 vdd.n2149 vdd.n2018 146.341
R2525 vdd.n2145 vdd.n2144 146.341
R2526 vdd.n2142 vdd.n2024 146.341
R2527 vdd.n2138 vdd.n2137 146.341
R2528 vdd.n2135 vdd.n2031 146.341
R2529 vdd.n2131 vdd.n2130 146.341
R2530 vdd.n2128 vdd.n2038 146.341
R2531 vdd.n2124 vdd.n2123 146.341
R2532 vdd.n2121 vdd.n2045 146.341
R2533 vdd.n2056 vdd.n2053 146.341
R2534 vdd.n2113 vdd.n2112 146.341
R2535 vdd.n2110 vdd.n2058 146.341
R2536 vdd.n2106 vdd.n2105 146.341
R2537 vdd.n2103 vdd.n2064 146.341
R2538 vdd.n2099 vdd.n2098 146.341
R2539 vdd.n2096 vdd.n2071 146.341
R2540 vdd.n2092 vdd.n2091 146.341
R2541 vdd.n2089 vdd.n2086 146.341
R2542 vdd.n2084 vdd.n2081 146.341
R2543 vdd.n2079 vdd.n1149 146.341
R2544 vdd.n1508 vdd.n1268 146.341
R2545 vdd.n1508 vdd.n1264 146.341
R2546 vdd.n1514 vdd.n1264 146.341
R2547 vdd.n1514 vdd.n1256 146.341
R2548 vdd.n1525 vdd.n1256 146.341
R2549 vdd.n1525 vdd.n1252 146.341
R2550 vdd.n1531 vdd.n1252 146.341
R2551 vdd.n1531 vdd.n1246 146.341
R2552 vdd.n1542 vdd.n1246 146.341
R2553 vdd.n1542 vdd.n1242 146.341
R2554 vdd.n1548 vdd.n1242 146.341
R2555 vdd.n1548 vdd.n1233 146.341
R2556 vdd.n1558 vdd.n1233 146.341
R2557 vdd.n1558 vdd.n1229 146.341
R2558 vdd.n1564 vdd.n1229 146.341
R2559 vdd.n1564 vdd.n1222 146.341
R2560 vdd.n1575 vdd.n1222 146.341
R2561 vdd.n1575 vdd.n1218 146.341
R2562 vdd.n1581 vdd.n1218 146.341
R2563 vdd.n1581 vdd.n1211 146.341
R2564 vdd.n1898 vdd.n1211 146.341
R2565 vdd.n1898 vdd.n1207 146.341
R2566 vdd.n1904 vdd.n1207 146.341
R2567 vdd.n1904 vdd.n1199 146.341
R2568 vdd.n1915 vdd.n1199 146.341
R2569 vdd.n1915 vdd.n1195 146.341
R2570 vdd.n1921 vdd.n1195 146.341
R2571 vdd.n1921 vdd.n1189 146.341
R2572 vdd.n1932 vdd.n1189 146.341
R2573 vdd.n1932 vdd.n1185 146.341
R2574 vdd.n1938 vdd.n1185 146.341
R2575 vdd.n1938 vdd.n1176 146.341
R2576 vdd.n1948 vdd.n1176 146.341
R2577 vdd.n1948 vdd.n1172 146.341
R2578 vdd.n1954 vdd.n1172 146.341
R2579 vdd.n1954 vdd.n1166 146.341
R2580 vdd.n1965 vdd.n1166 146.341
R2581 vdd.n1965 vdd.n1161 146.341
R2582 vdd.n1973 vdd.n1161 146.341
R2583 vdd.n1973 vdd.n1151 146.341
R2584 vdd.n2197 vdd.n1151 146.341
R2585 vdd.n1497 vdd.n1273 146.341
R2586 vdd.n1497 vdd.n1306 146.341
R2587 vdd.n1310 vdd.n1309 146.341
R2588 vdd.n1312 vdd.n1311 146.341
R2589 vdd.n1316 vdd.n1315 146.341
R2590 vdd.n1318 vdd.n1317 146.341
R2591 vdd.n1322 vdd.n1321 146.341
R2592 vdd.n1324 vdd.n1323 146.341
R2593 vdd.n1328 vdd.n1327 146.341
R2594 vdd.n1330 vdd.n1329 146.341
R2595 vdd.n1336 vdd.n1335 146.341
R2596 vdd.n1338 vdd.n1337 146.341
R2597 vdd.n1342 vdd.n1341 146.341
R2598 vdd.n1344 vdd.n1343 146.341
R2599 vdd.n1348 vdd.n1347 146.341
R2600 vdd.n1350 vdd.n1349 146.341
R2601 vdd.n1354 vdd.n1353 146.341
R2602 vdd.n1356 vdd.n1355 146.341
R2603 vdd.n1360 vdd.n1359 146.341
R2604 vdd.n1362 vdd.n1361 146.341
R2605 vdd.n1434 vdd.n1365 146.341
R2606 vdd.n1367 vdd.n1366 146.341
R2607 vdd.n1371 vdd.n1370 146.341
R2608 vdd.n1373 vdd.n1372 146.341
R2609 vdd.n1377 vdd.n1376 146.341
R2610 vdd.n1379 vdd.n1378 146.341
R2611 vdd.n1383 vdd.n1382 146.341
R2612 vdd.n1385 vdd.n1384 146.341
R2613 vdd.n1389 vdd.n1388 146.341
R2614 vdd.n1391 vdd.n1390 146.341
R2615 vdd.n1395 vdd.n1394 146.341
R2616 vdd.n1396 vdd.n1304 146.341
R2617 vdd.n1506 vdd.n1269 146.341
R2618 vdd.n1506 vdd.n1262 146.341
R2619 vdd.n1517 vdd.n1262 146.341
R2620 vdd.n1517 vdd.n1258 146.341
R2621 vdd.n1523 vdd.n1258 146.341
R2622 vdd.n1523 vdd.n1251 146.341
R2623 vdd.n1534 vdd.n1251 146.341
R2624 vdd.n1534 vdd.n1247 146.341
R2625 vdd.n1540 vdd.n1247 146.341
R2626 vdd.n1540 vdd.n1240 146.341
R2627 vdd.n1550 vdd.n1240 146.341
R2628 vdd.n1550 vdd.n1236 146.341
R2629 vdd.n1556 vdd.n1236 146.341
R2630 vdd.n1556 vdd.n1228 146.341
R2631 vdd.n1567 vdd.n1228 146.341
R2632 vdd.n1567 vdd.n1224 146.341
R2633 vdd.n1573 vdd.n1224 146.341
R2634 vdd.n1573 vdd.n1217 146.341
R2635 vdd.n1583 vdd.n1217 146.341
R2636 vdd.n1583 vdd.n1213 146.341
R2637 vdd.n1896 vdd.n1213 146.341
R2638 vdd.n1896 vdd.n1205 146.341
R2639 vdd.n1907 vdd.n1205 146.341
R2640 vdd.n1907 vdd.n1201 146.341
R2641 vdd.n1913 vdd.n1201 146.341
R2642 vdd.n1913 vdd.n1194 146.341
R2643 vdd.n1924 vdd.n1194 146.341
R2644 vdd.n1924 vdd.n1190 146.341
R2645 vdd.n1930 vdd.n1190 146.341
R2646 vdd.n1930 vdd.n1183 146.341
R2647 vdd.n1940 vdd.n1183 146.341
R2648 vdd.n1940 vdd.n1179 146.341
R2649 vdd.n1946 vdd.n1179 146.341
R2650 vdd.n1946 vdd.n1171 146.341
R2651 vdd.n1957 vdd.n1171 146.341
R2652 vdd.n1957 vdd.n1167 146.341
R2653 vdd.n1963 vdd.n1167 146.341
R2654 vdd.n1963 vdd.n1159 146.341
R2655 vdd.n1976 vdd.n1159 146.341
R2656 vdd.n1976 vdd.n1154 146.341
R2657 vdd.n2195 vdd.n1154 146.341
R2658 vdd.n1136 vdd.t32 127.284
R2659 vdd.n997 vdd.t69 127.284
R2660 vdd.n1130 vdd.t96 127.284
R2661 vdd.n988 vdd.t92 127.284
R2662 vdd.n885 vdd.t42 127.284
R2663 vdd.n885 vdd.t43 127.284
R2664 vdd.n2761 vdd.t87 127.284
R2665 vdd.n832 vdd.t55 127.284
R2666 vdd.n2830 vdd.t74 127.284
R2667 vdd.n799 vdd.t27 127.284
R2668 vdd.n1058 vdd.t83 127.284
R2669 vdd.n1058 vdd.t84 127.284
R2670 vdd.n22 vdd.n20 117.314
R2671 vdd.n17 vdd.n15 117.314
R2672 vdd.n27 vdd.n26 116.927
R2673 vdd.n24 vdd.n23 116.927
R2674 vdd.n22 vdd.n21 116.927
R2675 vdd.n17 vdd.n16 116.927
R2676 vdd.n19 vdd.n18 116.927
R2677 vdd.n27 vdd.n25 116.927
R2678 vdd.n1137 vdd.t31 111.188
R2679 vdd.n998 vdd.t70 111.188
R2680 vdd.n1131 vdd.t95 111.188
R2681 vdd.n989 vdd.t93 111.188
R2682 vdd.n2762 vdd.t86 111.188
R2683 vdd.n833 vdd.t56 111.188
R2684 vdd.n2831 vdd.t73 111.188
R2685 vdd.n800 vdd.t28 111.188
R2686 vdd.n3016 vdd.n938 99.5127
R2687 vdd.n3024 vdd.n938 99.5127
R2688 vdd.n3024 vdd.n936 99.5127
R2689 vdd.n3028 vdd.n936 99.5127
R2690 vdd.n3028 vdd.n926 99.5127
R2691 vdd.n3036 vdd.n926 99.5127
R2692 vdd.n3036 vdd.n924 99.5127
R2693 vdd.n3040 vdd.n924 99.5127
R2694 vdd.n3040 vdd.n916 99.5127
R2695 vdd.n3048 vdd.n916 99.5127
R2696 vdd.n3048 vdd.n914 99.5127
R2697 vdd.n3052 vdd.n914 99.5127
R2698 vdd.n3052 vdd.n904 99.5127
R2699 vdd.n3060 vdd.n904 99.5127
R2700 vdd.n3060 vdd.n902 99.5127
R2701 vdd.n3064 vdd.n902 99.5127
R2702 vdd.n3064 vdd.n893 99.5127
R2703 vdd.n3072 vdd.n893 99.5127
R2704 vdd.n3072 vdd.n891 99.5127
R2705 vdd.n3076 vdd.n891 99.5127
R2706 vdd.n3076 vdd.n880 99.5127
R2707 vdd.n3085 vdd.n880 99.5127
R2708 vdd.n3085 vdd.n878 99.5127
R2709 vdd.n3089 vdd.n878 99.5127
R2710 vdd.n3089 vdd.n867 99.5127
R2711 vdd.n3097 vdd.n867 99.5127
R2712 vdd.n3097 vdd.n865 99.5127
R2713 vdd.n3101 vdd.n865 99.5127
R2714 vdd.n3101 vdd.n856 99.5127
R2715 vdd.n3109 vdd.n856 99.5127
R2716 vdd.n3109 vdd.n854 99.5127
R2717 vdd.n3113 vdd.n854 99.5127
R2718 vdd.n3113 vdd.n842 99.5127
R2719 vdd.n3166 vdd.n842 99.5127
R2720 vdd.n3166 vdd.n840 99.5127
R2721 vdd.n3170 vdd.n840 99.5127
R2722 vdd.n3170 vdd.n808 99.5127
R2723 vdd.n3240 vdd.n808 99.5127
R2724 vdd.n3236 vdd.n809 99.5127
R2725 vdd.n3234 vdd.n3233 99.5127
R2726 vdd.n3231 vdd.n813 99.5127
R2727 vdd.n3227 vdd.n3226 99.5127
R2728 vdd.n3224 vdd.n816 99.5127
R2729 vdd.n3220 vdd.n3219 99.5127
R2730 vdd.n3217 vdd.n819 99.5127
R2731 vdd.n3213 vdd.n3212 99.5127
R2732 vdd.n3210 vdd.n3208 99.5127
R2733 vdd.n3206 vdd.n822 99.5127
R2734 vdd.n3202 vdd.n3201 99.5127
R2735 vdd.n3199 vdd.n825 99.5127
R2736 vdd.n3195 vdd.n3194 99.5127
R2737 vdd.n3192 vdd.n828 99.5127
R2738 vdd.n3188 vdd.n3187 99.5127
R2739 vdd.n3185 vdd.n831 99.5127
R2740 vdd.n3180 vdd.n3179 99.5127
R2741 vdd.n2898 vdd.n944 99.5127
R2742 vdd.n2898 vdd.n939 99.5127
R2743 vdd.n3000 vdd.n939 99.5127
R2744 vdd.n3000 vdd.n934 99.5127
R2745 vdd.n2996 vdd.n934 99.5127
R2746 vdd.n2996 vdd.n928 99.5127
R2747 vdd.n2993 vdd.n928 99.5127
R2748 vdd.n2993 vdd.n922 99.5127
R2749 vdd.n2990 vdd.n922 99.5127
R2750 vdd.n2990 vdd.n917 99.5127
R2751 vdd.n2940 vdd.n917 99.5127
R2752 vdd.n2940 vdd.n912 99.5127
R2753 vdd.n2943 vdd.n912 99.5127
R2754 vdd.n2943 vdd.n906 99.5127
R2755 vdd.n2976 vdd.n906 99.5127
R2756 vdd.n2976 vdd.n899 99.5127
R2757 vdd.n2972 vdd.n899 99.5127
R2758 vdd.n2972 vdd.n894 99.5127
R2759 vdd.n2969 vdd.n894 99.5127
R2760 vdd.n2969 vdd.n889 99.5127
R2761 vdd.n2966 vdd.n889 99.5127
R2762 vdd.n2966 vdd.n882 99.5127
R2763 vdd.n2963 vdd.n882 99.5127
R2764 vdd.n2963 vdd.n875 99.5127
R2765 vdd.n2960 vdd.n875 99.5127
R2766 vdd.n2960 vdd.n868 99.5127
R2767 vdd.n2957 vdd.n868 99.5127
R2768 vdd.n2957 vdd.n862 99.5127
R2769 vdd.n2954 vdd.n862 99.5127
R2770 vdd.n2954 vdd.n857 99.5127
R2771 vdd.n2951 vdd.n857 99.5127
R2772 vdd.n2951 vdd.n852 99.5127
R2773 vdd.n2948 vdd.n852 99.5127
R2774 vdd.n2948 vdd.n844 99.5127
R2775 vdd.n844 vdd.n837 99.5127
R2776 vdd.n3172 vdd.n837 99.5127
R2777 vdd.n3173 vdd.n3172 99.5127
R2778 vdd.n3173 vdd.n806 99.5127
R2779 vdd.n3012 vdd.n949 99.5127
R2780 vdd.n2832 vdd.n949 99.5127
R2781 vdd.n2836 vdd.n2835 99.5127
R2782 vdd.n2840 vdd.n2839 99.5127
R2783 vdd.n2844 vdd.n2843 99.5127
R2784 vdd.n2848 vdd.n2847 99.5127
R2785 vdd.n2852 vdd.n2851 99.5127
R2786 vdd.n2856 vdd.n2855 99.5127
R2787 vdd.n2860 vdd.n2859 99.5127
R2788 vdd.n2864 vdd.n2863 99.5127
R2789 vdd.n2868 vdd.n2867 99.5127
R2790 vdd.n2872 vdd.n2871 99.5127
R2791 vdd.n2876 vdd.n2875 99.5127
R2792 vdd.n2880 vdd.n2879 99.5127
R2793 vdd.n2884 vdd.n2883 99.5127
R2794 vdd.n2888 vdd.n2887 99.5127
R2795 vdd.n2893 vdd.n2892 99.5127
R2796 vdd.n2725 vdd.n986 99.5127
R2797 vdd.n2721 vdd.n2720 99.5127
R2798 vdd.n2717 vdd.n2716 99.5127
R2799 vdd.n2713 vdd.n2712 99.5127
R2800 vdd.n2709 vdd.n2708 99.5127
R2801 vdd.n2705 vdd.n2704 99.5127
R2802 vdd.n2701 vdd.n2700 99.5127
R2803 vdd.n2697 vdd.n2696 99.5127
R2804 vdd.n2693 vdd.n2692 99.5127
R2805 vdd.n2689 vdd.n2688 99.5127
R2806 vdd.n2685 vdd.n2684 99.5127
R2807 vdd.n2681 vdd.n2680 99.5127
R2808 vdd.n2677 vdd.n2676 99.5127
R2809 vdd.n2673 vdd.n2672 99.5127
R2810 vdd.n2669 vdd.n2668 99.5127
R2811 vdd.n2665 vdd.n2664 99.5127
R2812 vdd.n2660 vdd.n2659 99.5127
R2813 vdd.n2392 vdd.n1111 99.5127
R2814 vdd.n2392 vdd.n1105 99.5127
R2815 vdd.n2389 vdd.n1105 99.5127
R2816 vdd.n2389 vdd.n1099 99.5127
R2817 vdd.n2386 vdd.n1099 99.5127
R2818 vdd.n2386 vdd.n1093 99.5127
R2819 vdd.n2383 vdd.n1093 99.5127
R2820 vdd.n2383 vdd.n1087 99.5127
R2821 vdd.n2380 vdd.n1087 99.5127
R2822 vdd.n2380 vdd.n1081 99.5127
R2823 vdd.n2377 vdd.n1081 99.5127
R2824 vdd.n2377 vdd.n1075 99.5127
R2825 vdd.n2374 vdd.n1075 99.5127
R2826 vdd.n2374 vdd.n1068 99.5127
R2827 vdd.n2371 vdd.n1068 99.5127
R2828 vdd.n2371 vdd.n1061 99.5127
R2829 vdd.n2368 vdd.n1061 99.5127
R2830 vdd.n2368 vdd.n1055 99.5127
R2831 vdd.n2365 vdd.n1055 99.5127
R2832 vdd.n2365 vdd.n1050 99.5127
R2833 vdd.n2362 vdd.n1050 99.5127
R2834 vdd.n2362 vdd.n1044 99.5127
R2835 vdd.n2359 vdd.n1044 99.5127
R2836 vdd.n2359 vdd.n1037 99.5127
R2837 vdd.n2326 vdd.n1037 99.5127
R2838 vdd.n2326 vdd.n1031 99.5127
R2839 vdd.n2329 vdd.n1031 99.5127
R2840 vdd.n2329 vdd.n1026 99.5127
R2841 vdd.n2345 vdd.n1026 99.5127
R2842 vdd.n2345 vdd.n1021 99.5127
R2843 vdd.n2341 vdd.n1021 99.5127
R2844 vdd.n2341 vdd.n1016 99.5127
R2845 vdd.n2338 vdd.n1016 99.5127
R2846 vdd.n2338 vdd.n1009 99.5127
R2847 vdd.n2335 vdd.n1009 99.5127
R2848 vdd.n2335 vdd.n1002 99.5127
R2849 vdd.n1002 vdd.n991 99.5127
R2850 vdd.n2655 vdd.n991 99.5127
R2851 vdd.n2462 vdd.n2460 99.5127
R2852 vdd.n2460 vdd.n2459 99.5127
R2853 vdd.n2456 vdd.n2455 99.5127
R2854 vdd.n2453 vdd.n1117 99.5127
R2855 vdd.n2449 vdd.n2447 99.5127
R2856 vdd.n2445 vdd.n1119 99.5127
R2857 vdd.n2441 vdd.n2439 99.5127
R2858 vdd.n2437 vdd.n1121 99.5127
R2859 vdd.n2433 vdd.n2431 99.5127
R2860 vdd.n2429 vdd.n1123 99.5127
R2861 vdd.n2425 vdd.n2423 99.5127
R2862 vdd.n2421 vdd.n1125 99.5127
R2863 vdd.n2417 vdd.n2415 99.5127
R2864 vdd.n2413 vdd.n1127 99.5127
R2865 vdd.n2409 vdd.n2407 99.5127
R2866 vdd.n2405 vdd.n1129 99.5127
R2867 vdd.n2400 vdd.n2398 99.5127
R2868 vdd.n2466 vdd.n1103 99.5127
R2869 vdd.n2474 vdd.n1103 99.5127
R2870 vdd.n2474 vdd.n1101 99.5127
R2871 vdd.n2478 vdd.n1101 99.5127
R2872 vdd.n2478 vdd.n1091 99.5127
R2873 vdd.n2486 vdd.n1091 99.5127
R2874 vdd.n2486 vdd.n1089 99.5127
R2875 vdd.n2490 vdd.n1089 99.5127
R2876 vdd.n2490 vdd.n1079 99.5127
R2877 vdd.n2498 vdd.n1079 99.5127
R2878 vdd.n2498 vdd.n1077 99.5127
R2879 vdd.n2502 vdd.n1077 99.5127
R2880 vdd.n2502 vdd.n1066 99.5127
R2881 vdd.n2510 vdd.n1066 99.5127
R2882 vdd.n2510 vdd.n1064 99.5127
R2883 vdd.n2514 vdd.n1064 99.5127
R2884 vdd.n2514 vdd.n1054 99.5127
R2885 vdd.n2523 vdd.n1054 99.5127
R2886 vdd.n2523 vdd.n1052 99.5127
R2887 vdd.n2527 vdd.n1052 99.5127
R2888 vdd.n2527 vdd.n1042 99.5127
R2889 vdd.n2535 vdd.n1042 99.5127
R2890 vdd.n2535 vdd.n1040 99.5127
R2891 vdd.n2539 vdd.n1040 99.5127
R2892 vdd.n2539 vdd.n1030 99.5127
R2893 vdd.n2547 vdd.n1030 99.5127
R2894 vdd.n2547 vdd.n1028 99.5127
R2895 vdd.n2551 vdd.n1028 99.5127
R2896 vdd.n2551 vdd.n1020 99.5127
R2897 vdd.n2559 vdd.n1020 99.5127
R2898 vdd.n2559 vdd.n1018 99.5127
R2899 vdd.n2563 vdd.n1018 99.5127
R2900 vdd.n2563 vdd.n1007 99.5127
R2901 vdd.n2573 vdd.n1007 99.5127
R2902 vdd.n2573 vdd.n1004 99.5127
R2903 vdd.n2578 vdd.n1004 99.5127
R2904 vdd.n2578 vdd.n1005 99.5127
R2905 vdd.n1005 vdd.n985 99.5127
R2906 vdd.n3156 vdd.n3155 99.5127
R2907 vdd.n3153 vdd.n3119 99.5127
R2908 vdd.n3149 vdd.n3148 99.5127
R2909 vdd.n3146 vdd.n3122 99.5127
R2910 vdd.n3142 vdd.n3141 99.5127
R2911 vdd.n3139 vdd.n3125 99.5127
R2912 vdd.n3135 vdd.n3134 99.5127
R2913 vdd.n3132 vdd.n3129 99.5127
R2914 vdd.n3273 vdd.n787 99.5127
R2915 vdd.n3271 vdd.n3270 99.5127
R2916 vdd.n3268 vdd.n789 99.5127
R2917 vdd.n3264 vdd.n3263 99.5127
R2918 vdd.n3261 vdd.n792 99.5127
R2919 vdd.n3257 vdd.n3256 99.5127
R2920 vdd.n3254 vdd.n795 99.5127
R2921 vdd.n3250 vdd.n3249 99.5127
R2922 vdd.n3247 vdd.n798 99.5127
R2923 vdd.n3005 vdd.n945 99.5127
R2924 vdd.n3005 vdd.n940 99.5127
R2925 vdd.n3002 vdd.n940 99.5127
R2926 vdd.n3002 vdd.n935 99.5127
R2927 vdd.n2902 vdd.n935 99.5127
R2928 vdd.n2902 vdd.n929 99.5127
R2929 vdd.n2905 vdd.n929 99.5127
R2930 vdd.n2905 vdd.n923 99.5127
R2931 vdd.n2988 vdd.n923 99.5127
R2932 vdd.n2988 vdd.n918 99.5127
R2933 vdd.n2984 vdd.n918 99.5127
R2934 vdd.n2984 vdd.n913 99.5127
R2935 vdd.n2981 vdd.n913 99.5127
R2936 vdd.n2981 vdd.n907 99.5127
R2937 vdd.n2978 vdd.n907 99.5127
R2938 vdd.n2978 vdd.n900 99.5127
R2939 vdd.n2937 vdd.n900 99.5127
R2940 vdd.n2937 vdd.n895 99.5127
R2941 vdd.n2934 vdd.n895 99.5127
R2942 vdd.n2934 vdd.n890 99.5127
R2943 vdd.n2931 vdd.n890 99.5127
R2944 vdd.n2931 vdd.n883 99.5127
R2945 vdd.n2928 vdd.n883 99.5127
R2946 vdd.n2928 vdd.n876 99.5127
R2947 vdd.n2925 vdd.n876 99.5127
R2948 vdd.n2925 vdd.n869 99.5127
R2949 vdd.n2922 vdd.n869 99.5127
R2950 vdd.n2922 vdd.n863 99.5127
R2951 vdd.n2919 vdd.n863 99.5127
R2952 vdd.n2919 vdd.n858 99.5127
R2953 vdd.n2916 vdd.n858 99.5127
R2954 vdd.n2916 vdd.n853 99.5127
R2955 vdd.n2913 vdd.n853 99.5127
R2956 vdd.n2913 vdd.n845 99.5127
R2957 vdd.n2910 vdd.n845 99.5127
R2958 vdd.n2910 vdd.n838 99.5127
R2959 vdd.n838 vdd.n804 99.5127
R2960 vdd.n3242 vdd.n804 99.5127
R2961 vdd.n2766 vdd.n2765 99.5127
R2962 vdd.n2770 vdd.n2769 99.5127
R2963 vdd.n2774 vdd.n2773 99.5127
R2964 vdd.n2778 vdd.n2777 99.5127
R2965 vdd.n2782 vdd.n2781 99.5127
R2966 vdd.n2786 vdd.n2785 99.5127
R2967 vdd.n2790 vdd.n2789 99.5127
R2968 vdd.n2794 vdd.n2793 99.5127
R2969 vdd.n2798 vdd.n2797 99.5127
R2970 vdd.n2802 vdd.n2801 99.5127
R2971 vdd.n2806 vdd.n2805 99.5127
R2972 vdd.n2810 vdd.n2809 99.5127
R2973 vdd.n2814 vdd.n2813 99.5127
R2974 vdd.n2818 vdd.n2817 99.5127
R2975 vdd.n2822 vdd.n2821 99.5127
R2976 vdd.n2826 vdd.n2825 99.5127
R2977 vdd.n3009 vdd.n2760 99.5127
R2978 vdd.n3018 vdd.n941 99.5127
R2979 vdd.n3022 vdd.n941 99.5127
R2980 vdd.n3022 vdd.n933 99.5127
R2981 vdd.n3030 vdd.n933 99.5127
R2982 vdd.n3030 vdd.n931 99.5127
R2983 vdd.n3034 vdd.n931 99.5127
R2984 vdd.n3034 vdd.n921 99.5127
R2985 vdd.n3042 vdd.n921 99.5127
R2986 vdd.n3042 vdd.n919 99.5127
R2987 vdd.n3046 vdd.n919 99.5127
R2988 vdd.n3046 vdd.n910 99.5127
R2989 vdd.n3054 vdd.n910 99.5127
R2990 vdd.n3054 vdd.n908 99.5127
R2991 vdd.n3058 vdd.n908 99.5127
R2992 vdd.n3058 vdd.n898 99.5127
R2993 vdd.n3066 vdd.n898 99.5127
R2994 vdd.n3066 vdd.n896 99.5127
R2995 vdd.n3070 vdd.n896 99.5127
R2996 vdd.n3070 vdd.n887 99.5127
R2997 vdd.n3078 vdd.n887 99.5127
R2998 vdd.n3078 vdd.n884 99.5127
R2999 vdd.n3083 vdd.n884 99.5127
R3000 vdd.n3083 vdd.n873 99.5127
R3001 vdd.n3091 vdd.n873 99.5127
R3002 vdd.n3091 vdd.n871 99.5127
R3003 vdd.n3095 vdd.n871 99.5127
R3004 vdd.n3095 vdd.n861 99.5127
R3005 vdd.n3103 vdd.n861 99.5127
R3006 vdd.n3103 vdd.n859 99.5127
R3007 vdd.n3107 vdd.n859 99.5127
R3008 vdd.n3107 vdd.n850 99.5127
R3009 vdd.n3115 vdd.n850 99.5127
R3010 vdd.n3115 vdd.n847 99.5127
R3011 vdd.n3164 vdd.n847 99.5127
R3012 vdd.n3164 vdd.n848 99.5127
R3013 vdd.n848 vdd.n839 99.5127
R3014 vdd.n3159 vdd.n839 99.5127
R3015 vdd.n3159 vdd.n807 99.5127
R3016 vdd.n2649 vdd.n2648 99.5127
R3017 vdd.n2645 vdd.n2644 99.5127
R3018 vdd.n2641 vdd.n2640 99.5127
R3019 vdd.n2637 vdd.n2636 99.5127
R3020 vdd.n2633 vdd.n2632 99.5127
R3021 vdd.n2629 vdd.n2628 99.5127
R3022 vdd.n2625 vdd.n2624 99.5127
R3023 vdd.n2621 vdd.n2620 99.5127
R3024 vdd.n2617 vdd.n2616 99.5127
R3025 vdd.n2613 vdd.n2612 99.5127
R3026 vdd.n2609 vdd.n2608 99.5127
R3027 vdd.n2605 vdd.n2604 99.5127
R3028 vdd.n2601 vdd.n2600 99.5127
R3029 vdd.n2597 vdd.n2596 99.5127
R3030 vdd.n2593 vdd.n2592 99.5127
R3031 vdd.n2589 vdd.n2588 99.5127
R3032 vdd.n2585 vdd.n967 99.5127
R3033 vdd.n2285 vdd.n1112 99.5127
R3034 vdd.n2285 vdd.n1106 99.5127
R3035 vdd.n2288 vdd.n1106 99.5127
R3036 vdd.n2288 vdd.n1100 99.5127
R3037 vdd.n2291 vdd.n1100 99.5127
R3038 vdd.n2291 vdd.n1094 99.5127
R3039 vdd.n2294 vdd.n1094 99.5127
R3040 vdd.n2294 vdd.n1088 99.5127
R3041 vdd.n2297 vdd.n1088 99.5127
R3042 vdd.n2297 vdd.n1082 99.5127
R3043 vdd.n2300 vdd.n1082 99.5127
R3044 vdd.n2300 vdd.n1076 99.5127
R3045 vdd.n2303 vdd.n1076 99.5127
R3046 vdd.n2303 vdd.n1069 99.5127
R3047 vdd.n2306 vdd.n1069 99.5127
R3048 vdd.n2306 vdd.n1062 99.5127
R3049 vdd.n2309 vdd.n1062 99.5127
R3050 vdd.n2309 vdd.n1056 99.5127
R3051 vdd.n2312 vdd.n1056 99.5127
R3052 vdd.n2312 vdd.n1051 99.5127
R3053 vdd.n2315 vdd.n1051 99.5127
R3054 vdd.n2315 vdd.n1045 99.5127
R3055 vdd.n2357 vdd.n1045 99.5127
R3056 vdd.n2357 vdd.n1038 99.5127
R3057 vdd.n2353 vdd.n1038 99.5127
R3058 vdd.n2353 vdd.n1032 99.5127
R3059 vdd.n2350 vdd.n1032 99.5127
R3060 vdd.n2350 vdd.n1027 99.5127
R3061 vdd.n2347 vdd.n1027 99.5127
R3062 vdd.n2347 vdd.n1022 99.5127
R3063 vdd.n2323 vdd.n1022 99.5127
R3064 vdd.n2323 vdd.n1017 99.5127
R3065 vdd.n2320 vdd.n1017 99.5127
R3066 vdd.n2320 vdd.n1010 99.5127
R3067 vdd.n1010 vdd.n1001 99.5127
R3068 vdd.n2580 vdd.n1001 99.5127
R3069 vdd.n2581 vdd.n2580 99.5127
R3070 vdd.n2581 vdd.n993 99.5127
R3071 vdd.n2218 vdd.n2216 99.5127
R3072 vdd.n2222 vdd.n2213 99.5127
R3073 vdd.n2226 vdd.n2224 99.5127
R3074 vdd.n2230 vdd.n2211 99.5127
R3075 vdd.n2234 vdd.n2232 99.5127
R3076 vdd.n2238 vdd.n2209 99.5127
R3077 vdd.n2242 vdd.n2240 99.5127
R3078 vdd.n2246 vdd.n2207 99.5127
R3079 vdd.n2250 vdd.n2248 99.5127
R3080 vdd.n2254 vdd.n1143 99.5127
R3081 vdd.n2258 vdd.n2256 99.5127
R3082 vdd.n2262 vdd.n1141 99.5127
R3083 vdd.n2266 vdd.n2264 99.5127
R3084 vdd.n2270 vdd.n1139 99.5127
R3085 vdd.n2274 vdd.n2272 99.5127
R3086 vdd.n2279 vdd.n1135 99.5127
R3087 vdd.n2282 vdd.n2281 99.5127
R3088 vdd.n2468 vdd.n1107 99.5127
R3089 vdd.n2472 vdd.n1107 99.5127
R3090 vdd.n2472 vdd.n1097 99.5127
R3091 vdd.n2480 vdd.n1097 99.5127
R3092 vdd.n2480 vdd.n1095 99.5127
R3093 vdd.n2484 vdd.n1095 99.5127
R3094 vdd.n2484 vdd.n1085 99.5127
R3095 vdd.n2492 vdd.n1085 99.5127
R3096 vdd.n2492 vdd.n1083 99.5127
R3097 vdd.n2496 vdd.n1083 99.5127
R3098 vdd.n2496 vdd.n1073 99.5127
R3099 vdd.n2504 vdd.n1073 99.5127
R3100 vdd.n2504 vdd.n1071 99.5127
R3101 vdd.n2508 vdd.n1071 99.5127
R3102 vdd.n2508 vdd.n1060 99.5127
R3103 vdd.n2516 vdd.n1060 99.5127
R3104 vdd.n2516 vdd.n1057 99.5127
R3105 vdd.n2521 vdd.n1057 99.5127
R3106 vdd.n2521 vdd.n1048 99.5127
R3107 vdd.n2529 vdd.n1048 99.5127
R3108 vdd.n2529 vdd.n1046 99.5127
R3109 vdd.n2533 vdd.n1046 99.5127
R3110 vdd.n2533 vdd.n1036 99.5127
R3111 vdd.n2541 vdd.n1036 99.5127
R3112 vdd.n2541 vdd.n1034 99.5127
R3113 vdd.n2545 vdd.n1034 99.5127
R3114 vdd.n2545 vdd.n1025 99.5127
R3115 vdd.n2553 vdd.n1025 99.5127
R3116 vdd.n2553 vdd.n1023 99.5127
R3117 vdd.n2557 vdd.n1023 99.5127
R3118 vdd.n2557 vdd.n1014 99.5127
R3119 vdd.n2565 vdd.n1014 99.5127
R3120 vdd.n2565 vdd.n1011 99.5127
R3121 vdd.n2571 vdd.n1011 99.5127
R3122 vdd.n2571 vdd.n1012 99.5127
R3123 vdd.n1012 vdd.n1003 99.5127
R3124 vdd.n1003 vdd.n994 99.5127
R3125 vdd.n2653 vdd.n994 99.5127
R3126 vdd.n9 vdd.n7 98.9633
R3127 vdd.n2 vdd.n0 98.9633
R3128 vdd.n9 vdd.n8 98.6055
R3129 vdd.n11 vdd.n10 98.6055
R3130 vdd.n13 vdd.n12 98.6055
R3131 vdd.n6 vdd.n5 98.6055
R3132 vdd.n4 vdd.n3 98.6055
R3133 vdd.n2 vdd.n1 98.6055
R3134 vdd.t180 vdd.n303 85.8723
R3135 vdd.t221 vdd.n244 85.8723
R3136 vdd.t160 vdd.n201 85.8723
R3137 vdd.t201 vdd.n142 85.8723
R3138 vdd.t244 vdd.n100 85.8723
R3139 vdd.t270 vdd.n41 85.8723
R3140 vdd.t300 vdd.n1802 85.8723
R3141 vdd.t249 vdd.n1861 85.8723
R3142 vdd.t288 vdd.n1700 85.8723
R3143 vdd.t237 vdd.n1759 85.8723
R3144 vdd.t241 vdd.n1599 85.8723
R3145 vdd.t246 vdd.n1658 85.8723
R3146 vdd.n3080 vdd.n885 78.546
R3147 vdd.n2519 vdd.n1058 78.546
R3148 vdd.n290 vdd.n289 75.1835
R3149 vdd.n288 vdd.n287 75.1835
R3150 vdd.n286 vdd.n285 75.1835
R3151 vdd.n284 vdd.n283 75.1835
R3152 vdd.n282 vdd.n281 75.1835
R3153 vdd.n280 vdd.n279 75.1835
R3154 vdd.n278 vdd.n277 75.1835
R3155 vdd.n276 vdd.n275 75.1835
R3156 vdd.n274 vdd.n273 75.1835
R3157 vdd.n188 vdd.n187 75.1835
R3158 vdd.n186 vdd.n185 75.1835
R3159 vdd.n184 vdd.n183 75.1835
R3160 vdd.n182 vdd.n181 75.1835
R3161 vdd.n180 vdd.n179 75.1835
R3162 vdd.n178 vdd.n177 75.1835
R3163 vdd.n176 vdd.n175 75.1835
R3164 vdd.n174 vdd.n173 75.1835
R3165 vdd.n172 vdd.n171 75.1835
R3166 vdd.n87 vdd.n86 75.1835
R3167 vdd.n85 vdd.n84 75.1835
R3168 vdd.n83 vdd.n82 75.1835
R3169 vdd.n81 vdd.n80 75.1835
R3170 vdd.n79 vdd.n78 75.1835
R3171 vdd.n77 vdd.n76 75.1835
R3172 vdd.n75 vdd.n74 75.1835
R3173 vdd.n73 vdd.n72 75.1835
R3174 vdd.n71 vdd.n70 75.1835
R3175 vdd.n1832 vdd.n1831 75.1835
R3176 vdd.n1834 vdd.n1833 75.1835
R3177 vdd.n1836 vdd.n1835 75.1835
R3178 vdd.n1838 vdd.n1837 75.1835
R3179 vdd.n1840 vdd.n1839 75.1835
R3180 vdd.n1842 vdd.n1841 75.1835
R3181 vdd.n1844 vdd.n1843 75.1835
R3182 vdd.n1846 vdd.n1845 75.1835
R3183 vdd.n1848 vdd.n1847 75.1835
R3184 vdd.n1730 vdd.n1729 75.1835
R3185 vdd.n1732 vdd.n1731 75.1835
R3186 vdd.n1734 vdd.n1733 75.1835
R3187 vdd.n1736 vdd.n1735 75.1835
R3188 vdd.n1738 vdd.n1737 75.1835
R3189 vdd.n1740 vdd.n1739 75.1835
R3190 vdd.n1742 vdd.n1741 75.1835
R3191 vdd.n1744 vdd.n1743 75.1835
R3192 vdd.n1746 vdd.n1745 75.1835
R3193 vdd.n1629 vdd.n1628 75.1835
R3194 vdd.n1631 vdd.n1630 75.1835
R3195 vdd.n1633 vdd.n1632 75.1835
R3196 vdd.n1635 vdd.n1634 75.1835
R3197 vdd.n1637 vdd.n1636 75.1835
R3198 vdd.n1639 vdd.n1638 75.1835
R3199 vdd.n1641 vdd.n1640 75.1835
R3200 vdd.n1643 vdd.n1642 75.1835
R3201 vdd.n1645 vdd.n1644 75.1835
R3202 vdd.n3010 vdd.n2743 72.8958
R3203 vdd.n3010 vdd.n2744 72.8958
R3204 vdd.n3010 vdd.n2745 72.8958
R3205 vdd.n3010 vdd.n2746 72.8958
R3206 vdd.n3010 vdd.n2747 72.8958
R3207 vdd.n3010 vdd.n2748 72.8958
R3208 vdd.n3010 vdd.n2749 72.8958
R3209 vdd.n3010 vdd.n2750 72.8958
R3210 vdd.n3010 vdd.n2751 72.8958
R3211 vdd.n3010 vdd.n2752 72.8958
R3212 vdd.n3010 vdd.n2753 72.8958
R3213 vdd.n3010 vdd.n2754 72.8958
R3214 vdd.n3010 vdd.n2755 72.8958
R3215 vdd.n3010 vdd.n2756 72.8958
R3216 vdd.n3010 vdd.n2757 72.8958
R3217 vdd.n3010 vdd.n2758 72.8958
R3218 vdd.n3010 vdd.n2759 72.8958
R3219 vdd.n803 vdd.n692 72.8958
R3220 vdd.n3248 vdd.n692 72.8958
R3221 vdd.n797 vdd.n692 72.8958
R3222 vdd.n3255 vdd.n692 72.8958
R3223 vdd.n794 vdd.n692 72.8958
R3224 vdd.n3262 vdd.n692 72.8958
R3225 vdd.n791 vdd.n692 72.8958
R3226 vdd.n3269 vdd.n692 72.8958
R3227 vdd.n3272 vdd.n692 72.8958
R3228 vdd.n3128 vdd.n692 72.8958
R3229 vdd.n3133 vdd.n692 72.8958
R3230 vdd.n3127 vdd.n692 72.8958
R3231 vdd.n3140 vdd.n692 72.8958
R3232 vdd.n3124 vdd.n692 72.8958
R3233 vdd.n3147 vdd.n692 72.8958
R3234 vdd.n3121 vdd.n692 72.8958
R3235 vdd.n3154 vdd.n692 72.8958
R3236 vdd.n2461 vdd.n1110 72.8958
R3237 vdd.n1115 vdd.n1110 72.8958
R3238 vdd.n2454 vdd.n1110 72.8958
R3239 vdd.n2448 vdd.n1110 72.8958
R3240 vdd.n2446 vdd.n1110 72.8958
R3241 vdd.n2440 vdd.n1110 72.8958
R3242 vdd.n2438 vdd.n1110 72.8958
R3243 vdd.n2432 vdd.n1110 72.8958
R3244 vdd.n2430 vdd.n1110 72.8958
R3245 vdd.n2424 vdd.n1110 72.8958
R3246 vdd.n2422 vdd.n1110 72.8958
R3247 vdd.n2416 vdd.n1110 72.8958
R3248 vdd.n2414 vdd.n1110 72.8958
R3249 vdd.n2408 vdd.n1110 72.8958
R3250 vdd.n2406 vdd.n1110 72.8958
R3251 vdd.n2399 vdd.n1110 72.8958
R3252 vdd.n2397 vdd.n1110 72.8958
R3253 vdd.n2726 vdd.n968 72.8958
R3254 vdd.n2726 vdd.n969 72.8958
R3255 vdd.n2726 vdd.n970 72.8958
R3256 vdd.n2726 vdd.n971 72.8958
R3257 vdd.n2726 vdd.n972 72.8958
R3258 vdd.n2726 vdd.n973 72.8958
R3259 vdd.n2726 vdd.n974 72.8958
R3260 vdd.n2726 vdd.n975 72.8958
R3261 vdd.n2726 vdd.n976 72.8958
R3262 vdd.n2726 vdd.n977 72.8958
R3263 vdd.n2726 vdd.n978 72.8958
R3264 vdd.n2726 vdd.n979 72.8958
R3265 vdd.n2726 vdd.n980 72.8958
R3266 vdd.n2726 vdd.n981 72.8958
R3267 vdd.n2726 vdd.n982 72.8958
R3268 vdd.n2726 vdd.n983 72.8958
R3269 vdd.n2726 vdd.n984 72.8958
R3270 vdd.n3011 vdd.n3010 72.8958
R3271 vdd.n3010 vdd.n2727 72.8958
R3272 vdd.n3010 vdd.n2728 72.8958
R3273 vdd.n3010 vdd.n2729 72.8958
R3274 vdd.n3010 vdd.n2730 72.8958
R3275 vdd.n3010 vdd.n2731 72.8958
R3276 vdd.n3010 vdd.n2732 72.8958
R3277 vdd.n3010 vdd.n2733 72.8958
R3278 vdd.n3010 vdd.n2734 72.8958
R3279 vdd.n3010 vdd.n2735 72.8958
R3280 vdd.n3010 vdd.n2736 72.8958
R3281 vdd.n3010 vdd.n2737 72.8958
R3282 vdd.n3010 vdd.n2738 72.8958
R3283 vdd.n3010 vdd.n2739 72.8958
R3284 vdd.n3010 vdd.n2740 72.8958
R3285 vdd.n3010 vdd.n2741 72.8958
R3286 vdd.n3010 vdd.n2742 72.8958
R3287 vdd.n3178 vdd.n692 72.8958
R3288 vdd.n835 vdd.n692 72.8958
R3289 vdd.n3186 vdd.n692 72.8958
R3290 vdd.n830 vdd.n692 72.8958
R3291 vdd.n3193 vdd.n692 72.8958
R3292 vdd.n827 vdd.n692 72.8958
R3293 vdd.n3200 vdd.n692 72.8958
R3294 vdd.n824 vdd.n692 72.8958
R3295 vdd.n3207 vdd.n692 72.8958
R3296 vdd.n3211 vdd.n692 72.8958
R3297 vdd.n821 vdd.n692 72.8958
R3298 vdd.n3218 vdd.n692 72.8958
R3299 vdd.n818 vdd.n692 72.8958
R3300 vdd.n3225 vdd.n692 72.8958
R3301 vdd.n815 vdd.n692 72.8958
R3302 vdd.n3232 vdd.n692 72.8958
R3303 vdd.n3235 vdd.n692 72.8958
R3304 vdd.n2726 vdd.n966 72.8958
R3305 vdd.n2726 vdd.n965 72.8958
R3306 vdd.n2726 vdd.n964 72.8958
R3307 vdd.n2726 vdd.n963 72.8958
R3308 vdd.n2726 vdd.n962 72.8958
R3309 vdd.n2726 vdd.n961 72.8958
R3310 vdd.n2726 vdd.n960 72.8958
R3311 vdd.n2726 vdd.n959 72.8958
R3312 vdd.n2726 vdd.n958 72.8958
R3313 vdd.n2726 vdd.n957 72.8958
R3314 vdd.n2726 vdd.n956 72.8958
R3315 vdd.n2726 vdd.n955 72.8958
R3316 vdd.n2726 vdd.n954 72.8958
R3317 vdd.n2726 vdd.n953 72.8958
R3318 vdd.n2726 vdd.n952 72.8958
R3319 vdd.n2726 vdd.n951 72.8958
R3320 vdd.n2726 vdd.n950 72.8958
R3321 vdd.n2215 vdd.n1110 72.8958
R3322 vdd.n2217 vdd.n1110 72.8958
R3323 vdd.n2223 vdd.n1110 72.8958
R3324 vdd.n2225 vdd.n1110 72.8958
R3325 vdd.n2231 vdd.n1110 72.8958
R3326 vdd.n2233 vdd.n1110 72.8958
R3327 vdd.n2239 vdd.n1110 72.8958
R3328 vdd.n2241 vdd.n1110 72.8958
R3329 vdd.n2247 vdd.n1110 72.8958
R3330 vdd.n2249 vdd.n1110 72.8958
R3331 vdd.n2255 vdd.n1110 72.8958
R3332 vdd.n2257 vdd.n1110 72.8958
R3333 vdd.n2263 vdd.n1110 72.8958
R3334 vdd.n2265 vdd.n1110 72.8958
R3335 vdd.n2271 vdd.n1110 72.8958
R3336 vdd.n2273 vdd.n1110 72.8958
R3337 vdd.n2280 vdd.n1110 72.8958
R3338 vdd.n1499 vdd.n1498 66.2847
R3339 vdd.n1498 vdd.n1274 66.2847
R3340 vdd.n1498 vdd.n1275 66.2847
R3341 vdd.n1498 vdd.n1276 66.2847
R3342 vdd.n1498 vdd.n1277 66.2847
R3343 vdd.n1498 vdd.n1278 66.2847
R3344 vdd.n1498 vdd.n1279 66.2847
R3345 vdd.n1498 vdd.n1280 66.2847
R3346 vdd.n1498 vdd.n1281 66.2847
R3347 vdd.n1498 vdd.n1282 66.2847
R3348 vdd.n1498 vdd.n1283 66.2847
R3349 vdd.n1498 vdd.n1284 66.2847
R3350 vdd.n1498 vdd.n1285 66.2847
R3351 vdd.n1498 vdd.n1286 66.2847
R3352 vdd.n1498 vdd.n1287 66.2847
R3353 vdd.n1498 vdd.n1288 66.2847
R3354 vdd.n1498 vdd.n1289 66.2847
R3355 vdd.n1498 vdd.n1290 66.2847
R3356 vdd.n1498 vdd.n1291 66.2847
R3357 vdd.n1498 vdd.n1292 66.2847
R3358 vdd.n1498 vdd.n1293 66.2847
R3359 vdd.n1498 vdd.n1294 66.2847
R3360 vdd.n1498 vdd.n1295 66.2847
R3361 vdd.n1498 vdd.n1296 66.2847
R3362 vdd.n1498 vdd.n1297 66.2847
R3363 vdd.n1498 vdd.n1298 66.2847
R3364 vdd.n1498 vdd.n1299 66.2847
R3365 vdd.n1498 vdd.n1300 66.2847
R3366 vdd.n1498 vdd.n1301 66.2847
R3367 vdd.n1498 vdd.n1302 66.2847
R3368 vdd.n1498 vdd.n1303 66.2847
R3369 vdd.n1153 vdd.n1150 66.2847
R3370 vdd.n2080 vdd.n1153 66.2847
R3371 vdd.n2085 vdd.n1153 66.2847
R3372 vdd.n2090 vdd.n1153 66.2847
R3373 vdd.n2078 vdd.n1153 66.2847
R3374 vdd.n2097 vdd.n1153 66.2847
R3375 vdd.n2070 vdd.n1153 66.2847
R3376 vdd.n2104 vdd.n1153 66.2847
R3377 vdd.n2063 vdd.n1153 66.2847
R3378 vdd.n2111 vdd.n1153 66.2847
R3379 vdd.n2057 vdd.n1153 66.2847
R3380 vdd.n2052 vdd.n1153 66.2847
R3381 vdd.n2122 vdd.n1153 66.2847
R3382 vdd.n2044 vdd.n1153 66.2847
R3383 vdd.n2129 vdd.n1153 66.2847
R3384 vdd.n2037 vdd.n1153 66.2847
R3385 vdd.n2136 vdd.n1153 66.2847
R3386 vdd.n2030 vdd.n1153 66.2847
R3387 vdd.n2143 vdd.n1153 66.2847
R3388 vdd.n2023 vdd.n1153 66.2847
R3389 vdd.n2150 vdd.n1153 66.2847
R3390 vdd.n2017 vdd.n1153 66.2847
R3391 vdd.n2012 vdd.n1153 66.2847
R3392 vdd.n2161 vdd.n1153 66.2847
R3393 vdd.n2004 vdd.n1153 66.2847
R3394 vdd.n2168 vdd.n1153 66.2847
R3395 vdd.n1997 vdd.n1153 66.2847
R3396 vdd.n2175 vdd.n1153 66.2847
R3397 vdd.n2178 vdd.n1153 66.2847
R3398 vdd.n1988 vdd.n1153 66.2847
R3399 vdd.n2187 vdd.n1153 66.2847
R3400 vdd.n1982 vdd.n1153 66.2847
R3401 vdd.n3405 vdd.n3404 66.2847
R3402 vdd.n3405 vdd.n693 66.2847
R3403 vdd.n3405 vdd.n694 66.2847
R3404 vdd.n3405 vdd.n695 66.2847
R3405 vdd.n3405 vdd.n696 66.2847
R3406 vdd.n3405 vdd.n697 66.2847
R3407 vdd.n3405 vdd.n698 66.2847
R3408 vdd.n3405 vdd.n699 66.2847
R3409 vdd.n3405 vdd.n700 66.2847
R3410 vdd.n3405 vdd.n701 66.2847
R3411 vdd.n3405 vdd.n702 66.2847
R3412 vdd.n3405 vdd.n703 66.2847
R3413 vdd.n3405 vdd.n704 66.2847
R3414 vdd.n3405 vdd.n705 66.2847
R3415 vdd.n3405 vdd.n706 66.2847
R3416 vdd.n3405 vdd.n707 66.2847
R3417 vdd.n3405 vdd.n708 66.2847
R3418 vdd.n3405 vdd.n709 66.2847
R3419 vdd.n3405 vdd.n710 66.2847
R3420 vdd.n3405 vdd.n711 66.2847
R3421 vdd.n3405 vdd.n712 66.2847
R3422 vdd.n3405 vdd.n713 66.2847
R3423 vdd.n3405 vdd.n714 66.2847
R3424 vdd.n3405 vdd.n715 66.2847
R3425 vdd.n3405 vdd.n716 66.2847
R3426 vdd.n3405 vdd.n717 66.2847
R3427 vdd.n3405 vdd.n718 66.2847
R3428 vdd.n3405 vdd.n719 66.2847
R3429 vdd.n3405 vdd.n720 66.2847
R3430 vdd.n3405 vdd.n721 66.2847
R3431 vdd.n3405 vdd.n722 66.2847
R3432 vdd.n3536 vdd.n3535 66.2847
R3433 vdd.n3536 vdd.n424 66.2847
R3434 vdd.n3536 vdd.n423 66.2847
R3435 vdd.n3536 vdd.n422 66.2847
R3436 vdd.n3536 vdd.n421 66.2847
R3437 vdd.n3536 vdd.n420 66.2847
R3438 vdd.n3536 vdd.n419 66.2847
R3439 vdd.n3536 vdd.n418 66.2847
R3440 vdd.n3536 vdd.n417 66.2847
R3441 vdd.n3536 vdd.n416 66.2847
R3442 vdd.n3536 vdd.n415 66.2847
R3443 vdd.n3536 vdd.n414 66.2847
R3444 vdd.n3536 vdd.n413 66.2847
R3445 vdd.n3536 vdd.n412 66.2847
R3446 vdd.n3536 vdd.n411 66.2847
R3447 vdd.n3536 vdd.n410 66.2847
R3448 vdd.n3536 vdd.n409 66.2847
R3449 vdd.n3536 vdd.n408 66.2847
R3450 vdd.n3536 vdd.n407 66.2847
R3451 vdd.n3536 vdd.n406 66.2847
R3452 vdd.n3536 vdd.n405 66.2847
R3453 vdd.n3536 vdd.n404 66.2847
R3454 vdd.n3536 vdd.n403 66.2847
R3455 vdd.n3536 vdd.n402 66.2847
R3456 vdd.n3536 vdd.n401 66.2847
R3457 vdd.n3536 vdd.n400 66.2847
R3458 vdd.n3536 vdd.n399 66.2847
R3459 vdd.n3536 vdd.n398 66.2847
R3460 vdd.n3536 vdd.n397 66.2847
R3461 vdd.n3536 vdd.n396 66.2847
R3462 vdd.n3536 vdd.n395 66.2847
R3463 vdd.n3536 vdd.n394 66.2847
R3464 vdd.n467 vdd.n394 52.4337
R3465 vdd.n473 vdd.n395 52.4337
R3466 vdd.n477 vdd.n396 52.4337
R3467 vdd.n483 vdd.n397 52.4337
R3468 vdd.n487 vdd.n398 52.4337
R3469 vdd.n493 vdd.n399 52.4337
R3470 vdd.n497 vdd.n400 52.4337
R3471 vdd.n503 vdd.n401 52.4337
R3472 vdd.n507 vdd.n402 52.4337
R3473 vdd.n513 vdd.n403 52.4337
R3474 vdd.n517 vdd.n404 52.4337
R3475 vdd.n523 vdd.n405 52.4337
R3476 vdd.n527 vdd.n406 52.4337
R3477 vdd.n533 vdd.n407 52.4337
R3478 vdd.n537 vdd.n408 52.4337
R3479 vdd.n543 vdd.n409 52.4337
R3480 vdd.n547 vdd.n410 52.4337
R3481 vdd.n553 vdd.n411 52.4337
R3482 vdd.n557 vdd.n412 52.4337
R3483 vdd.n563 vdd.n413 52.4337
R3484 vdd.n567 vdd.n414 52.4337
R3485 vdd.n573 vdd.n415 52.4337
R3486 vdd.n577 vdd.n416 52.4337
R3487 vdd.n583 vdd.n417 52.4337
R3488 vdd.n587 vdd.n418 52.4337
R3489 vdd.n593 vdd.n419 52.4337
R3490 vdd.n597 vdd.n420 52.4337
R3491 vdd.n603 vdd.n421 52.4337
R3492 vdd.n607 vdd.n422 52.4337
R3493 vdd.n613 vdd.n423 52.4337
R3494 vdd.n616 vdd.n424 52.4337
R3495 vdd.n3535 vdd.n3534 52.4337
R3496 vdd.n3404 vdd.n3403 52.4337
R3497 vdd.n728 vdd.n693 52.4337
R3498 vdd.n734 vdd.n694 52.4337
R3499 vdd.n3393 vdd.n695 52.4337
R3500 vdd.n3389 vdd.n696 52.4337
R3501 vdd.n3385 vdd.n697 52.4337
R3502 vdd.n3381 vdd.n698 52.4337
R3503 vdd.n3377 vdd.n699 52.4337
R3504 vdd.n3373 vdd.n700 52.4337
R3505 vdd.n3369 vdd.n701 52.4337
R3506 vdd.n3361 vdd.n702 52.4337
R3507 vdd.n3357 vdd.n703 52.4337
R3508 vdd.n3353 vdd.n704 52.4337
R3509 vdd.n3349 vdd.n705 52.4337
R3510 vdd.n3345 vdd.n706 52.4337
R3511 vdd.n3341 vdd.n707 52.4337
R3512 vdd.n3337 vdd.n708 52.4337
R3513 vdd.n3333 vdd.n709 52.4337
R3514 vdd.n3329 vdd.n710 52.4337
R3515 vdd.n3325 vdd.n711 52.4337
R3516 vdd.n3321 vdd.n712 52.4337
R3517 vdd.n3315 vdd.n713 52.4337
R3518 vdd.n3311 vdd.n714 52.4337
R3519 vdd.n3307 vdd.n715 52.4337
R3520 vdd.n3303 vdd.n716 52.4337
R3521 vdd.n3299 vdd.n717 52.4337
R3522 vdd.n3295 vdd.n718 52.4337
R3523 vdd.n3291 vdd.n719 52.4337
R3524 vdd.n3287 vdd.n720 52.4337
R3525 vdd.n3283 vdd.n721 52.4337
R3526 vdd.n3279 vdd.n722 52.4337
R3527 vdd.n2189 vdd.n1982 52.4337
R3528 vdd.n2187 vdd.n2186 52.4337
R3529 vdd.n1989 vdd.n1988 52.4337
R3530 vdd.n2178 vdd.n2177 52.4337
R3531 vdd.n2175 vdd.n2174 52.4337
R3532 vdd.n2170 vdd.n1997 52.4337
R3533 vdd.n2168 vdd.n2167 52.4337
R3534 vdd.n2163 vdd.n2004 52.4337
R3535 vdd.n2161 vdd.n2160 52.4337
R3536 vdd.n2013 vdd.n2012 52.4337
R3537 vdd.n2152 vdd.n2017 52.4337
R3538 vdd.n2150 vdd.n2149 52.4337
R3539 vdd.n2145 vdd.n2023 52.4337
R3540 vdd.n2143 vdd.n2142 52.4337
R3541 vdd.n2138 vdd.n2030 52.4337
R3542 vdd.n2136 vdd.n2135 52.4337
R3543 vdd.n2131 vdd.n2037 52.4337
R3544 vdd.n2129 vdd.n2128 52.4337
R3545 vdd.n2124 vdd.n2044 52.4337
R3546 vdd.n2122 vdd.n2121 52.4337
R3547 vdd.n2053 vdd.n2052 52.4337
R3548 vdd.n2113 vdd.n2057 52.4337
R3549 vdd.n2111 vdd.n2110 52.4337
R3550 vdd.n2106 vdd.n2063 52.4337
R3551 vdd.n2104 vdd.n2103 52.4337
R3552 vdd.n2099 vdd.n2070 52.4337
R3553 vdd.n2097 vdd.n2096 52.4337
R3554 vdd.n2092 vdd.n2078 52.4337
R3555 vdd.n2090 vdd.n2089 52.4337
R3556 vdd.n2085 vdd.n2084 52.4337
R3557 vdd.n2080 vdd.n2079 52.4337
R3558 vdd.n2198 vdd.n1150 52.4337
R3559 vdd.n1500 vdd.n1499 52.4337
R3560 vdd.n1306 vdd.n1274 52.4337
R3561 vdd.n1310 vdd.n1275 52.4337
R3562 vdd.n1312 vdd.n1276 52.4337
R3563 vdd.n1316 vdd.n1277 52.4337
R3564 vdd.n1318 vdd.n1278 52.4337
R3565 vdd.n1322 vdd.n1279 52.4337
R3566 vdd.n1324 vdd.n1280 52.4337
R3567 vdd.n1328 vdd.n1281 52.4337
R3568 vdd.n1330 vdd.n1282 52.4337
R3569 vdd.n1336 vdd.n1283 52.4337
R3570 vdd.n1338 vdd.n1284 52.4337
R3571 vdd.n1342 vdd.n1285 52.4337
R3572 vdd.n1344 vdd.n1286 52.4337
R3573 vdd.n1348 vdd.n1287 52.4337
R3574 vdd.n1350 vdd.n1288 52.4337
R3575 vdd.n1354 vdd.n1289 52.4337
R3576 vdd.n1356 vdd.n1290 52.4337
R3577 vdd.n1360 vdd.n1291 52.4337
R3578 vdd.n1362 vdd.n1292 52.4337
R3579 vdd.n1434 vdd.n1293 52.4337
R3580 vdd.n1367 vdd.n1294 52.4337
R3581 vdd.n1371 vdd.n1295 52.4337
R3582 vdd.n1373 vdd.n1296 52.4337
R3583 vdd.n1377 vdd.n1297 52.4337
R3584 vdd.n1379 vdd.n1298 52.4337
R3585 vdd.n1383 vdd.n1299 52.4337
R3586 vdd.n1385 vdd.n1300 52.4337
R3587 vdd.n1389 vdd.n1301 52.4337
R3588 vdd.n1391 vdd.n1302 52.4337
R3589 vdd.n1395 vdd.n1303 52.4337
R3590 vdd.n1499 vdd.n1273 52.4337
R3591 vdd.n1309 vdd.n1274 52.4337
R3592 vdd.n1311 vdd.n1275 52.4337
R3593 vdd.n1315 vdd.n1276 52.4337
R3594 vdd.n1317 vdd.n1277 52.4337
R3595 vdd.n1321 vdd.n1278 52.4337
R3596 vdd.n1323 vdd.n1279 52.4337
R3597 vdd.n1327 vdd.n1280 52.4337
R3598 vdd.n1329 vdd.n1281 52.4337
R3599 vdd.n1335 vdd.n1282 52.4337
R3600 vdd.n1337 vdd.n1283 52.4337
R3601 vdd.n1341 vdd.n1284 52.4337
R3602 vdd.n1343 vdd.n1285 52.4337
R3603 vdd.n1347 vdd.n1286 52.4337
R3604 vdd.n1349 vdd.n1287 52.4337
R3605 vdd.n1353 vdd.n1288 52.4337
R3606 vdd.n1355 vdd.n1289 52.4337
R3607 vdd.n1359 vdd.n1290 52.4337
R3608 vdd.n1361 vdd.n1291 52.4337
R3609 vdd.n1365 vdd.n1292 52.4337
R3610 vdd.n1366 vdd.n1293 52.4337
R3611 vdd.n1370 vdd.n1294 52.4337
R3612 vdd.n1372 vdd.n1295 52.4337
R3613 vdd.n1376 vdd.n1296 52.4337
R3614 vdd.n1378 vdd.n1297 52.4337
R3615 vdd.n1382 vdd.n1298 52.4337
R3616 vdd.n1384 vdd.n1299 52.4337
R3617 vdd.n1388 vdd.n1300 52.4337
R3618 vdd.n1390 vdd.n1301 52.4337
R3619 vdd.n1394 vdd.n1302 52.4337
R3620 vdd.n1396 vdd.n1303 52.4337
R3621 vdd.n1150 vdd.n1149 52.4337
R3622 vdd.n2081 vdd.n2080 52.4337
R3623 vdd.n2086 vdd.n2085 52.4337
R3624 vdd.n2091 vdd.n2090 52.4337
R3625 vdd.n2078 vdd.n2071 52.4337
R3626 vdd.n2098 vdd.n2097 52.4337
R3627 vdd.n2070 vdd.n2064 52.4337
R3628 vdd.n2105 vdd.n2104 52.4337
R3629 vdd.n2063 vdd.n2058 52.4337
R3630 vdd.n2112 vdd.n2111 52.4337
R3631 vdd.n2057 vdd.n2056 52.4337
R3632 vdd.n2052 vdd.n2045 52.4337
R3633 vdd.n2123 vdd.n2122 52.4337
R3634 vdd.n2044 vdd.n2038 52.4337
R3635 vdd.n2130 vdd.n2129 52.4337
R3636 vdd.n2037 vdd.n2031 52.4337
R3637 vdd.n2137 vdd.n2136 52.4337
R3638 vdd.n2030 vdd.n2024 52.4337
R3639 vdd.n2144 vdd.n2143 52.4337
R3640 vdd.n2023 vdd.n2018 52.4337
R3641 vdd.n2151 vdd.n2150 52.4337
R3642 vdd.n2017 vdd.n2016 52.4337
R3643 vdd.n2012 vdd.n2005 52.4337
R3644 vdd.n2162 vdd.n2161 52.4337
R3645 vdd.n2004 vdd.n1998 52.4337
R3646 vdd.n2169 vdd.n2168 52.4337
R3647 vdd.n1997 vdd.n1991 52.4337
R3648 vdd.n2176 vdd.n2175 52.4337
R3649 vdd.n2179 vdd.n2178 52.4337
R3650 vdd.n1988 vdd.n1983 52.4337
R3651 vdd.n2188 vdd.n2187 52.4337
R3652 vdd.n1982 vdd.n1155 52.4337
R3653 vdd.n3404 vdd.n725 52.4337
R3654 vdd.n733 vdd.n693 52.4337
R3655 vdd.n3394 vdd.n694 52.4337
R3656 vdd.n3390 vdd.n695 52.4337
R3657 vdd.n3386 vdd.n696 52.4337
R3658 vdd.n3382 vdd.n697 52.4337
R3659 vdd.n3378 vdd.n698 52.4337
R3660 vdd.n3374 vdd.n699 52.4337
R3661 vdd.n3370 vdd.n700 52.4337
R3662 vdd.n3360 vdd.n701 52.4337
R3663 vdd.n3358 vdd.n702 52.4337
R3664 vdd.n3354 vdd.n703 52.4337
R3665 vdd.n3350 vdd.n704 52.4337
R3666 vdd.n3346 vdd.n705 52.4337
R3667 vdd.n3342 vdd.n706 52.4337
R3668 vdd.n3338 vdd.n707 52.4337
R3669 vdd.n3334 vdd.n708 52.4337
R3670 vdd.n3330 vdd.n709 52.4337
R3671 vdd.n3326 vdd.n710 52.4337
R3672 vdd.n3322 vdd.n711 52.4337
R3673 vdd.n3314 vdd.n712 52.4337
R3674 vdd.n3312 vdd.n713 52.4337
R3675 vdd.n3308 vdd.n714 52.4337
R3676 vdd.n3304 vdd.n715 52.4337
R3677 vdd.n3300 vdd.n716 52.4337
R3678 vdd.n3296 vdd.n717 52.4337
R3679 vdd.n3292 vdd.n718 52.4337
R3680 vdd.n3288 vdd.n719 52.4337
R3681 vdd.n3284 vdd.n720 52.4337
R3682 vdd.n3280 vdd.n721 52.4337
R3683 vdd.n722 vdd.n691 52.4337
R3684 vdd.n3535 vdd.n425 52.4337
R3685 vdd.n614 vdd.n424 52.4337
R3686 vdd.n608 vdd.n423 52.4337
R3687 vdd.n604 vdd.n422 52.4337
R3688 vdd.n598 vdd.n421 52.4337
R3689 vdd.n594 vdd.n420 52.4337
R3690 vdd.n588 vdd.n419 52.4337
R3691 vdd.n584 vdd.n418 52.4337
R3692 vdd.n578 vdd.n417 52.4337
R3693 vdd.n574 vdd.n416 52.4337
R3694 vdd.n568 vdd.n415 52.4337
R3695 vdd.n564 vdd.n414 52.4337
R3696 vdd.n558 vdd.n413 52.4337
R3697 vdd.n554 vdd.n412 52.4337
R3698 vdd.n548 vdd.n411 52.4337
R3699 vdd.n544 vdd.n410 52.4337
R3700 vdd.n538 vdd.n409 52.4337
R3701 vdd.n534 vdd.n408 52.4337
R3702 vdd.n528 vdd.n407 52.4337
R3703 vdd.n524 vdd.n406 52.4337
R3704 vdd.n518 vdd.n405 52.4337
R3705 vdd.n514 vdd.n404 52.4337
R3706 vdd.n508 vdd.n403 52.4337
R3707 vdd.n504 vdd.n402 52.4337
R3708 vdd.n498 vdd.n401 52.4337
R3709 vdd.n494 vdd.n400 52.4337
R3710 vdd.n488 vdd.n399 52.4337
R3711 vdd.n484 vdd.n398 52.4337
R3712 vdd.n478 vdd.n397 52.4337
R3713 vdd.n474 vdd.n396 52.4337
R3714 vdd.n468 vdd.n395 52.4337
R3715 vdd.n394 vdd.n392 52.4337
R3716 vdd.t125 vdd.t128 51.4683
R3717 vdd.n274 vdd.n272 42.0461
R3718 vdd.n172 vdd.n170 42.0461
R3719 vdd.n71 vdd.n69 42.0461
R3720 vdd.n1832 vdd.n1830 42.0461
R3721 vdd.n1730 vdd.n1728 42.0461
R3722 vdd.n1629 vdd.n1627 42.0461
R3723 vdd.n332 vdd.n331 41.6884
R3724 vdd.n230 vdd.n229 41.6884
R3725 vdd.n129 vdd.n128 41.6884
R3726 vdd.n1890 vdd.n1889 41.6884
R3727 vdd.n1788 vdd.n1787 41.6884
R3728 vdd.n1687 vdd.n1686 41.6884
R3729 vdd.n1399 vdd.n1398 41.1157
R3730 vdd.n1437 vdd.n1436 41.1157
R3731 vdd.n1333 vdd.n1332 41.1157
R3732 vdd.n428 vdd.n427 41.1157
R3733 vdd.n566 vdd.n441 41.1157
R3734 vdd.n454 vdd.n453 41.1157
R3735 vdd.n3235 vdd.n3234 39.2114
R3736 vdd.n3232 vdd.n3231 39.2114
R3737 vdd.n3227 vdd.n815 39.2114
R3738 vdd.n3225 vdd.n3224 39.2114
R3739 vdd.n3220 vdd.n818 39.2114
R3740 vdd.n3218 vdd.n3217 39.2114
R3741 vdd.n3213 vdd.n821 39.2114
R3742 vdd.n3211 vdd.n3210 39.2114
R3743 vdd.n3207 vdd.n3206 39.2114
R3744 vdd.n3202 vdd.n824 39.2114
R3745 vdd.n3200 vdd.n3199 39.2114
R3746 vdd.n3195 vdd.n827 39.2114
R3747 vdd.n3193 vdd.n3192 39.2114
R3748 vdd.n3188 vdd.n830 39.2114
R3749 vdd.n3186 vdd.n3185 39.2114
R3750 vdd.n3180 vdd.n835 39.2114
R3751 vdd.n3178 vdd.n3177 39.2114
R3752 vdd.n3011 vdd.n947 39.2114
R3753 vdd.n2832 vdd.n2727 39.2114
R3754 vdd.n2836 vdd.n2728 39.2114
R3755 vdd.n2840 vdd.n2729 39.2114
R3756 vdd.n2844 vdd.n2730 39.2114
R3757 vdd.n2848 vdd.n2731 39.2114
R3758 vdd.n2852 vdd.n2732 39.2114
R3759 vdd.n2856 vdd.n2733 39.2114
R3760 vdd.n2860 vdd.n2734 39.2114
R3761 vdd.n2864 vdd.n2735 39.2114
R3762 vdd.n2868 vdd.n2736 39.2114
R3763 vdd.n2872 vdd.n2737 39.2114
R3764 vdd.n2876 vdd.n2738 39.2114
R3765 vdd.n2880 vdd.n2739 39.2114
R3766 vdd.n2884 vdd.n2740 39.2114
R3767 vdd.n2888 vdd.n2741 39.2114
R3768 vdd.n2893 vdd.n2742 39.2114
R3769 vdd.n2721 vdd.n984 39.2114
R3770 vdd.n2717 vdd.n983 39.2114
R3771 vdd.n2713 vdd.n982 39.2114
R3772 vdd.n2709 vdd.n981 39.2114
R3773 vdd.n2705 vdd.n980 39.2114
R3774 vdd.n2701 vdd.n979 39.2114
R3775 vdd.n2697 vdd.n978 39.2114
R3776 vdd.n2693 vdd.n977 39.2114
R3777 vdd.n2689 vdd.n976 39.2114
R3778 vdd.n2685 vdd.n975 39.2114
R3779 vdd.n2681 vdd.n974 39.2114
R3780 vdd.n2677 vdd.n973 39.2114
R3781 vdd.n2673 vdd.n972 39.2114
R3782 vdd.n2669 vdd.n971 39.2114
R3783 vdd.n2665 vdd.n970 39.2114
R3784 vdd.n2660 vdd.n969 39.2114
R3785 vdd.n2656 vdd.n968 39.2114
R3786 vdd.n2461 vdd.n1113 39.2114
R3787 vdd.n2459 vdd.n1115 39.2114
R3788 vdd.n2455 vdd.n2454 39.2114
R3789 vdd.n2448 vdd.n1117 39.2114
R3790 vdd.n2447 vdd.n2446 39.2114
R3791 vdd.n2440 vdd.n1119 39.2114
R3792 vdd.n2439 vdd.n2438 39.2114
R3793 vdd.n2432 vdd.n1121 39.2114
R3794 vdd.n2431 vdd.n2430 39.2114
R3795 vdd.n2424 vdd.n1123 39.2114
R3796 vdd.n2423 vdd.n2422 39.2114
R3797 vdd.n2416 vdd.n1125 39.2114
R3798 vdd.n2415 vdd.n2414 39.2114
R3799 vdd.n2408 vdd.n1127 39.2114
R3800 vdd.n2407 vdd.n2406 39.2114
R3801 vdd.n2399 vdd.n1129 39.2114
R3802 vdd.n2398 vdd.n2397 39.2114
R3803 vdd.n3154 vdd.n3153 39.2114
R3804 vdd.n3149 vdd.n3121 39.2114
R3805 vdd.n3147 vdd.n3146 39.2114
R3806 vdd.n3142 vdd.n3124 39.2114
R3807 vdd.n3140 vdd.n3139 39.2114
R3808 vdd.n3135 vdd.n3127 39.2114
R3809 vdd.n3133 vdd.n3132 39.2114
R3810 vdd.n3128 vdd.n787 39.2114
R3811 vdd.n3272 vdd.n3271 39.2114
R3812 vdd.n3269 vdd.n3268 39.2114
R3813 vdd.n3264 vdd.n791 39.2114
R3814 vdd.n3262 vdd.n3261 39.2114
R3815 vdd.n3257 vdd.n794 39.2114
R3816 vdd.n3255 vdd.n3254 39.2114
R3817 vdd.n3250 vdd.n797 39.2114
R3818 vdd.n3248 vdd.n3247 39.2114
R3819 vdd.n3243 vdd.n803 39.2114
R3820 vdd.n2743 vdd.n943 39.2114
R3821 vdd.n2766 vdd.n2744 39.2114
R3822 vdd.n2770 vdd.n2745 39.2114
R3823 vdd.n2774 vdd.n2746 39.2114
R3824 vdd.n2778 vdd.n2747 39.2114
R3825 vdd.n2782 vdd.n2748 39.2114
R3826 vdd.n2786 vdd.n2749 39.2114
R3827 vdd.n2790 vdd.n2750 39.2114
R3828 vdd.n2794 vdd.n2751 39.2114
R3829 vdd.n2798 vdd.n2752 39.2114
R3830 vdd.n2802 vdd.n2753 39.2114
R3831 vdd.n2806 vdd.n2754 39.2114
R3832 vdd.n2810 vdd.n2755 39.2114
R3833 vdd.n2814 vdd.n2756 39.2114
R3834 vdd.n2818 vdd.n2757 39.2114
R3835 vdd.n2822 vdd.n2758 39.2114
R3836 vdd.n2826 vdd.n2759 39.2114
R3837 vdd.n2765 vdd.n2743 39.2114
R3838 vdd.n2769 vdd.n2744 39.2114
R3839 vdd.n2773 vdd.n2745 39.2114
R3840 vdd.n2777 vdd.n2746 39.2114
R3841 vdd.n2781 vdd.n2747 39.2114
R3842 vdd.n2785 vdd.n2748 39.2114
R3843 vdd.n2789 vdd.n2749 39.2114
R3844 vdd.n2793 vdd.n2750 39.2114
R3845 vdd.n2797 vdd.n2751 39.2114
R3846 vdd.n2801 vdd.n2752 39.2114
R3847 vdd.n2805 vdd.n2753 39.2114
R3848 vdd.n2809 vdd.n2754 39.2114
R3849 vdd.n2813 vdd.n2755 39.2114
R3850 vdd.n2817 vdd.n2756 39.2114
R3851 vdd.n2821 vdd.n2757 39.2114
R3852 vdd.n2825 vdd.n2758 39.2114
R3853 vdd.n2760 vdd.n2759 39.2114
R3854 vdd.n803 vdd.n798 39.2114
R3855 vdd.n3249 vdd.n3248 39.2114
R3856 vdd.n797 vdd.n795 39.2114
R3857 vdd.n3256 vdd.n3255 39.2114
R3858 vdd.n794 vdd.n792 39.2114
R3859 vdd.n3263 vdd.n3262 39.2114
R3860 vdd.n791 vdd.n789 39.2114
R3861 vdd.n3270 vdd.n3269 39.2114
R3862 vdd.n3273 vdd.n3272 39.2114
R3863 vdd.n3129 vdd.n3128 39.2114
R3864 vdd.n3134 vdd.n3133 39.2114
R3865 vdd.n3127 vdd.n3125 39.2114
R3866 vdd.n3141 vdd.n3140 39.2114
R3867 vdd.n3124 vdd.n3122 39.2114
R3868 vdd.n3148 vdd.n3147 39.2114
R3869 vdd.n3121 vdd.n3119 39.2114
R3870 vdd.n3155 vdd.n3154 39.2114
R3871 vdd.n2462 vdd.n2461 39.2114
R3872 vdd.n2456 vdd.n1115 39.2114
R3873 vdd.n2454 vdd.n2453 39.2114
R3874 vdd.n2449 vdd.n2448 39.2114
R3875 vdd.n2446 vdd.n2445 39.2114
R3876 vdd.n2441 vdd.n2440 39.2114
R3877 vdd.n2438 vdd.n2437 39.2114
R3878 vdd.n2433 vdd.n2432 39.2114
R3879 vdd.n2430 vdd.n2429 39.2114
R3880 vdd.n2425 vdd.n2424 39.2114
R3881 vdd.n2422 vdd.n2421 39.2114
R3882 vdd.n2417 vdd.n2416 39.2114
R3883 vdd.n2414 vdd.n2413 39.2114
R3884 vdd.n2409 vdd.n2408 39.2114
R3885 vdd.n2406 vdd.n2405 39.2114
R3886 vdd.n2400 vdd.n2399 39.2114
R3887 vdd.n2397 vdd.n2396 39.2114
R3888 vdd.n2659 vdd.n968 39.2114
R3889 vdd.n2664 vdd.n969 39.2114
R3890 vdd.n2668 vdd.n970 39.2114
R3891 vdd.n2672 vdd.n971 39.2114
R3892 vdd.n2676 vdd.n972 39.2114
R3893 vdd.n2680 vdd.n973 39.2114
R3894 vdd.n2684 vdd.n974 39.2114
R3895 vdd.n2688 vdd.n975 39.2114
R3896 vdd.n2692 vdd.n976 39.2114
R3897 vdd.n2696 vdd.n977 39.2114
R3898 vdd.n2700 vdd.n978 39.2114
R3899 vdd.n2704 vdd.n979 39.2114
R3900 vdd.n2708 vdd.n980 39.2114
R3901 vdd.n2712 vdd.n981 39.2114
R3902 vdd.n2716 vdd.n982 39.2114
R3903 vdd.n2720 vdd.n983 39.2114
R3904 vdd.n986 vdd.n984 39.2114
R3905 vdd.n3012 vdd.n3011 39.2114
R3906 vdd.n2835 vdd.n2727 39.2114
R3907 vdd.n2839 vdd.n2728 39.2114
R3908 vdd.n2843 vdd.n2729 39.2114
R3909 vdd.n2847 vdd.n2730 39.2114
R3910 vdd.n2851 vdd.n2731 39.2114
R3911 vdd.n2855 vdd.n2732 39.2114
R3912 vdd.n2859 vdd.n2733 39.2114
R3913 vdd.n2863 vdd.n2734 39.2114
R3914 vdd.n2867 vdd.n2735 39.2114
R3915 vdd.n2871 vdd.n2736 39.2114
R3916 vdd.n2875 vdd.n2737 39.2114
R3917 vdd.n2879 vdd.n2738 39.2114
R3918 vdd.n2883 vdd.n2739 39.2114
R3919 vdd.n2887 vdd.n2740 39.2114
R3920 vdd.n2892 vdd.n2741 39.2114
R3921 vdd.n2895 vdd.n2742 39.2114
R3922 vdd.n3179 vdd.n3178 39.2114
R3923 vdd.n835 vdd.n831 39.2114
R3924 vdd.n3187 vdd.n3186 39.2114
R3925 vdd.n830 vdd.n828 39.2114
R3926 vdd.n3194 vdd.n3193 39.2114
R3927 vdd.n827 vdd.n825 39.2114
R3928 vdd.n3201 vdd.n3200 39.2114
R3929 vdd.n824 vdd.n822 39.2114
R3930 vdd.n3208 vdd.n3207 39.2114
R3931 vdd.n3212 vdd.n3211 39.2114
R3932 vdd.n821 vdd.n819 39.2114
R3933 vdd.n3219 vdd.n3218 39.2114
R3934 vdd.n818 vdd.n816 39.2114
R3935 vdd.n3226 vdd.n3225 39.2114
R3936 vdd.n815 vdd.n813 39.2114
R3937 vdd.n3233 vdd.n3232 39.2114
R3938 vdd.n3236 vdd.n3235 39.2114
R3939 vdd.n995 vdd.n950 39.2114
R3940 vdd.n2648 vdd.n951 39.2114
R3941 vdd.n2644 vdd.n952 39.2114
R3942 vdd.n2640 vdd.n953 39.2114
R3943 vdd.n2636 vdd.n954 39.2114
R3944 vdd.n2632 vdd.n955 39.2114
R3945 vdd.n2628 vdd.n956 39.2114
R3946 vdd.n2624 vdd.n957 39.2114
R3947 vdd.n2620 vdd.n958 39.2114
R3948 vdd.n2616 vdd.n959 39.2114
R3949 vdd.n2612 vdd.n960 39.2114
R3950 vdd.n2608 vdd.n961 39.2114
R3951 vdd.n2604 vdd.n962 39.2114
R3952 vdd.n2600 vdd.n963 39.2114
R3953 vdd.n2596 vdd.n964 39.2114
R3954 vdd.n2592 vdd.n965 39.2114
R3955 vdd.n2588 vdd.n966 39.2114
R3956 vdd.n2215 vdd.n1109 39.2114
R3957 vdd.n2218 vdd.n2217 39.2114
R3958 vdd.n2223 vdd.n2222 39.2114
R3959 vdd.n2226 vdd.n2225 39.2114
R3960 vdd.n2231 vdd.n2230 39.2114
R3961 vdd.n2234 vdd.n2233 39.2114
R3962 vdd.n2239 vdd.n2238 39.2114
R3963 vdd.n2242 vdd.n2241 39.2114
R3964 vdd.n2247 vdd.n2246 39.2114
R3965 vdd.n2250 vdd.n2249 39.2114
R3966 vdd.n2255 vdd.n2254 39.2114
R3967 vdd.n2258 vdd.n2257 39.2114
R3968 vdd.n2263 vdd.n2262 39.2114
R3969 vdd.n2266 vdd.n2265 39.2114
R3970 vdd.n2271 vdd.n2270 39.2114
R3971 vdd.n2274 vdd.n2273 39.2114
R3972 vdd.n2280 vdd.n2279 39.2114
R3973 vdd.n2585 vdd.n966 39.2114
R3974 vdd.n2589 vdd.n965 39.2114
R3975 vdd.n2593 vdd.n964 39.2114
R3976 vdd.n2597 vdd.n963 39.2114
R3977 vdd.n2601 vdd.n962 39.2114
R3978 vdd.n2605 vdd.n961 39.2114
R3979 vdd.n2609 vdd.n960 39.2114
R3980 vdd.n2613 vdd.n959 39.2114
R3981 vdd.n2617 vdd.n958 39.2114
R3982 vdd.n2621 vdd.n957 39.2114
R3983 vdd.n2625 vdd.n956 39.2114
R3984 vdd.n2629 vdd.n955 39.2114
R3985 vdd.n2633 vdd.n954 39.2114
R3986 vdd.n2637 vdd.n953 39.2114
R3987 vdd.n2641 vdd.n952 39.2114
R3988 vdd.n2645 vdd.n951 39.2114
R3989 vdd.n2649 vdd.n950 39.2114
R3990 vdd.n2216 vdd.n2215 39.2114
R3991 vdd.n2217 vdd.n2213 39.2114
R3992 vdd.n2224 vdd.n2223 39.2114
R3993 vdd.n2225 vdd.n2211 39.2114
R3994 vdd.n2232 vdd.n2231 39.2114
R3995 vdd.n2233 vdd.n2209 39.2114
R3996 vdd.n2240 vdd.n2239 39.2114
R3997 vdd.n2241 vdd.n2207 39.2114
R3998 vdd.n2248 vdd.n2247 39.2114
R3999 vdd.n2249 vdd.n1143 39.2114
R4000 vdd.n2256 vdd.n2255 39.2114
R4001 vdd.n2257 vdd.n1141 39.2114
R4002 vdd.n2264 vdd.n2263 39.2114
R4003 vdd.n2265 vdd.n1139 39.2114
R4004 vdd.n2272 vdd.n2271 39.2114
R4005 vdd.n2273 vdd.n1135 39.2114
R4006 vdd.n2281 vdd.n2280 39.2114
R4007 vdd.n2202 vdd.n2201 37.2369
R4008 vdd.n2118 vdd.n2051 37.2369
R4009 vdd.n2157 vdd.n2011 37.2369
R4010 vdd.n3320 vdd.n769 37.2369
R4011 vdd.n3368 vdd.n3367 37.2369
R4012 vdd.n690 vdd.n689 37.2369
R4013 vdd.n2277 vdd.n1137 30.449
R4014 vdd.n999 vdd.n998 30.449
R4015 vdd.n2402 vdd.n1131 30.449
R4016 vdd.n2662 vdd.n989 30.449
R4017 vdd.n2763 vdd.n2762 30.449
R4018 vdd.n3182 vdd.n833 30.449
R4019 vdd.n2890 vdd.n2831 30.449
R4020 vdd.n801 vdd.n800 30.449
R4021 vdd.n2465 vdd.n2464 30.4395
R4022 vdd.n2724 vdd.n987 30.4395
R4023 vdd.n2657 vdd.n990 30.4395
R4024 vdd.n2395 vdd.n2394 30.4395
R4025 vdd.n2897 vdd.n2896 30.4395
R4026 vdd.n3176 vdd.n3175 30.4395
R4027 vdd.n3015 vdd.n3014 30.4395
R4028 vdd.n3239 vdd.n3238 30.4395
R4029 vdd.n3158 vdd.n3157 30.4395
R4030 vdd.n3244 vdd.n802 30.4395
R4031 vdd.n3008 vdd.n3007 30.4395
R4032 vdd.n3019 vdd.n942 30.4395
R4033 vdd.n2469 vdd.n1108 30.4395
R4034 vdd.n2652 vdd.n2651 30.4395
R4035 vdd.n2584 vdd.n2583 30.4395
R4036 vdd.n2284 vdd.n2283 30.4395
R4037 vdd.n1498 vdd.n1305 22.2201
R4038 vdd.n2196 vdd.n1153 22.2201
R4039 vdd.n3405 vdd.n723 22.2201
R4040 vdd.n3537 vdd.n3536 22.2201
R4041 vdd.n1509 vdd.n1267 19.3944
R4042 vdd.n1509 vdd.n1265 19.3944
R4043 vdd.n1513 vdd.n1265 19.3944
R4044 vdd.n1513 vdd.n1255 19.3944
R4045 vdd.n1526 vdd.n1255 19.3944
R4046 vdd.n1526 vdd.n1253 19.3944
R4047 vdd.n1530 vdd.n1253 19.3944
R4048 vdd.n1530 vdd.n1245 19.3944
R4049 vdd.n1543 vdd.n1245 19.3944
R4050 vdd.n1543 vdd.n1243 19.3944
R4051 vdd.n1547 vdd.n1243 19.3944
R4052 vdd.n1547 vdd.n1232 19.3944
R4053 vdd.n1559 vdd.n1232 19.3944
R4054 vdd.n1559 vdd.n1230 19.3944
R4055 vdd.n1563 vdd.n1230 19.3944
R4056 vdd.n1563 vdd.n1221 19.3944
R4057 vdd.n1576 vdd.n1221 19.3944
R4058 vdd.n1576 vdd.n1219 19.3944
R4059 vdd.n1580 vdd.n1219 19.3944
R4060 vdd.n1580 vdd.n1210 19.3944
R4061 vdd.n1899 vdd.n1210 19.3944
R4062 vdd.n1899 vdd.n1208 19.3944
R4063 vdd.n1903 vdd.n1208 19.3944
R4064 vdd.n1903 vdd.n1198 19.3944
R4065 vdd.n1916 vdd.n1198 19.3944
R4066 vdd.n1916 vdd.n1196 19.3944
R4067 vdd.n1920 vdd.n1196 19.3944
R4068 vdd.n1920 vdd.n1188 19.3944
R4069 vdd.n1933 vdd.n1188 19.3944
R4070 vdd.n1933 vdd.n1186 19.3944
R4071 vdd.n1937 vdd.n1186 19.3944
R4072 vdd.n1937 vdd.n1175 19.3944
R4073 vdd.n1949 vdd.n1175 19.3944
R4074 vdd.n1949 vdd.n1173 19.3944
R4075 vdd.n1953 vdd.n1173 19.3944
R4076 vdd.n1953 vdd.n1165 19.3944
R4077 vdd.n1966 vdd.n1165 19.3944
R4078 vdd.n1966 vdd.n1162 19.3944
R4079 vdd.n1972 vdd.n1162 19.3944
R4080 vdd.n1972 vdd.n1163 19.3944
R4081 vdd.n1163 vdd.n1152 19.3944
R4082 vdd.n1433 vdd.n1368 19.3944
R4083 vdd.n1429 vdd.n1368 19.3944
R4084 vdd.n1429 vdd.n1428 19.3944
R4085 vdd.n1428 vdd.n1427 19.3944
R4086 vdd.n1427 vdd.n1374 19.3944
R4087 vdd.n1423 vdd.n1374 19.3944
R4088 vdd.n1423 vdd.n1422 19.3944
R4089 vdd.n1422 vdd.n1421 19.3944
R4090 vdd.n1421 vdd.n1380 19.3944
R4091 vdd.n1417 vdd.n1380 19.3944
R4092 vdd.n1417 vdd.n1416 19.3944
R4093 vdd.n1416 vdd.n1415 19.3944
R4094 vdd.n1415 vdd.n1386 19.3944
R4095 vdd.n1411 vdd.n1386 19.3944
R4096 vdd.n1411 vdd.n1410 19.3944
R4097 vdd.n1410 vdd.n1409 19.3944
R4098 vdd.n1409 vdd.n1392 19.3944
R4099 vdd.n1405 vdd.n1392 19.3944
R4100 vdd.n1405 vdd.n1404 19.3944
R4101 vdd.n1404 vdd.n1403 19.3944
R4102 vdd.n1468 vdd.n1467 19.3944
R4103 vdd.n1467 vdd.n1466 19.3944
R4104 vdd.n1466 vdd.n1339 19.3944
R4105 vdd.n1462 vdd.n1339 19.3944
R4106 vdd.n1462 vdd.n1461 19.3944
R4107 vdd.n1461 vdd.n1460 19.3944
R4108 vdd.n1460 vdd.n1345 19.3944
R4109 vdd.n1456 vdd.n1345 19.3944
R4110 vdd.n1456 vdd.n1455 19.3944
R4111 vdd.n1455 vdd.n1454 19.3944
R4112 vdd.n1454 vdd.n1351 19.3944
R4113 vdd.n1450 vdd.n1351 19.3944
R4114 vdd.n1450 vdd.n1449 19.3944
R4115 vdd.n1449 vdd.n1448 19.3944
R4116 vdd.n1448 vdd.n1357 19.3944
R4117 vdd.n1444 vdd.n1357 19.3944
R4118 vdd.n1444 vdd.n1443 19.3944
R4119 vdd.n1443 vdd.n1442 19.3944
R4120 vdd.n1442 vdd.n1363 19.3944
R4121 vdd.n1438 vdd.n1363 19.3944
R4122 vdd.n1501 vdd.n1272 19.3944
R4123 vdd.n1496 vdd.n1272 19.3944
R4124 vdd.n1496 vdd.n1307 19.3944
R4125 vdd.n1492 vdd.n1307 19.3944
R4126 vdd.n1492 vdd.n1491 19.3944
R4127 vdd.n1491 vdd.n1490 19.3944
R4128 vdd.n1490 vdd.n1313 19.3944
R4129 vdd.n1486 vdd.n1313 19.3944
R4130 vdd.n1486 vdd.n1485 19.3944
R4131 vdd.n1485 vdd.n1484 19.3944
R4132 vdd.n1484 vdd.n1319 19.3944
R4133 vdd.n1480 vdd.n1319 19.3944
R4134 vdd.n1480 vdd.n1479 19.3944
R4135 vdd.n1479 vdd.n1478 19.3944
R4136 vdd.n1478 vdd.n1325 19.3944
R4137 vdd.n1474 vdd.n1325 19.3944
R4138 vdd.n1474 vdd.n1473 19.3944
R4139 vdd.n1473 vdd.n1472 19.3944
R4140 vdd.n2114 vdd.n2049 19.3944
R4141 vdd.n2114 vdd.n2055 19.3944
R4142 vdd.n2109 vdd.n2055 19.3944
R4143 vdd.n2109 vdd.n2108 19.3944
R4144 vdd.n2108 vdd.n2107 19.3944
R4145 vdd.n2107 vdd.n2062 19.3944
R4146 vdd.n2102 vdd.n2062 19.3944
R4147 vdd.n2102 vdd.n2101 19.3944
R4148 vdd.n2101 vdd.n2100 19.3944
R4149 vdd.n2100 vdd.n2069 19.3944
R4150 vdd.n2095 vdd.n2069 19.3944
R4151 vdd.n2095 vdd.n2094 19.3944
R4152 vdd.n2094 vdd.n2093 19.3944
R4153 vdd.n2093 vdd.n2077 19.3944
R4154 vdd.n2088 vdd.n2077 19.3944
R4155 vdd.n2088 vdd.n2087 19.3944
R4156 vdd.n2083 vdd.n2082 19.3944
R4157 vdd.n2203 vdd.n1148 19.3944
R4158 vdd.n2153 vdd.n2009 19.3944
R4159 vdd.n2153 vdd.n2015 19.3944
R4160 vdd.n2148 vdd.n2015 19.3944
R4161 vdd.n2148 vdd.n2147 19.3944
R4162 vdd.n2147 vdd.n2146 19.3944
R4163 vdd.n2146 vdd.n2022 19.3944
R4164 vdd.n2141 vdd.n2022 19.3944
R4165 vdd.n2141 vdd.n2140 19.3944
R4166 vdd.n2140 vdd.n2139 19.3944
R4167 vdd.n2139 vdd.n2029 19.3944
R4168 vdd.n2134 vdd.n2029 19.3944
R4169 vdd.n2134 vdd.n2133 19.3944
R4170 vdd.n2133 vdd.n2132 19.3944
R4171 vdd.n2132 vdd.n2036 19.3944
R4172 vdd.n2127 vdd.n2036 19.3944
R4173 vdd.n2127 vdd.n2126 19.3944
R4174 vdd.n2126 vdd.n2125 19.3944
R4175 vdd.n2125 vdd.n2043 19.3944
R4176 vdd.n2120 vdd.n2043 19.3944
R4177 vdd.n2120 vdd.n2119 19.3944
R4178 vdd.n2191 vdd.n2190 19.3944
R4179 vdd.n2190 vdd.n1981 19.3944
R4180 vdd.n2185 vdd.n2184 19.3944
R4181 vdd.n2180 vdd.n1985 19.3944
R4182 vdd.n2180 vdd.n1987 19.3944
R4183 vdd.n1990 vdd.n1987 19.3944
R4184 vdd.n2173 vdd.n1990 19.3944
R4185 vdd.n2173 vdd.n2172 19.3944
R4186 vdd.n2172 vdd.n2171 19.3944
R4187 vdd.n2171 vdd.n1996 19.3944
R4188 vdd.n2166 vdd.n1996 19.3944
R4189 vdd.n2166 vdd.n2165 19.3944
R4190 vdd.n2165 vdd.n2164 19.3944
R4191 vdd.n2164 vdd.n2003 19.3944
R4192 vdd.n2159 vdd.n2003 19.3944
R4193 vdd.n2159 vdd.n2158 19.3944
R4194 vdd.n1505 vdd.n1270 19.3944
R4195 vdd.n1505 vdd.n1261 19.3944
R4196 vdd.n1518 vdd.n1261 19.3944
R4197 vdd.n1518 vdd.n1259 19.3944
R4198 vdd.n1522 vdd.n1259 19.3944
R4199 vdd.n1522 vdd.n1250 19.3944
R4200 vdd.n1535 vdd.n1250 19.3944
R4201 vdd.n1535 vdd.n1248 19.3944
R4202 vdd.n1539 vdd.n1248 19.3944
R4203 vdd.n1539 vdd.n1239 19.3944
R4204 vdd.n1551 vdd.n1239 19.3944
R4205 vdd.n1551 vdd.n1237 19.3944
R4206 vdd.n1555 vdd.n1237 19.3944
R4207 vdd.n1555 vdd.n1227 19.3944
R4208 vdd.n1568 vdd.n1227 19.3944
R4209 vdd.n1568 vdd.n1225 19.3944
R4210 vdd.n1572 vdd.n1225 19.3944
R4211 vdd.n1572 vdd.n1216 19.3944
R4212 vdd.n1584 vdd.n1216 19.3944
R4213 vdd.n1584 vdd.n1214 19.3944
R4214 vdd.n1895 vdd.n1214 19.3944
R4215 vdd.n1895 vdd.n1204 19.3944
R4216 vdd.n1908 vdd.n1204 19.3944
R4217 vdd.n1908 vdd.n1202 19.3944
R4218 vdd.n1912 vdd.n1202 19.3944
R4219 vdd.n1912 vdd.n1193 19.3944
R4220 vdd.n1925 vdd.n1193 19.3944
R4221 vdd.n1925 vdd.n1191 19.3944
R4222 vdd.n1929 vdd.n1191 19.3944
R4223 vdd.n1929 vdd.n1182 19.3944
R4224 vdd.n1941 vdd.n1182 19.3944
R4225 vdd.n1941 vdd.n1180 19.3944
R4226 vdd.n1945 vdd.n1180 19.3944
R4227 vdd.n1945 vdd.n1170 19.3944
R4228 vdd.n1958 vdd.n1170 19.3944
R4229 vdd.n1958 vdd.n1168 19.3944
R4230 vdd.n1962 vdd.n1168 19.3944
R4231 vdd.n1962 vdd.n1158 19.3944
R4232 vdd.n1977 vdd.n1158 19.3944
R4233 vdd.n1977 vdd.n1156 19.3944
R4234 vdd.n2194 vdd.n1156 19.3944
R4235 vdd.n3411 vdd.n686 19.3944
R4236 vdd.n3411 vdd.n676 19.3944
R4237 vdd.n3423 vdd.n676 19.3944
R4238 vdd.n3423 vdd.n674 19.3944
R4239 vdd.n3427 vdd.n674 19.3944
R4240 vdd.n3427 vdd.n666 19.3944
R4241 vdd.n3440 vdd.n666 19.3944
R4242 vdd.n3440 vdd.n664 19.3944
R4243 vdd.n3444 vdd.n664 19.3944
R4244 vdd.n3444 vdd.n653 19.3944
R4245 vdd.n3456 vdd.n653 19.3944
R4246 vdd.n3456 vdd.n651 19.3944
R4247 vdd.n3460 vdd.n651 19.3944
R4248 vdd.n3460 vdd.n642 19.3944
R4249 vdd.n3473 vdd.n642 19.3944
R4250 vdd.n3473 vdd.n640 19.3944
R4251 vdd.n3480 vdd.n640 19.3944
R4252 vdd.n3480 vdd.n3479 19.3944
R4253 vdd.n3479 vdd.n631 19.3944
R4254 vdd.n3493 vdd.n631 19.3944
R4255 vdd.n3494 vdd.n3493 19.3944
R4256 vdd.n3494 vdd.n629 19.3944
R4257 vdd.n3498 vdd.n629 19.3944
R4258 vdd.n3500 vdd.n3498 19.3944
R4259 vdd.n3501 vdd.n3500 19.3944
R4260 vdd.n3501 vdd.n627 19.3944
R4261 vdd.n3505 vdd.n627 19.3944
R4262 vdd.n3507 vdd.n3505 19.3944
R4263 vdd.n3508 vdd.n3507 19.3944
R4264 vdd.n3508 vdd.n625 19.3944
R4265 vdd.n3512 vdd.n625 19.3944
R4266 vdd.n3515 vdd.n3512 19.3944
R4267 vdd.n3516 vdd.n3515 19.3944
R4268 vdd.n3516 vdd.n623 19.3944
R4269 vdd.n3520 vdd.n623 19.3944
R4270 vdd.n3522 vdd.n3520 19.3944
R4271 vdd.n3523 vdd.n3522 19.3944
R4272 vdd.n3523 vdd.n621 19.3944
R4273 vdd.n3527 vdd.n621 19.3944
R4274 vdd.n3529 vdd.n3527 19.3944
R4275 vdd.n3530 vdd.n3529 19.3944
R4276 vdd.n569 vdd.n438 19.3944
R4277 vdd.n575 vdd.n438 19.3944
R4278 vdd.n576 vdd.n575 19.3944
R4279 vdd.n579 vdd.n576 19.3944
R4280 vdd.n579 vdd.n436 19.3944
R4281 vdd.n585 vdd.n436 19.3944
R4282 vdd.n586 vdd.n585 19.3944
R4283 vdd.n589 vdd.n586 19.3944
R4284 vdd.n589 vdd.n434 19.3944
R4285 vdd.n595 vdd.n434 19.3944
R4286 vdd.n596 vdd.n595 19.3944
R4287 vdd.n599 vdd.n596 19.3944
R4288 vdd.n599 vdd.n432 19.3944
R4289 vdd.n605 vdd.n432 19.3944
R4290 vdd.n606 vdd.n605 19.3944
R4291 vdd.n609 vdd.n606 19.3944
R4292 vdd.n609 vdd.n430 19.3944
R4293 vdd.n615 vdd.n430 19.3944
R4294 vdd.n617 vdd.n615 19.3944
R4295 vdd.n618 vdd.n617 19.3944
R4296 vdd.n516 vdd.n515 19.3944
R4297 vdd.n519 vdd.n516 19.3944
R4298 vdd.n519 vdd.n450 19.3944
R4299 vdd.n525 vdd.n450 19.3944
R4300 vdd.n526 vdd.n525 19.3944
R4301 vdd.n529 vdd.n526 19.3944
R4302 vdd.n529 vdd.n448 19.3944
R4303 vdd.n535 vdd.n448 19.3944
R4304 vdd.n536 vdd.n535 19.3944
R4305 vdd.n539 vdd.n536 19.3944
R4306 vdd.n539 vdd.n446 19.3944
R4307 vdd.n545 vdd.n446 19.3944
R4308 vdd.n546 vdd.n545 19.3944
R4309 vdd.n549 vdd.n546 19.3944
R4310 vdd.n549 vdd.n444 19.3944
R4311 vdd.n555 vdd.n444 19.3944
R4312 vdd.n556 vdd.n555 19.3944
R4313 vdd.n559 vdd.n556 19.3944
R4314 vdd.n559 vdd.n442 19.3944
R4315 vdd.n565 vdd.n442 19.3944
R4316 vdd.n466 vdd.n465 19.3944
R4317 vdd.n469 vdd.n466 19.3944
R4318 vdd.n469 vdd.n462 19.3944
R4319 vdd.n475 vdd.n462 19.3944
R4320 vdd.n476 vdd.n475 19.3944
R4321 vdd.n479 vdd.n476 19.3944
R4322 vdd.n479 vdd.n460 19.3944
R4323 vdd.n485 vdd.n460 19.3944
R4324 vdd.n486 vdd.n485 19.3944
R4325 vdd.n489 vdd.n486 19.3944
R4326 vdd.n489 vdd.n458 19.3944
R4327 vdd.n495 vdd.n458 19.3944
R4328 vdd.n496 vdd.n495 19.3944
R4329 vdd.n499 vdd.n496 19.3944
R4330 vdd.n499 vdd.n456 19.3944
R4331 vdd.n505 vdd.n456 19.3944
R4332 vdd.n506 vdd.n505 19.3944
R4333 vdd.n509 vdd.n506 19.3944
R4334 vdd.n3415 vdd.n683 19.3944
R4335 vdd.n3415 vdd.n681 19.3944
R4336 vdd.n3419 vdd.n681 19.3944
R4337 vdd.n3419 vdd.n671 19.3944
R4338 vdd.n3432 vdd.n671 19.3944
R4339 vdd.n3432 vdd.n669 19.3944
R4340 vdd.n3436 vdd.n669 19.3944
R4341 vdd.n3436 vdd.n660 19.3944
R4342 vdd.n3448 vdd.n660 19.3944
R4343 vdd.n3448 vdd.n658 19.3944
R4344 vdd.n3452 vdd.n658 19.3944
R4345 vdd.n3452 vdd.n648 19.3944
R4346 vdd.n3465 vdd.n648 19.3944
R4347 vdd.n3465 vdd.n646 19.3944
R4348 vdd.n3469 vdd.n646 19.3944
R4349 vdd.n3469 vdd.n637 19.3944
R4350 vdd.n3484 vdd.n637 19.3944
R4351 vdd.n3484 vdd.n635 19.3944
R4352 vdd.n3488 vdd.n635 19.3944
R4353 vdd.n3488 vdd.n336 19.3944
R4354 vdd.n3579 vdd.n336 19.3944
R4355 vdd.n3579 vdd.n337 19.3944
R4356 vdd.n3573 vdd.n337 19.3944
R4357 vdd.n3573 vdd.n3572 19.3944
R4358 vdd.n3572 vdd.n3571 19.3944
R4359 vdd.n3571 vdd.n349 19.3944
R4360 vdd.n3565 vdd.n349 19.3944
R4361 vdd.n3565 vdd.n3564 19.3944
R4362 vdd.n3564 vdd.n3563 19.3944
R4363 vdd.n3563 vdd.n359 19.3944
R4364 vdd.n3557 vdd.n359 19.3944
R4365 vdd.n3557 vdd.n3556 19.3944
R4366 vdd.n3556 vdd.n3555 19.3944
R4367 vdd.n3555 vdd.n370 19.3944
R4368 vdd.n3549 vdd.n370 19.3944
R4369 vdd.n3549 vdd.n3548 19.3944
R4370 vdd.n3548 vdd.n3547 19.3944
R4371 vdd.n3547 vdd.n381 19.3944
R4372 vdd.n3541 vdd.n381 19.3944
R4373 vdd.n3541 vdd.n3540 19.3944
R4374 vdd.n3540 vdd.n3539 19.3944
R4375 vdd.n3362 vdd.n747 19.3944
R4376 vdd.n3362 vdd.n3359 19.3944
R4377 vdd.n3359 vdd.n3356 19.3944
R4378 vdd.n3356 vdd.n3355 19.3944
R4379 vdd.n3355 vdd.n3352 19.3944
R4380 vdd.n3352 vdd.n3351 19.3944
R4381 vdd.n3351 vdd.n3348 19.3944
R4382 vdd.n3348 vdd.n3347 19.3944
R4383 vdd.n3347 vdd.n3344 19.3944
R4384 vdd.n3344 vdd.n3343 19.3944
R4385 vdd.n3343 vdd.n3340 19.3944
R4386 vdd.n3340 vdd.n3339 19.3944
R4387 vdd.n3339 vdd.n3336 19.3944
R4388 vdd.n3336 vdd.n3335 19.3944
R4389 vdd.n3335 vdd.n3332 19.3944
R4390 vdd.n3332 vdd.n3331 19.3944
R4391 vdd.n3331 vdd.n3328 19.3944
R4392 vdd.n3328 vdd.n3327 19.3944
R4393 vdd.n3327 vdd.n3324 19.3944
R4394 vdd.n3324 vdd.n3323 19.3944
R4395 vdd.n3402 vdd.n3401 19.3944
R4396 vdd.n3401 vdd.n3400 19.3944
R4397 vdd.n732 vdd.n729 19.3944
R4398 vdd.n3396 vdd.n3395 19.3944
R4399 vdd.n3395 vdd.n3392 19.3944
R4400 vdd.n3392 vdd.n3391 19.3944
R4401 vdd.n3391 vdd.n3388 19.3944
R4402 vdd.n3388 vdd.n3387 19.3944
R4403 vdd.n3387 vdd.n3384 19.3944
R4404 vdd.n3384 vdd.n3383 19.3944
R4405 vdd.n3383 vdd.n3380 19.3944
R4406 vdd.n3380 vdd.n3379 19.3944
R4407 vdd.n3379 vdd.n3376 19.3944
R4408 vdd.n3376 vdd.n3375 19.3944
R4409 vdd.n3375 vdd.n3372 19.3944
R4410 vdd.n3372 vdd.n3371 19.3944
R4411 vdd.n3316 vdd.n767 19.3944
R4412 vdd.n3316 vdd.n3313 19.3944
R4413 vdd.n3313 vdd.n3310 19.3944
R4414 vdd.n3310 vdd.n3309 19.3944
R4415 vdd.n3309 vdd.n3306 19.3944
R4416 vdd.n3306 vdd.n3305 19.3944
R4417 vdd.n3305 vdd.n3302 19.3944
R4418 vdd.n3302 vdd.n3301 19.3944
R4419 vdd.n3301 vdd.n3298 19.3944
R4420 vdd.n3298 vdd.n3297 19.3944
R4421 vdd.n3297 vdd.n3294 19.3944
R4422 vdd.n3294 vdd.n3293 19.3944
R4423 vdd.n3293 vdd.n3290 19.3944
R4424 vdd.n3290 vdd.n3289 19.3944
R4425 vdd.n3289 vdd.n3286 19.3944
R4426 vdd.n3286 vdd.n3285 19.3944
R4427 vdd.n3282 vdd.n3281 19.3944
R4428 vdd.n3278 vdd.n3277 19.3944
R4429 vdd.n1437 vdd.n1433 19.0066
R4430 vdd.n2118 vdd.n2049 19.0066
R4431 vdd.n569 vdd.n566 19.0066
R4432 vdd.n3320 vdd.n767 19.0066
R4433 vdd.n1137 vdd.n1136 16.0975
R4434 vdd.n998 vdd.n997 16.0975
R4435 vdd.n1398 vdd.n1397 16.0975
R4436 vdd.n1436 vdd.n1435 16.0975
R4437 vdd.n1332 vdd.n1331 16.0975
R4438 vdd.n2201 vdd.n2200 16.0975
R4439 vdd.n2051 vdd.n2050 16.0975
R4440 vdd.n2011 vdd.n2010 16.0975
R4441 vdd.n1131 vdd.n1130 16.0975
R4442 vdd.n989 vdd.n988 16.0975
R4443 vdd.n2762 vdd.n2761 16.0975
R4444 vdd.n427 vdd.n426 16.0975
R4445 vdd.n441 vdd.n440 16.0975
R4446 vdd.n453 vdd.n452 16.0975
R4447 vdd.n769 vdd.n768 16.0975
R4448 vdd.n3367 vdd.n3366 16.0975
R4449 vdd.n833 vdd.n832 16.0975
R4450 vdd.n2831 vdd.n2830 16.0975
R4451 vdd.n689 vdd.n688 16.0975
R4452 vdd.n800 vdd.n799 16.0975
R4453 vdd.t128 vdd.n2726 15.4182
R4454 vdd.n3010 vdd.t125 15.4182
R4455 vdd.n28 vdd.n27 14.8356
R4456 vdd.n2467 vdd.n1110 13.6043
R4457 vdd.n3241 vdd.n692 13.6043
R4458 vdd.n328 vdd.n293 13.1884
R4459 vdd.n269 vdd.n234 13.1884
R4460 vdd.n226 vdd.n191 13.1884
R4461 vdd.n167 vdd.n132 13.1884
R4462 vdd.n125 vdd.n90 13.1884
R4463 vdd.n66 vdd.n31 13.1884
R4464 vdd.n1827 vdd.n1792 13.1884
R4465 vdd.n1886 vdd.n1851 13.1884
R4466 vdd.n1725 vdd.n1690 13.1884
R4467 vdd.n1784 vdd.n1749 13.1884
R4468 vdd.n1624 vdd.n1589 13.1884
R4469 vdd.n1683 vdd.n1648 13.1884
R4470 vdd.n1468 vdd.n1333 12.9944
R4471 vdd.n1472 vdd.n1333 12.9944
R4472 vdd.n2157 vdd.n2009 12.9944
R4473 vdd.n2158 vdd.n2157 12.9944
R4474 vdd.n515 vdd.n454 12.9944
R4475 vdd.n509 vdd.n454 12.9944
R4476 vdd.n3368 vdd.n747 12.9944
R4477 vdd.n3371 vdd.n3368 12.9944
R4478 vdd.n329 vdd.n291 12.8005
R4479 vdd.n324 vdd.n295 12.8005
R4480 vdd.n270 vdd.n232 12.8005
R4481 vdd.n265 vdd.n236 12.8005
R4482 vdd.n227 vdd.n189 12.8005
R4483 vdd.n222 vdd.n193 12.8005
R4484 vdd.n168 vdd.n130 12.8005
R4485 vdd.n163 vdd.n134 12.8005
R4486 vdd.n126 vdd.n88 12.8005
R4487 vdd.n121 vdd.n92 12.8005
R4488 vdd.n67 vdd.n29 12.8005
R4489 vdd.n62 vdd.n33 12.8005
R4490 vdd.n1828 vdd.n1790 12.8005
R4491 vdd.n1823 vdd.n1794 12.8005
R4492 vdd.n1887 vdd.n1849 12.8005
R4493 vdd.n1882 vdd.n1853 12.8005
R4494 vdd.n1726 vdd.n1688 12.8005
R4495 vdd.n1721 vdd.n1692 12.8005
R4496 vdd.n1785 vdd.n1747 12.8005
R4497 vdd.n1780 vdd.n1751 12.8005
R4498 vdd.n1625 vdd.n1587 12.8005
R4499 vdd.n1620 vdd.n1591 12.8005
R4500 vdd.n1684 vdd.n1646 12.8005
R4501 vdd.n1679 vdd.n1650 12.8005
R4502 vdd.n323 vdd.n296 12.0247
R4503 vdd.n264 vdd.n237 12.0247
R4504 vdd.n221 vdd.n194 12.0247
R4505 vdd.n162 vdd.n135 12.0247
R4506 vdd.n120 vdd.n93 12.0247
R4507 vdd.n61 vdd.n34 12.0247
R4508 vdd.n1822 vdd.n1795 12.0247
R4509 vdd.n1881 vdd.n1854 12.0247
R4510 vdd.n1720 vdd.n1693 12.0247
R4511 vdd.n1779 vdd.n1752 12.0247
R4512 vdd.n1619 vdd.n1592 12.0247
R4513 vdd.n1678 vdd.n1651 12.0247
R4514 vdd.n1507 vdd.n1263 11.337
R4515 vdd.n1516 vdd.n1263 11.337
R4516 vdd.n1516 vdd.n1515 11.337
R4517 vdd.n1524 vdd.n1257 11.337
R4518 vdd.n1533 vdd.n1532 11.337
R4519 vdd.n1549 vdd.n1241 11.337
R4520 vdd.n1557 vdd.n1234 11.337
R4521 vdd.n1566 vdd.n1565 11.337
R4522 vdd.n1574 vdd.n1223 11.337
R4523 vdd.n1897 vdd.n1212 11.337
R4524 vdd.n1906 vdd.n1206 11.337
R4525 vdd.n1914 vdd.n1200 11.337
R4526 vdd.n1923 vdd.n1922 11.337
R4527 vdd.n1939 vdd.n1184 11.337
R4528 vdd.n1947 vdd.n1177 11.337
R4529 vdd.n1956 vdd.n1955 11.337
R4530 vdd.n1964 vdd.n1160 11.337
R4531 vdd.n1975 vdd.n1160 11.337
R4532 vdd.n1975 vdd.n1974 11.337
R4533 vdd.n3413 vdd.n678 11.337
R4534 vdd.n3421 vdd.n678 11.337
R4535 vdd.n3421 vdd.n679 11.337
R4536 vdd.n3430 vdd.n3429 11.337
R4537 vdd.n3446 vdd.n662 11.337
R4538 vdd.n3454 vdd.n655 11.337
R4539 vdd.n3463 vdd.n3462 11.337
R4540 vdd.n3471 vdd.n644 11.337
R4541 vdd.n3490 vdd.n633 11.337
R4542 vdd.n3577 vdd.n340 11.337
R4543 vdd.n3575 vdd.n344 11.337
R4544 vdd.n3569 vdd.n3568 11.337
R4545 vdd.n3561 vdd.n361 11.337
R4546 vdd.n3560 vdd.n3559 11.337
R4547 vdd.n3553 vdd.n3552 11.337
R4548 vdd.n3551 vdd.n375 11.337
R4549 vdd.n3545 vdd.n3544 11.337
R4550 vdd.n3544 vdd.n3543 11.337
R4551 vdd.n3543 vdd.n386 11.337
R4552 vdd.n320 vdd.n319 11.249
R4553 vdd.n261 vdd.n260 11.249
R4554 vdd.n218 vdd.n217 11.249
R4555 vdd.n159 vdd.n158 11.249
R4556 vdd.n117 vdd.n116 11.249
R4557 vdd.n58 vdd.n57 11.249
R4558 vdd.n1819 vdd.n1818 11.249
R4559 vdd.n1878 vdd.n1877 11.249
R4560 vdd.n1717 vdd.n1716 11.249
R4561 vdd.n1776 vdd.n1775 11.249
R4562 vdd.n1616 vdd.n1615 11.249
R4563 vdd.n1675 vdd.n1674 11.249
R4564 vdd.n1305 vdd.t64 11.2237
R4565 vdd.n3537 vdd.t34 11.2237
R4566 vdd.t204 vdd.n1178 10.7702
R4567 vdd.n3438 vdd.t187 10.7702
R4568 vdd.n305 vdd.n304 10.7238
R4569 vdd.n246 vdd.n245 10.7238
R4570 vdd.n203 vdd.n202 10.7238
R4571 vdd.n144 vdd.n143 10.7238
R4572 vdd.n102 vdd.n101 10.7238
R4573 vdd.n43 vdd.n42 10.7238
R4574 vdd.n1804 vdd.n1803 10.7238
R4575 vdd.n1863 vdd.n1862 10.7238
R4576 vdd.n1702 vdd.n1701 10.7238
R4577 vdd.n1761 vdd.n1760 10.7238
R4578 vdd.n1601 vdd.n1600 10.7238
R4579 vdd.n1660 vdd.n1659 10.7238
R4580 vdd.n2465 vdd.n1102 10.6151
R4581 vdd.n2475 vdd.n1102 10.6151
R4582 vdd.n2476 vdd.n2475 10.6151
R4583 vdd.n2477 vdd.n2476 10.6151
R4584 vdd.n2477 vdd.n1090 10.6151
R4585 vdd.n2487 vdd.n1090 10.6151
R4586 vdd.n2488 vdd.n2487 10.6151
R4587 vdd.n2489 vdd.n2488 10.6151
R4588 vdd.n2489 vdd.n1078 10.6151
R4589 vdd.n2499 vdd.n1078 10.6151
R4590 vdd.n2500 vdd.n2499 10.6151
R4591 vdd.n2501 vdd.n2500 10.6151
R4592 vdd.n2501 vdd.n1065 10.6151
R4593 vdd.n2511 vdd.n1065 10.6151
R4594 vdd.n2512 vdd.n2511 10.6151
R4595 vdd.n2513 vdd.n2512 10.6151
R4596 vdd.n2513 vdd.n1053 10.6151
R4597 vdd.n2524 vdd.n1053 10.6151
R4598 vdd.n2525 vdd.n2524 10.6151
R4599 vdd.n2526 vdd.n2525 10.6151
R4600 vdd.n2526 vdd.n1041 10.6151
R4601 vdd.n2536 vdd.n1041 10.6151
R4602 vdd.n2537 vdd.n2536 10.6151
R4603 vdd.n2538 vdd.n2537 10.6151
R4604 vdd.n2538 vdd.n1029 10.6151
R4605 vdd.n2548 vdd.n1029 10.6151
R4606 vdd.n2549 vdd.n2548 10.6151
R4607 vdd.n2550 vdd.n2549 10.6151
R4608 vdd.n2550 vdd.n1019 10.6151
R4609 vdd.n2560 vdd.n1019 10.6151
R4610 vdd.n2561 vdd.n2560 10.6151
R4611 vdd.n2562 vdd.n2561 10.6151
R4612 vdd.n2562 vdd.n1006 10.6151
R4613 vdd.n2574 vdd.n1006 10.6151
R4614 vdd.n2575 vdd.n2574 10.6151
R4615 vdd.n2577 vdd.n2575 10.6151
R4616 vdd.n2577 vdd.n2576 10.6151
R4617 vdd.n2576 vdd.n987 10.6151
R4618 vdd.n2724 vdd.n2723 10.6151
R4619 vdd.n2723 vdd.n2722 10.6151
R4620 vdd.n2722 vdd.n2719 10.6151
R4621 vdd.n2719 vdd.n2718 10.6151
R4622 vdd.n2718 vdd.n2715 10.6151
R4623 vdd.n2715 vdd.n2714 10.6151
R4624 vdd.n2714 vdd.n2711 10.6151
R4625 vdd.n2711 vdd.n2710 10.6151
R4626 vdd.n2710 vdd.n2707 10.6151
R4627 vdd.n2707 vdd.n2706 10.6151
R4628 vdd.n2706 vdd.n2703 10.6151
R4629 vdd.n2703 vdd.n2702 10.6151
R4630 vdd.n2702 vdd.n2699 10.6151
R4631 vdd.n2699 vdd.n2698 10.6151
R4632 vdd.n2698 vdd.n2695 10.6151
R4633 vdd.n2695 vdd.n2694 10.6151
R4634 vdd.n2694 vdd.n2691 10.6151
R4635 vdd.n2691 vdd.n2690 10.6151
R4636 vdd.n2690 vdd.n2687 10.6151
R4637 vdd.n2687 vdd.n2686 10.6151
R4638 vdd.n2686 vdd.n2683 10.6151
R4639 vdd.n2683 vdd.n2682 10.6151
R4640 vdd.n2682 vdd.n2679 10.6151
R4641 vdd.n2679 vdd.n2678 10.6151
R4642 vdd.n2678 vdd.n2675 10.6151
R4643 vdd.n2675 vdd.n2674 10.6151
R4644 vdd.n2674 vdd.n2671 10.6151
R4645 vdd.n2671 vdd.n2670 10.6151
R4646 vdd.n2670 vdd.n2667 10.6151
R4647 vdd.n2667 vdd.n2666 10.6151
R4648 vdd.n2666 vdd.n2663 10.6151
R4649 vdd.n2661 vdd.n2658 10.6151
R4650 vdd.n2658 vdd.n2657 10.6151
R4651 vdd.n2394 vdd.n2393 10.6151
R4652 vdd.n2393 vdd.n2391 10.6151
R4653 vdd.n2391 vdd.n2390 10.6151
R4654 vdd.n2390 vdd.n2388 10.6151
R4655 vdd.n2388 vdd.n2387 10.6151
R4656 vdd.n2387 vdd.n2385 10.6151
R4657 vdd.n2385 vdd.n2384 10.6151
R4658 vdd.n2384 vdd.n2382 10.6151
R4659 vdd.n2382 vdd.n2381 10.6151
R4660 vdd.n2381 vdd.n2379 10.6151
R4661 vdd.n2379 vdd.n2378 10.6151
R4662 vdd.n2378 vdd.n2376 10.6151
R4663 vdd.n2376 vdd.n2375 10.6151
R4664 vdd.n2375 vdd.n2373 10.6151
R4665 vdd.n2373 vdd.n2372 10.6151
R4666 vdd.n2372 vdd.n2370 10.6151
R4667 vdd.n2370 vdd.n2369 10.6151
R4668 vdd.n2369 vdd.n2367 10.6151
R4669 vdd.n2367 vdd.n2366 10.6151
R4670 vdd.n2366 vdd.n2364 10.6151
R4671 vdd.n2364 vdd.n2363 10.6151
R4672 vdd.n2363 vdd.n2361 10.6151
R4673 vdd.n2361 vdd.n2360 10.6151
R4674 vdd.n2360 vdd.n1133 10.6151
R4675 vdd.n2327 vdd.n1133 10.6151
R4676 vdd.n2328 vdd.n2327 10.6151
R4677 vdd.n2330 vdd.n2328 10.6151
R4678 vdd.n2331 vdd.n2330 10.6151
R4679 vdd.n2344 vdd.n2331 10.6151
R4680 vdd.n2344 vdd.n2343 10.6151
R4681 vdd.n2343 vdd.n2342 10.6151
R4682 vdd.n2342 vdd.n2340 10.6151
R4683 vdd.n2340 vdd.n2339 10.6151
R4684 vdd.n2339 vdd.n2337 10.6151
R4685 vdd.n2337 vdd.n2336 10.6151
R4686 vdd.n2336 vdd.n2333 10.6151
R4687 vdd.n2333 vdd.n2332 10.6151
R4688 vdd.n2332 vdd.n990 10.6151
R4689 vdd.n2464 vdd.n2463 10.6151
R4690 vdd.n2463 vdd.n1114 10.6151
R4691 vdd.n2458 vdd.n1114 10.6151
R4692 vdd.n2458 vdd.n2457 10.6151
R4693 vdd.n2457 vdd.n1116 10.6151
R4694 vdd.n2452 vdd.n1116 10.6151
R4695 vdd.n2452 vdd.n2451 10.6151
R4696 vdd.n2451 vdd.n2450 10.6151
R4697 vdd.n2450 vdd.n1118 10.6151
R4698 vdd.n2444 vdd.n1118 10.6151
R4699 vdd.n2444 vdd.n2443 10.6151
R4700 vdd.n2443 vdd.n2442 10.6151
R4701 vdd.n2442 vdd.n1120 10.6151
R4702 vdd.n2436 vdd.n1120 10.6151
R4703 vdd.n2436 vdd.n2435 10.6151
R4704 vdd.n2435 vdd.n2434 10.6151
R4705 vdd.n2434 vdd.n1122 10.6151
R4706 vdd.n2428 vdd.n1122 10.6151
R4707 vdd.n2428 vdd.n2427 10.6151
R4708 vdd.n2427 vdd.n2426 10.6151
R4709 vdd.n2426 vdd.n1124 10.6151
R4710 vdd.n2420 vdd.n1124 10.6151
R4711 vdd.n2420 vdd.n2419 10.6151
R4712 vdd.n2419 vdd.n2418 10.6151
R4713 vdd.n2418 vdd.n1126 10.6151
R4714 vdd.n2412 vdd.n1126 10.6151
R4715 vdd.n2412 vdd.n2411 10.6151
R4716 vdd.n2411 vdd.n2410 10.6151
R4717 vdd.n2410 vdd.n1128 10.6151
R4718 vdd.n2404 vdd.n1128 10.6151
R4719 vdd.n2404 vdd.n2403 10.6151
R4720 vdd.n2401 vdd.n1132 10.6151
R4721 vdd.n2395 vdd.n1132 10.6151
R4722 vdd.n2899 vdd.n2897 10.6151
R4723 vdd.n2900 vdd.n2899 10.6151
R4724 vdd.n2999 vdd.n2900 10.6151
R4725 vdd.n2999 vdd.n2998 10.6151
R4726 vdd.n2998 vdd.n2997 10.6151
R4727 vdd.n2997 vdd.n2995 10.6151
R4728 vdd.n2995 vdd.n2994 10.6151
R4729 vdd.n2994 vdd.n2992 10.6151
R4730 vdd.n2992 vdd.n2991 10.6151
R4731 vdd.n2991 vdd.n2901 10.6151
R4732 vdd.n2941 vdd.n2901 10.6151
R4733 vdd.n2942 vdd.n2941 10.6151
R4734 vdd.n2944 vdd.n2942 10.6151
R4735 vdd.n2945 vdd.n2944 10.6151
R4736 vdd.n2975 vdd.n2945 10.6151
R4737 vdd.n2975 vdd.n2974 10.6151
R4738 vdd.n2974 vdd.n2973 10.6151
R4739 vdd.n2973 vdd.n2971 10.6151
R4740 vdd.n2971 vdd.n2970 10.6151
R4741 vdd.n2970 vdd.n2968 10.6151
R4742 vdd.n2968 vdd.n2967 10.6151
R4743 vdd.n2967 vdd.n2965 10.6151
R4744 vdd.n2965 vdd.n2964 10.6151
R4745 vdd.n2964 vdd.n2962 10.6151
R4746 vdd.n2962 vdd.n2961 10.6151
R4747 vdd.n2961 vdd.n2959 10.6151
R4748 vdd.n2959 vdd.n2958 10.6151
R4749 vdd.n2958 vdd.n2956 10.6151
R4750 vdd.n2956 vdd.n2955 10.6151
R4751 vdd.n2955 vdd.n2953 10.6151
R4752 vdd.n2953 vdd.n2952 10.6151
R4753 vdd.n2952 vdd.n2950 10.6151
R4754 vdd.n2950 vdd.n2949 10.6151
R4755 vdd.n2949 vdd.n2947 10.6151
R4756 vdd.n2947 vdd.n2946 10.6151
R4757 vdd.n2946 vdd.n836 10.6151
R4758 vdd.n3174 vdd.n836 10.6151
R4759 vdd.n3175 vdd.n3174 10.6151
R4760 vdd.n3014 vdd.n3013 10.6151
R4761 vdd.n3013 vdd.n948 10.6151
R4762 vdd.n2833 vdd.n948 10.6151
R4763 vdd.n2834 vdd.n2833 10.6151
R4764 vdd.n2837 vdd.n2834 10.6151
R4765 vdd.n2838 vdd.n2837 10.6151
R4766 vdd.n2841 vdd.n2838 10.6151
R4767 vdd.n2842 vdd.n2841 10.6151
R4768 vdd.n2845 vdd.n2842 10.6151
R4769 vdd.n2846 vdd.n2845 10.6151
R4770 vdd.n2849 vdd.n2846 10.6151
R4771 vdd.n2850 vdd.n2849 10.6151
R4772 vdd.n2853 vdd.n2850 10.6151
R4773 vdd.n2854 vdd.n2853 10.6151
R4774 vdd.n2857 vdd.n2854 10.6151
R4775 vdd.n2858 vdd.n2857 10.6151
R4776 vdd.n2861 vdd.n2858 10.6151
R4777 vdd.n2862 vdd.n2861 10.6151
R4778 vdd.n2865 vdd.n2862 10.6151
R4779 vdd.n2866 vdd.n2865 10.6151
R4780 vdd.n2869 vdd.n2866 10.6151
R4781 vdd.n2870 vdd.n2869 10.6151
R4782 vdd.n2873 vdd.n2870 10.6151
R4783 vdd.n2874 vdd.n2873 10.6151
R4784 vdd.n2877 vdd.n2874 10.6151
R4785 vdd.n2878 vdd.n2877 10.6151
R4786 vdd.n2881 vdd.n2878 10.6151
R4787 vdd.n2882 vdd.n2881 10.6151
R4788 vdd.n2885 vdd.n2882 10.6151
R4789 vdd.n2886 vdd.n2885 10.6151
R4790 vdd.n2889 vdd.n2886 10.6151
R4791 vdd.n2894 vdd.n2891 10.6151
R4792 vdd.n2896 vdd.n2894 10.6151
R4793 vdd.n3015 vdd.n937 10.6151
R4794 vdd.n3025 vdd.n937 10.6151
R4795 vdd.n3026 vdd.n3025 10.6151
R4796 vdd.n3027 vdd.n3026 10.6151
R4797 vdd.n3027 vdd.n925 10.6151
R4798 vdd.n3037 vdd.n925 10.6151
R4799 vdd.n3038 vdd.n3037 10.6151
R4800 vdd.n3039 vdd.n3038 10.6151
R4801 vdd.n3039 vdd.n915 10.6151
R4802 vdd.n3049 vdd.n915 10.6151
R4803 vdd.n3050 vdd.n3049 10.6151
R4804 vdd.n3051 vdd.n3050 10.6151
R4805 vdd.n3051 vdd.n903 10.6151
R4806 vdd.n3061 vdd.n903 10.6151
R4807 vdd.n3062 vdd.n3061 10.6151
R4808 vdd.n3063 vdd.n3062 10.6151
R4809 vdd.n3063 vdd.n892 10.6151
R4810 vdd.n3073 vdd.n892 10.6151
R4811 vdd.n3074 vdd.n3073 10.6151
R4812 vdd.n3075 vdd.n3074 10.6151
R4813 vdd.n3075 vdd.n879 10.6151
R4814 vdd.n3086 vdd.n879 10.6151
R4815 vdd.n3087 vdd.n3086 10.6151
R4816 vdd.n3088 vdd.n3087 10.6151
R4817 vdd.n3088 vdd.n866 10.6151
R4818 vdd.n3098 vdd.n866 10.6151
R4819 vdd.n3099 vdd.n3098 10.6151
R4820 vdd.n3100 vdd.n3099 10.6151
R4821 vdd.n3100 vdd.n855 10.6151
R4822 vdd.n3110 vdd.n855 10.6151
R4823 vdd.n3111 vdd.n3110 10.6151
R4824 vdd.n3112 vdd.n3111 10.6151
R4825 vdd.n3112 vdd.n841 10.6151
R4826 vdd.n3167 vdd.n841 10.6151
R4827 vdd.n3168 vdd.n3167 10.6151
R4828 vdd.n3169 vdd.n3168 10.6151
R4829 vdd.n3169 vdd.n810 10.6151
R4830 vdd.n3239 vdd.n810 10.6151
R4831 vdd.n3238 vdd.n3237 10.6151
R4832 vdd.n3237 vdd.n811 10.6151
R4833 vdd.n812 vdd.n811 10.6151
R4834 vdd.n3230 vdd.n812 10.6151
R4835 vdd.n3230 vdd.n3229 10.6151
R4836 vdd.n3229 vdd.n3228 10.6151
R4837 vdd.n3228 vdd.n814 10.6151
R4838 vdd.n3223 vdd.n814 10.6151
R4839 vdd.n3223 vdd.n3222 10.6151
R4840 vdd.n3222 vdd.n3221 10.6151
R4841 vdd.n3221 vdd.n817 10.6151
R4842 vdd.n3216 vdd.n817 10.6151
R4843 vdd.n3216 vdd.n3215 10.6151
R4844 vdd.n3215 vdd.n3214 10.6151
R4845 vdd.n3214 vdd.n820 10.6151
R4846 vdd.n3209 vdd.n820 10.6151
R4847 vdd.n3209 vdd.n731 10.6151
R4848 vdd.n3205 vdd.n731 10.6151
R4849 vdd.n3205 vdd.n3204 10.6151
R4850 vdd.n3204 vdd.n3203 10.6151
R4851 vdd.n3203 vdd.n823 10.6151
R4852 vdd.n3198 vdd.n823 10.6151
R4853 vdd.n3198 vdd.n3197 10.6151
R4854 vdd.n3197 vdd.n3196 10.6151
R4855 vdd.n3196 vdd.n826 10.6151
R4856 vdd.n3191 vdd.n826 10.6151
R4857 vdd.n3191 vdd.n3190 10.6151
R4858 vdd.n3190 vdd.n3189 10.6151
R4859 vdd.n3189 vdd.n829 10.6151
R4860 vdd.n3184 vdd.n829 10.6151
R4861 vdd.n3184 vdd.n3183 10.6151
R4862 vdd.n3181 vdd.n834 10.6151
R4863 vdd.n3176 vdd.n834 10.6151
R4864 vdd.n3157 vdd.n3118 10.6151
R4865 vdd.n3152 vdd.n3118 10.6151
R4866 vdd.n3152 vdd.n3151 10.6151
R4867 vdd.n3151 vdd.n3150 10.6151
R4868 vdd.n3150 vdd.n3120 10.6151
R4869 vdd.n3145 vdd.n3120 10.6151
R4870 vdd.n3145 vdd.n3144 10.6151
R4871 vdd.n3144 vdd.n3143 10.6151
R4872 vdd.n3143 vdd.n3123 10.6151
R4873 vdd.n3138 vdd.n3123 10.6151
R4874 vdd.n3138 vdd.n3137 10.6151
R4875 vdd.n3137 vdd.n3136 10.6151
R4876 vdd.n3136 vdd.n3126 10.6151
R4877 vdd.n3131 vdd.n3126 10.6151
R4878 vdd.n3131 vdd.n3130 10.6151
R4879 vdd.n3130 vdd.n785 10.6151
R4880 vdd.n3274 vdd.n785 10.6151
R4881 vdd.n3274 vdd.n786 10.6151
R4882 vdd.n788 vdd.n786 10.6151
R4883 vdd.n3267 vdd.n788 10.6151
R4884 vdd.n3267 vdd.n3266 10.6151
R4885 vdd.n3266 vdd.n3265 10.6151
R4886 vdd.n3265 vdd.n790 10.6151
R4887 vdd.n3260 vdd.n790 10.6151
R4888 vdd.n3260 vdd.n3259 10.6151
R4889 vdd.n3259 vdd.n3258 10.6151
R4890 vdd.n3258 vdd.n793 10.6151
R4891 vdd.n3253 vdd.n793 10.6151
R4892 vdd.n3253 vdd.n3252 10.6151
R4893 vdd.n3252 vdd.n3251 10.6151
R4894 vdd.n3251 vdd.n796 10.6151
R4895 vdd.n3246 vdd.n3245 10.6151
R4896 vdd.n3245 vdd.n3244 10.6151
R4897 vdd.n3007 vdd.n3006 10.6151
R4898 vdd.n3006 vdd.n3004 10.6151
R4899 vdd.n3004 vdd.n3003 10.6151
R4900 vdd.n3003 vdd.n2829 10.6151
R4901 vdd.n2903 vdd.n2829 10.6151
R4902 vdd.n2904 vdd.n2903 10.6151
R4903 vdd.n2906 vdd.n2904 10.6151
R4904 vdd.n2907 vdd.n2906 10.6151
R4905 vdd.n2987 vdd.n2907 10.6151
R4906 vdd.n2987 vdd.n2986 10.6151
R4907 vdd.n2986 vdd.n2985 10.6151
R4908 vdd.n2985 vdd.n2983 10.6151
R4909 vdd.n2983 vdd.n2982 10.6151
R4910 vdd.n2982 vdd.n2980 10.6151
R4911 vdd.n2980 vdd.n2979 10.6151
R4912 vdd.n2979 vdd.n2939 10.6151
R4913 vdd.n2939 vdd.n2938 10.6151
R4914 vdd.n2938 vdd.n2936 10.6151
R4915 vdd.n2936 vdd.n2935 10.6151
R4916 vdd.n2935 vdd.n2933 10.6151
R4917 vdd.n2933 vdd.n2932 10.6151
R4918 vdd.n2932 vdd.n2930 10.6151
R4919 vdd.n2930 vdd.n2929 10.6151
R4920 vdd.n2929 vdd.n2927 10.6151
R4921 vdd.n2927 vdd.n2926 10.6151
R4922 vdd.n2926 vdd.n2924 10.6151
R4923 vdd.n2924 vdd.n2923 10.6151
R4924 vdd.n2923 vdd.n2921 10.6151
R4925 vdd.n2921 vdd.n2920 10.6151
R4926 vdd.n2920 vdd.n2918 10.6151
R4927 vdd.n2918 vdd.n2917 10.6151
R4928 vdd.n2917 vdd.n2915 10.6151
R4929 vdd.n2915 vdd.n2914 10.6151
R4930 vdd.n2914 vdd.n2912 10.6151
R4931 vdd.n2912 vdd.n2911 10.6151
R4932 vdd.n2911 vdd.n2909 10.6151
R4933 vdd.n2909 vdd.n2908 10.6151
R4934 vdd.n2908 vdd.n802 10.6151
R4935 vdd.n2764 vdd.n942 10.6151
R4936 vdd.n2767 vdd.n2764 10.6151
R4937 vdd.n2768 vdd.n2767 10.6151
R4938 vdd.n2771 vdd.n2768 10.6151
R4939 vdd.n2772 vdd.n2771 10.6151
R4940 vdd.n2775 vdd.n2772 10.6151
R4941 vdd.n2776 vdd.n2775 10.6151
R4942 vdd.n2779 vdd.n2776 10.6151
R4943 vdd.n2780 vdd.n2779 10.6151
R4944 vdd.n2783 vdd.n2780 10.6151
R4945 vdd.n2784 vdd.n2783 10.6151
R4946 vdd.n2787 vdd.n2784 10.6151
R4947 vdd.n2788 vdd.n2787 10.6151
R4948 vdd.n2791 vdd.n2788 10.6151
R4949 vdd.n2792 vdd.n2791 10.6151
R4950 vdd.n2795 vdd.n2792 10.6151
R4951 vdd.n2796 vdd.n2795 10.6151
R4952 vdd.n2799 vdd.n2796 10.6151
R4953 vdd.n2800 vdd.n2799 10.6151
R4954 vdd.n2803 vdd.n2800 10.6151
R4955 vdd.n2804 vdd.n2803 10.6151
R4956 vdd.n2807 vdd.n2804 10.6151
R4957 vdd.n2808 vdd.n2807 10.6151
R4958 vdd.n2811 vdd.n2808 10.6151
R4959 vdd.n2812 vdd.n2811 10.6151
R4960 vdd.n2815 vdd.n2812 10.6151
R4961 vdd.n2816 vdd.n2815 10.6151
R4962 vdd.n2819 vdd.n2816 10.6151
R4963 vdd.n2820 vdd.n2819 10.6151
R4964 vdd.n2823 vdd.n2820 10.6151
R4965 vdd.n2824 vdd.n2823 10.6151
R4966 vdd.n2828 vdd.n2827 10.6151
R4967 vdd.n3008 vdd.n2828 10.6151
R4968 vdd.n3020 vdd.n3019 10.6151
R4969 vdd.n3021 vdd.n3020 10.6151
R4970 vdd.n3021 vdd.n932 10.6151
R4971 vdd.n3031 vdd.n932 10.6151
R4972 vdd.n3032 vdd.n3031 10.6151
R4973 vdd.n3033 vdd.n3032 10.6151
R4974 vdd.n3033 vdd.n920 10.6151
R4975 vdd.n3043 vdd.n920 10.6151
R4976 vdd.n3044 vdd.n3043 10.6151
R4977 vdd.n3045 vdd.n3044 10.6151
R4978 vdd.n3045 vdd.n909 10.6151
R4979 vdd.n3055 vdd.n909 10.6151
R4980 vdd.n3056 vdd.n3055 10.6151
R4981 vdd.n3057 vdd.n3056 10.6151
R4982 vdd.n3057 vdd.n897 10.6151
R4983 vdd.n3067 vdd.n897 10.6151
R4984 vdd.n3068 vdd.n3067 10.6151
R4985 vdd.n3069 vdd.n3068 10.6151
R4986 vdd.n3069 vdd.n886 10.6151
R4987 vdd.n3079 vdd.n886 10.6151
R4988 vdd.n3082 vdd.n3081 10.6151
R4989 vdd.n3082 vdd.n872 10.6151
R4990 vdd.n3092 vdd.n872 10.6151
R4991 vdd.n3093 vdd.n3092 10.6151
R4992 vdd.n3094 vdd.n3093 10.6151
R4993 vdd.n3094 vdd.n860 10.6151
R4994 vdd.n3104 vdd.n860 10.6151
R4995 vdd.n3105 vdd.n3104 10.6151
R4996 vdd.n3106 vdd.n3105 10.6151
R4997 vdd.n3106 vdd.n849 10.6151
R4998 vdd.n3116 vdd.n849 10.6151
R4999 vdd.n3117 vdd.n3116 10.6151
R5000 vdd.n3163 vdd.n3117 10.6151
R5001 vdd.n3163 vdd.n3162 10.6151
R5002 vdd.n3162 vdd.n3161 10.6151
R5003 vdd.n3161 vdd.n3160 10.6151
R5004 vdd.n3160 vdd.n3158 10.6151
R5005 vdd.n2470 vdd.n2469 10.6151
R5006 vdd.n2471 vdd.n2470 10.6151
R5007 vdd.n2471 vdd.n1096 10.6151
R5008 vdd.n2481 vdd.n1096 10.6151
R5009 vdd.n2482 vdd.n2481 10.6151
R5010 vdd.n2483 vdd.n2482 10.6151
R5011 vdd.n2483 vdd.n1084 10.6151
R5012 vdd.n2493 vdd.n1084 10.6151
R5013 vdd.n2494 vdd.n2493 10.6151
R5014 vdd.n2495 vdd.n2494 10.6151
R5015 vdd.n2495 vdd.n1072 10.6151
R5016 vdd.n2505 vdd.n1072 10.6151
R5017 vdd.n2506 vdd.n2505 10.6151
R5018 vdd.n2507 vdd.n2506 10.6151
R5019 vdd.n2507 vdd.n1059 10.6151
R5020 vdd.n2517 vdd.n1059 10.6151
R5021 vdd.n2518 vdd.n2517 10.6151
R5022 vdd.n2520 vdd.n1047 10.6151
R5023 vdd.n2530 vdd.n1047 10.6151
R5024 vdd.n2531 vdd.n2530 10.6151
R5025 vdd.n2532 vdd.n2531 10.6151
R5026 vdd.n2532 vdd.n1035 10.6151
R5027 vdd.n2542 vdd.n1035 10.6151
R5028 vdd.n2543 vdd.n2542 10.6151
R5029 vdd.n2544 vdd.n2543 10.6151
R5030 vdd.n2544 vdd.n1024 10.6151
R5031 vdd.n2554 vdd.n1024 10.6151
R5032 vdd.n2555 vdd.n2554 10.6151
R5033 vdd.n2556 vdd.n2555 10.6151
R5034 vdd.n2556 vdd.n1013 10.6151
R5035 vdd.n2566 vdd.n1013 10.6151
R5036 vdd.n2567 vdd.n2566 10.6151
R5037 vdd.n2570 vdd.n2567 10.6151
R5038 vdd.n2570 vdd.n2569 10.6151
R5039 vdd.n2569 vdd.n2568 10.6151
R5040 vdd.n2568 vdd.n996 10.6151
R5041 vdd.n2652 vdd.n996 10.6151
R5042 vdd.n2651 vdd.n2650 10.6151
R5043 vdd.n2650 vdd.n2647 10.6151
R5044 vdd.n2647 vdd.n2646 10.6151
R5045 vdd.n2646 vdd.n2643 10.6151
R5046 vdd.n2643 vdd.n2642 10.6151
R5047 vdd.n2642 vdd.n2639 10.6151
R5048 vdd.n2639 vdd.n2638 10.6151
R5049 vdd.n2638 vdd.n2635 10.6151
R5050 vdd.n2635 vdd.n2634 10.6151
R5051 vdd.n2634 vdd.n2631 10.6151
R5052 vdd.n2631 vdd.n2630 10.6151
R5053 vdd.n2630 vdd.n2627 10.6151
R5054 vdd.n2627 vdd.n2626 10.6151
R5055 vdd.n2626 vdd.n2623 10.6151
R5056 vdd.n2623 vdd.n2622 10.6151
R5057 vdd.n2622 vdd.n2619 10.6151
R5058 vdd.n2619 vdd.n2618 10.6151
R5059 vdd.n2618 vdd.n2615 10.6151
R5060 vdd.n2615 vdd.n2614 10.6151
R5061 vdd.n2614 vdd.n2611 10.6151
R5062 vdd.n2611 vdd.n2610 10.6151
R5063 vdd.n2610 vdd.n2607 10.6151
R5064 vdd.n2607 vdd.n2606 10.6151
R5065 vdd.n2606 vdd.n2603 10.6151
R5066 vdd.n2603 vdd.n2602 10.6151
R5067 vdd.n2602 vdd.n2599 10.6151
R5068 vdd.n2599 vdd.n2598 10.6151
R5069 vdd.n2598 vdd.n2595 10.6151
R5070 vdd.n2595 vdd.n2594 10.6151
R5071 vdd.n2594 vdd.n2591 10.6151
R5072 vdd.n2591 vdd.n2590 10.6151
R5073 vdd.n2587 vdd.n2586 10.6151
R5074 vdd.n2586 vdd.n2584 10.6151
R5075 vdd.n2286 vdd.n2284 10.6151
R5076 vdd.n2287 vdd.n2286 10.6151
R5077 vdd.n2289 vdd.n2287 10.6151
R5078 vdd.n2290 vdd.n2289 10.6151
R5079 vdd.n2292 vdd.n2290 10.6151
R5080 vdd.n2293 vdd.n2292 10.6151
R5081 vdd.n2295 vdd.n2293 10.6151
R5082 vdd.n2296 vdd.n2295 10.6151
R5083 vdd.n2298 vdd.n2296 10.6151
R5084 vdd.n2299 vdd.n2298 10.6151
R5085 vdd.n2301 vdd.n2299 10.6151
R5086 vdd.n2302 vdd.n2301 10.6151
R5087 vdd.n2304 vdd.n2302 10.6151
R5088 vdd.n2305 vdd.n2304 10.6151
R5089 vdd.n2307 vdd.n2305 10.6151
R5090 vdd.n2308 vdd.n2307 10.6151
R5091 vdd.n2310 vdd.n2308 10.6151
R5092 vdd.n2311 vdd.n2310 10.6151
R5093 vdd.n2313 vdd.n2311 10.6151
R5094 vdd.n2314 vdd.n2313 10.6151
R5095 vdd.n2316 vdd.n2314 10.6151
R5096 vdd.n2317 vdd.n2316 10.6151
R5097 vdd.n2356 vdd.n2317 10.6151
R5098 vdd.n2356 vdd.n2355 10.6151
R5099 vdd.n2355 vdd.n2354 10.6151
R5100 vdd.n2354 vdd.n2352 10.6151
R5101 vdd.n2352 vdd.n2351 10.6151
R5102 vdd.n2351 vdd.n2349 10.6151
R5103 vdd.n2349 vdd.n2348 10.6151
R5104 vdd.n2348 vdd.n2325 10.6151
R5105 vdd.n2325 vdd.n2324 10.6151
R5106 vdd.n2324 vdd.n2322 10.6151
R5107 vdd.n2322 vdd.n2321 10.6151
R5108 vdd.n2321 vdd.n2319 10.6151
R5109 vdd.n2319 vdd.n2318 10.6151
R5110 vdd.n2318 vdd.n1000 10.6151
R5111 vdd.n2582 vdd.n1000 10.6151
R5112 vdd.n2583 vdd.n2582 10.6151
R5113 vdd.n2214 vdd.n1108 10.6151
R5114 vdd.n2219 vdd.n2214 10.6151
R5115 vdd.n2220 vdd.n2219 10.6151
R5116 vdd.n2221 vdd.n2220 10.6151
R5117 vdd.n2221 vdd.n2212 10.6151
R5118 vdd.n2227 vdd.n2212 10.6151
R5119 vdd.n2228 vdd.n2227 10.6151
R5120 vdd.n2229 vdd.n2228 10.6151
R5121 vdd.n2229 vdd.n2210 10.6151
R5122 vdd.n2235 vdd.n2210 10.6151
R5123 vdd.n2236 vdd.n2235 10.6151
R5124 vdd.n2237 vdd.n2236 10.6151
R5125 vdd.n2237 vdd.n2208 10.6151
R5126 vdd.n2243 vdd.n2208 10.6151
R5127 vdd.n2244 vdd.n2243 10.6151
R5128 vdd.n2245 vdd.n2244 10.6151
R5129 vdd.n2245 vdd.n2206 10.6151
R5130 vdd.n2251 vdd.n2206 10.6151
R5131 vdd.n2252 vdd.n2251 10.6151
R5132 vdd.n2253 vdd.n2252 10.6151
R5133 vdd.n2253 vdd.n1142 10.6151
R5134 vdd.n2259 vdd.n1142 10.6151
R5135 vdd.n2260 vdd.n2259 10.6151
R5136 vdd.n2261 vdd.n2260 10.6151
R5137 vdd.n2261 vdd.n1140 10.6151
R5138 vdd.n2267 vdd.n1140 10.6151
R5139 vdd.n2268 vdd.n2267 10.6151
R5140 vdd.n2269 vdd.n2268 10.6151
R5141 vdd.n2269 vdd.n1138 10.6151
R5142 vdd.n2275 vdd.n1138 10.6151
R5143 vdd.n2276 vdd.n2275 10.6151
R5144 vdd.n2278 vdd.n1134 10.6151
R5145 vdd.n2283 vdd.n1134 10.6151
R5146 vdd.n1931 vdd.t234 10.5435
R5147 vdd.n656 vdd.t192 10.5435
R5148 vdd.n316 vdd.n298 10.4732
R5149 vdd.n257 vdd.n239 10.4732
R5150 vdd.n214 vdd.n196 10.4732
R5151 vdd.n155 vdd.n137 10.4732
R5152 vdd.n113 vdd.n95 10.4732
R5153 vdd.n54 vdd.n36 10.4732
R5154 vdd.n1815 vdd.n1797 10.4732
R5155 vdd.n1874 vdd.n1856 10.4732
R5156 vdd.n1713 vdd.n1695 10.4732
R5157 vdd.n1772 vdd.n1754 10.4732
R5158 vdd.n1612 vdd.n1594 10.4732
R5159 vdd.n1671 vdd.n1653 10.4732
R5160 vdd.t176 vdd.n1905 10.3167
R5161 vdd.n3482 vdd.t256 10.3167
R5162 vdd.n2654 vdd.t139 10.2034
R5163 vdd.n3017 vdd.t5 10.2034
R5164 vdd.n1582 vdd.t147 10.09
R5165 vdd.n3576 vdd.t210 10.09
R5166 vdd.n2182 vdd.n1122 9.88581
R5167 vdd.n3398 vdd.n731 9.88581
R5168 vdd.n3275 vdd.n3274 9.88581
R5169 vdd.n2206 vdd.n2205 9.88581
R5170 vdd.t141 vdd.n1235 9.86327
R5171 vdd.n3567 vdd.t260 9.86327
R5172 vdd.n315 vdd.n300 9.69747
R5173 vdd.n256 vdd.n241 9.69747
R5174 vdd.n213 vdd.n198 9.69747
R5175 vdd.n154 vdd.n139 9.69747
R5176 vdd.n112 vdd.n97 9.69747
R5177 vdd.n53 vdd.n38 9.69747
R5178 vdd.n1814 vdd.n1799 9.69747
R5179 vdd.n1873 vdd.n1858 9.69747
R5180 vdd.n1712 vdd.n1697 9.69747
R5181 vdd.n1771 vdd.n1756 9.69747
R5182 vdd.n1611 vdd.n1596 9.69747
R5183 vdd.n1670 vdd.n1655 9.69747
R5184 vdd.n1541 vdd.t222 9.63654
R5185 vdd.n3513 vdd.t219 9.63654
R5186 vdd.n331 vdd.n330 9.45567
R5187 vdd.n272 vdd.n271 9.45567
R5188 vdd.n229 vdd.n228 9.45567
R5189 vdd.n170 vdd.n169 9.45567
R5190 vdd.n128 vdd.n127 9.45567
R5191 vdd.n69 vdd.n68 9.45567
R5192 vdd.n1830 vdd.n1829 9.45567
R5193 vdd.n1889 vdd.n1888 9.45567
R5194 vdd.n1728 vdd.n1727 9.45567
R5195 vdd.n1787 vdd.n1786 9.45567
R5196 vdd.n1627 vdd.n1626 9.45567
R5197 vdd.n1686 vdd.n1685 9.45567
R5198 vdd.n1515 vdd.t236 9.40981
R5199 vdd.n3545 vdd.t159 9.40981
R5200 vdd.n2155 vdd.n2009 9.3005
R5201 vdd.n2154 vdd.n2153 9.3005
R5202 vdd.n2015 vdd.n2014 9.3005
R5203 vdd.n2148 vdd.n2019 9.3005
R5204 vdd.n2147 vdd.n2020 9.3005
R5205 vdd.n2146 vdd.n2021 9.3005
R5206 vdd.n2025 vdd.n2022 9.3005
R5207 vdd.n2141 vdd.n2026 9.3005
R5208 vdd.n2140 vdd.n2027 9.3005
R5209 vdd.n2139 vdd.n2028 9.3005
R5210 vdd.n2032 vdd.n2029 9.3005
R5211 vdd.n2134 vdd.n2033 9.3005
R5212 vdd.n2133 vdd.n2034 9.3005
R5213 vdd.n2132 vdd.n2035 9.3005
R5214 vdd.n2039 vdd.n2036 9.3005
R5215 vdd.n2127 vdd.n2040 9.3005
R5216 vdd.n2126 vdd.n2041 9.3005
R5217 vdd.n2125 vdd.n2042 9.3005
R5218 vdd.n2046 vdd.n2043 9.3005
R5219 vdd.n2120 vdd.n2047 9.3005
R5220 vdd.n2119 vdd.n2048 9.3005
R5221 vdd.n2118 vdd.n2117 9.3005
R5222 vdd.n2116 vdd.n2049 9.3005
R5223 vdd.n2115 vdd.n2114 9.3005
R5224 vdd.n2055 vdd.n2054 9.3005
R5225 vdd.n2109 vdd.n2059 9.3005
R5226 vdd.n2108 vdd.n2060 9.3005
R5227 vdd.n2107 vdd.n2061 9.3005
R5228 vdd.n2065 vdd.n2062 9.3005
R5229 vdd.n2102 vdd.n2066 9.3005
R5230 vdd.n2101 vdd.n2067 9.3005
R5231 vdd.n2100 vdd.n2068 9.3005
R5232 vdd.n2072 vdd.n2069 9.3005
R5233 vdd.n2095 vdd.n2073 9.3005
R5234 vdd.n2094 vdd.n2074 9.3005
R5235 vdd.n2093 vdd.n2075 9.3005
R5236 vdd.n2077 vdd.n2076 9.3005
R5237 vdd.n2088 vdd.n1144 9.3005
R5238 vdd.n2157 vdd.n2156 9.3005
R5239 vdd.n2181 vdd.n2180 9.3005
R5240 vdd.n1987 vdd.n1986 9.3005
R5241 vdd.n1992 vdd.n1990 9.3005
R5242 vdd.n2173 vdd.n1993 9.3005
R5243 vdd.n2172 vdd.n1994 9.3005
R5244 vdd.n2171 vdd.n1995 9.3005
R5245 vdd.n1999 vdd.n1996 9.3005
R5246 vdd.n2166 vdd.n2000 9.3005
R5247 vdd.n2165 vdd.n2001 9.3005
R5248 vdd.n2164 vdd.n2002 9.3005
R5249 vdd.n2006 vdd.n2003 9.3005
R5250 vdd.n2159 vdd.n2007 9.3005
R5251 vdd.n2158 vdd.n2008 9.3005
R5252 vdd.n2190 vdd.n1980 9.3005
R5253 vdd.n2192 vdd.n2191 9.3005
R5254 vdd.n1895 vdd.n1894 9.3005
R5255 vdd.n1204 vdd.n1203 9.3005
R5256 vdd.n1909 vdd.n1908 9.3005
R5257 vdd.n1910 vdd.n1202 9.3005
R5258 vdd.n1912 vdd.n1911 9.3005
R5259 vdd.n1193 vdd.n1192 9.3005
R5260 vdd.n1926 vdd.n1925 9.3005
R5261 vdd.n1927 vdd.n1191 9.3005
R5262 vdd.n1929 vdd.n1928 9.3005
R5263 vdd.n1182 vdd.n1181 9.3005
R5264 vdd.n1942 vdd.n1941 9.3005
R5265 vdd.n1943 vdd.n1180 9.3005
R5266 vdd.n1945 vdd.n1944 9.3005
R5267 vdd.n1170 vdd.n1169 9.3005
R5268 vdd.n1959 vdd.n1958 9.3005
R5269 vdd.n1960 vdd.n1168 9.3005
R5270 vdd.n1962 vdd.n1961 9.3005
R5271 vdd.n1158 vdd.n1157 9.3005
R5272 vdd.n1978 vdd.n1977 9.3005
R5273 vdd.n1979 vdd.n1156 9.3005
R5274 vdd.n2194 vdd.n2193 9.3005
R5275 vdd.n307 vdd.n306 9.3005
R5276 vdd.n302 vdd.n301 9.3005
R5277 vdd.n313 vdd.n312 9.3005
R5278 vdd.n315 vdd.n314 9.3005
R5279 vdd.n298 vdd.n297 9.3005
R5280 vdd.n321 vdd.n320 9.3005
R5281 vdd.n323 vdd.n322 9.3005
R5282 vdd.n295 vdd.n292 9.3005
R5283 vdd.n330 vdd.n329 9.3005
R5284 vdd.n248 vdd.n247 9.3005
R5285 vdd.n243 vdd.n242 9.3005
R5286 vdd.n254 vdd.n253 9.3005
R5287 vdd.n256 vdd.n255 9.3005
R5288 vdd.n239 vdd.n238 9.3005
R5289 vdd.n262 vdd.n261 9.3005
R5290 vdd.n264 vdd.n263 9.3005
R5291 vdd.n236 vdd.n233 9.3005
R5292 vdd.n271 vdd.n270 9.3005
R5293 vdd.n205 vdd.n204 9.3005
R5294 vdd.n200 vdd.n199 9.3005
R5295 vdd.n211 vdd.n210 9.3005
R5296 vdd.n213 vdd.n212 9.3005
R5297 vdd.n196 vdd.n195 9.3005
R5298 vdd.n219 vdd.n218 9.3005
R5299 vdd.n221 vdd.n220 9.3005
R5300 vdd.n193 vdd.n190 9.3005
R5301 vdd.n228 vdd.n227 9.3005
R5302 vdd.n146 vdd.n145 9.3005
R5303 vdd.n141 vdd.n140 9.3005
R5304 vdd.n152 vdd.n151 9.3005
R5305 vdd.n154 vdd.n153 9.3005
R5306 vdd.n137 vdd.n136 9.3005
R5307 vdd.n160 vdd.n159 9.3005
R5308 vdd.n162 vdd.n161 9.3005
R5309 vdd.n134 vdd.n131 9.3005
R5310 vdd.n169 vdd.n168 9.3005
R5311 vdd.n104 vdd.n103 9.3005
R5312 vdd.n99 vdd.n98 9.3005
R5313 vdd.n110 vdd.n109 9.3005
R5314 vdd.n112 vdd.n111 9.3005
R5315 vdd.n95 vdd.n94 9.3005
R5316 vdd.n118 vdd.n117 9.3005
R5317 vdd.n120 vdd.n119 9.3005
R5318 vdd.n92 vdd.n89 9.3005
R5319 vdd.n127 vdd.n126 9.3005
R5320 vdd.n45 vdd.n44 9.3005
R5321 vdd.n40 vdd.n39 9.3005
R5322 vdd.n51 vdd.n50 9.3005
R5323 vdd.n53 vdd.n52 9.3005
R5324 vdd.n36 vdd.n35 9.3005
R5325 vdd.n59 vdd.n58 9.3005
R5326 vdd.n61 vdd.n60 9.3005
R5327 vdd.n33 vdd.n30 9.3005
R5328 vdd.n68 vdd.n67 9.3005
R5329 vdd.n3320 vdd.n3319 9.3005
R5330 vdd.n3323 vdd.n766 9.3005
R5331 vdd.n3324 vdd.n765 9.3005
R5332 vdd.n3327 vdd.n764 9.3005
R5333 vdd.n3328 vdd.n763 9.3005
R5334 vdd.n3331 vdd.n762 9.3005
R5335 vdd.n3332 vdd.n761 9.3005
R5336 vdd.n3335 vdd.n760 9.3005
R5337 vdd.n3336 vdd.n759 9.3005
R5338 vdd.n3339 vdd.n758 9.3005
R5339 vdd.n3340 vdd.n757 9.3005
R5340 vdd.n3343 vdd.n756 9.3005
R5341 vdd.n3344 vdd.n755 9.3005
R5342 vdd.n3347 vdd.n754 9.3005
R5343 vdd.n3348 vdd.n753 9.3005
R5344 vdd.n3351 vdd.n752 9.3005
R5345 vdd.n3352 vdd.n751 9.3005
R5346 vdd.n3355 vdd.n750 9.3005
R5347 vdd.n3356 vdd.n749 9.3005
R5348 vdd.n3359 vdd.n748 9.3005
R5349 vdd.n3363 vdd.n3362 9.3005
R5350 vdd.n3364 vdd.n747 9.3005
R5351 vdd.n3368 vdd.n3365 9.3005
R5352 vdd.n3371 vdd.n746 9.3005
R5353 vdd.n3372 vdd.n745 9.3005
R5354 vdd.n3375 vdd.n744 9.3005
R5355 vdd.n3376 vdd.n743 9.3005
R5356 vdd.n3379 vdd.n742 9.3005
R5357 vdd.n3380 vdd.n741 9.3005
R5358 vdd.n3383 vdd.n740 9.3005
R5359 vdd.n3384 vdd.n739 9.3005
R5360 vdd.n3387 vdd.n738 9.3005
R5361 vdd.n3388 vdd.n737 9.3005
R5362 vdd.n3391 vdd.n736 9.3005
R5363 vdd.n3392 vdd.n735 9.3005
R5364 vdd.n3395 vdd.n730 9.3005
R5365 vdd.n3401 vdd.n727 9.3005
R5366 vdd.n3402 vdd.n726 9.3005
R5367 vdd.n3416 vdd.n3415 9.3005
R5368 vdd.n3417 vdd.n681 9.3005
R5369 vdd.n3419 vdd.n3418 9.3005
R5370 vdd.n671 vdd.n670 9.3005
R5371 vdd.n3433 vdd.n3432 9.3005
R5372 vdd.n3434 vdd.n669 9.3005
R5373 vdd.n3436 vdd.n3435 9.3005
R5374 vdd.n660 vdd.n659 9.3005
R5375 vdd.n3449 vdd.n3448 9.3005
R5376 vdd.n3450 vdd.n658 9.3005
R5377 vdd.n3452 vdd.n3451 9.3005
R5378 vdd.n648 vdd.n647 9.3005
R5379 vdd.n3466 vdd.n3465 9.3005
R5380 vdd.n3467 vdd.n646 9.3005
R5381 vdd.n3469 vdd.n3468 9.3005
R5382 vdd.n637 vdd.n636 9.3005
R5383 vdd.n3485 vdd.n3484 9.3005
R5384 vdd.n3486 vdd.n635 9.3005
R5385 vdd.n3488 vdd.n3487 9.3005
R5386 vdd.n336 vdd.n334 9.3005
R5387 vdd.n683 vdd.n682 9.3005
R5388 vdd.n3580 vdd.n3579 9.3005
R5389 vdd.n337 vdd.n335 9.3005
R5390 vdd.n3573 vdd.n346 9.3005
R5391 vdd.n3572 vdd.n347 9.3005
R5392 vdd.n3571 vdd.n348 9.3005
R5393 vdd.n355 vdd.n349 9.3005
R5394 vdd.n3565 vdd.n356 9.3005
R5395 vdd.n3564 vdd.n357 9.3005
R5396 vdd.n3563 vdd.n358 9.3005
R5397 vdd.n366 vdd.n359 9.3005
R5398 vdd.n3557 vdd.n367 9.3005
R5399 vdd.n3556 vdd.n368 9.3005
R5400 vdd.n3555 vdd.n369 9.3005
R5401 vdd.n377 vdd.n370 9.3005
R5402 vdd.n3549 vdd.n378 9.3005
R5403 vdd.n3548 vdd.n379 9.3005
R5404 vdd.n3547 vdd.n380 9.3005
R5405 vdd.n388 vdd.n381 9.3005
R5406 vdd.n3541 vdd.n389 9.3005
R5407 vdd.n3540 vdd.n390 9.3005
R5408 vdd.n3539 vdd.n391 9.3005
R5409 vdd.n466 vdd.n463 9.3005
R5410 vdd.n470 vdd.n469 9.3005
R5411 vdd.n471 vdd.n462 9.3005
R5412 vdd.n475 vdd.n472 9.3005
R5413 vdd.n476 vdd.n461 9.3005
R5414 vdd.n480 vdd.n479 9.3005
R5415 vdd.n481 vdd.n460 9.3005
R5416 vdd.n485 vdd.n482 9.3005
R5417 vdd.n486 vdd.n459 9.3005
R5418 vdd.n490 vdd.n489 9.3005
R5419 vdd.n491 vdd.n458 9.3005
R5420 vdd.n495 vdd.n492 9.3005
R5421 vdd.n496 vdd.n457 9.3005
R5422 vdd.n500 vdd.n499 9.3005
R5423 vdd.n501 vdd.n456 9.3005
R5424 vdd.n505 vdd.n502 9.3005
R5425 vdd.n506 vdd.n455 9.3005
R5426 vdd.n510 vdd.n509 9.3005
R5427 vdd.n511 vdd.n454 9.3005
R5428 vdd.n515 vdd.n512 9.3005
R5429 vdd.n516 vdd.n451 9.3005
R5430 vdd.n520 vdd.n519 9.3005
R5431 vdd.n521 vdd.n450 9.3005
R5432 vdd.n525 vdd.n522 9.3005
R5433 vdd.n526 vdd.n449 9.3005
R5434 vdd.n530 vdd.n529 9.3005
R5435 vdd.n531 vdd.n448 9.3005
R5436 vdd.n535 vdd.n532 9.3005
R5437 vdd.n536 vdd.n447 9.3005
R5438 vdd.n540 vdd.n539 9.3005
R5439 vdd.n541 vdd.n446 9.3005
R5440 vdd.n545 vdd.n542 9.3005
R5441 vdd.n546 vdd.n445 9.3005
R5442 vdd.n550 vdd.n549 9.3005
R5443 vdd.n551 vdd.n444 9.3005
R5444 vdd.n555 vdd.n552 9.3005
R5445 vdd.n556 vdd.n443 9.3005
R5446 vdd.n560 vdd.n559 9.3005
R5447 vdd.n561 vdd.n442 9.3005
R5448 vdd.n565 vdd.n562 9.3005
R5449 vdd.n566 vdd.n439 9.3005
R5450 vdd.n570 vdd.n569 9.3005
R5451 vdd.n571 vdd.n438 9.3005
R5452 vdd.n575 vdd.n572 9.3005
R5453 vdd.n576 vdd.n437 9.3005
R5454 vdd.n580 vdd.n579 9.3005
R5455 vdd.n581 vdd.n436 9.3005
R5456 vdd.n585 vdd.n582 9.3005
R5457 vdd.n586 vdd.n435 9.3005
R5458 vdd.n590 vdd.n589 9.3005
R5459 vdd.n591 vdd.n434 9.3005
R5460 vdd.n595 vdd.n592 9.3005
R5461 vdd.n596 vdd.n433 9.3005
R5462 vdd.n600 vdd.n599 9.3005
R5463 vdd.n601 vdd.n432 9.3005
R5464 vdd.n605 vdd.n602 9.3005
R5465 vdd.n606 vdd.n431 9.3005
R5466 vdd.n610 vdd.n609 9.3005
R5467 vdd.n611 vdd.n430 9.3005
R5468 vdd.n615 vdd.n612 9.3005
R5469 vdd.n617 vdd.n429 9.3005
R5470 vdd.n619 vdd.n618 9.3005
R5471 vdd.n3533 vdd.n3532 9.3005
R5472 vdd.n465 vdd.n464 9.3005
R5473 vdd.n3411 vdd.n3410 9.3005
R5474 vdd.n676 vdd.n675 9.3005
R5475 vdd.n3424 vdd.n3423 9.3005
R5476 vdd.n3425 vdd.n674 9.3005
R5477 vdd.n3427 vdd.n3426 9.3005
R5478 vdd.n666 vdd.n665 9.3005
R5479 vdd.n3441 vdd.n3440 9.3005
R5480 vdd.n3442 vdd.n664 9.3005
R5481 vdd.n3444 vdd.n3443 9.3005
R5482 vdd.n653 vdd.n652 9.3005
R5483 vdd.n3457 vdd.n3456 9.3005
R5484 vdd.n3458 vdd.n651 9.3005
R5485 vdd.n3460 vdd.n3459 9.3005
R5486 vdd.n642 vdd.n641 9.3005
R5487 vdd.n3474 vdd.n3473 9.3005
R5488 vdd.n3475 vdd.n640 9.3005
R5489 vdd.n3480 vdd.n3476 9.3005
R5490 vdd.n3479 vdd.n3478 9.3005
R5491 vdd.n3477 vdd.n631 9.3005
R5492 vdd.n3493 vdd.n630 9.3005
R5493 vdd.n3495 vdd.n3494 9.3005
R5494 vdd.n3496 vdd.n629 9.3005
R5495 vdd.n3498 vdd.n3497 9.3005
R5496 vdd.n3500 vdd.n628 9.3005
R5497 vdd.n3502 vdd.n3501 9.3005
R5498 vdd.n3503 vdd.n627 9.3005
R5499 vdd.n3505 vdd.n3504 9.3005
R5500 vdd.n3507 vdd.n626 9.3005
R5501 vdd.n3509 vdd.n3508 9.3005
R5502 vdd.n3510 vdd.n625 9.3005
R5503 vdd.n3512 vdd.n3511 9.3005
R5504 vdd.n3515 vdd.n624 9.3005
R5505 vdd.n3517 vdd.n3516 9.3005
R5506 vdd.n3518 vdd.n623 9.3005
R5507 vdd.n3520 vdd.n3519 9.3005
R5508 vdd.n3522 vdd.n622 9.3005
R5509 vdd.n3524 vdd.n3523 9.3005
R5510 vdd.n3525 vdd.n621 9.3005
R5511 vdd.n3527 vdd.n3526 9.3005
R5512 vdd.n3529 vdd.n620 9.3005
R5513 vdd.n3531 vdd.n3530 9.3005
R5514 vdd.n3409 vdd.n686 9.3005
R5515 vdd.n3408 vdd.n3407 9.3005
R5516 vdd.n3277 vdd.n687 9.3005
R5517 vdd.n3286 vdd.n783 9.3005
R5518 vdd.n3289 vdd.n782 9.3005
R5519 vdd.n3290 vdd.n781 9.3005
R5520 vdd.n3293 vdd.n780 9.3005
R5521 vdd.n3294 vdd.n779 9.3005
R5522 vdd.n3297 vdd.n778 9.3005
R5523 vdd.n3298 vdd.n777 9.3005
R5524 vdd.n3301 vdd.n776 9.3005
R5525 vdd.n3302 vdd.n775 9.3005
R5526 vdd.n3305 vdd.n774 9.3005
R5527 vdd.n3306 vdd.n773 9.3005
R5528 vdd.n3309 vdd.n772 9.3005
R5529 vdd.n3310 vdd.n771 9.3005
R5530 vdd.n3313 vdd.n770 9.3005
R5531 vdd.n3317 vdd.n3316 9.3005
R5532 vdd.n3318 vdd.n767 9.3005
R5533 vdd.n2204 vdd.n2203 9.3005
R5534 vdd.n2199 vdd.n1147 9.3005
R5535 vdd.n1510 vdd.n1509 9.3005
R5536 vdd.n1511 vdd.n1265 9.3005
R5537 vdd.n1513 vdd.n1512 9.3005
R5538 vdd.n1255 vdd.n1254 9.3005
R5539 vdd.n1527 vdd.n1526 9.3005
R5540 vdd.n1528 vdd.n1253 9.3005
R5541 vdd.n1530 vdd.n1529 9.3005
R5542 vdd.n1245 vdd.n1244 9.3005
R5543 vdd.n1544 vdd.n1543 9.3005
R5544 vdd.n1545 vdd.n1243 9.3005
R5545 vdd.n1547 vdd.n1546 9.3005
R5546 vdd.n1232 vdd.n1231 9.3005
R5547 vdd.n1560 vdd.n1559 9.3005
R5548 vdd.n1561 vdd.n1230 9.3005
R5549 vdd.n1563 vdd.n1562 9.3005
R5550 vdd.n1221 vdd.n1220 9.3005
R5551 vdd.n1577 vdd.n1576 9.3005
R5552 vdd.n1578 vdd.n1219 9.3005
R5553 vdd.n1580 vdd.n1579 9.3005
R5554 vdd.n1210 vdd.n1209 9.3005
R5555 vdd.n1900 vdd.n1899 9.3005
R5556 vdd.n1901 vdd.n1208 9.3005
R5557 vdd.n1903 vdd.n1902 9.3005
R5558 vdd.n1198 vdd.n1197 9.3005
R5559 vdd.n1917 vdd.n1916 9.3005
R5560 vdd.n1918 vdd.n1196 9.3005
R5561 vdd.n1920 vdd.n1919 9.3005
R5562 vdd.n1188 vdd.n1187 9.3005
R5563 vdd.n1934 vdd.n1933 9.3005
R5564 vdd.n1935 vdd.n1186 9.3005
R5565 vdd.n1937 vdd.n1936 9.3005
R5566 vdd.n1175 vdd.n1174 9.3005
R5567 vdd.n1950 vdd.n1949 9.3005
R5568 vdd.n1951 vdd.n1173 9.3005
R5569 vdd.n1953 vdd.n1952 9.3005
R5570 vdd.n1165 vdd.n1164 9.3005
R5571 vdd.n1967 vdd.n1966 9.3005
R5572 vdd.n1968 vdd.n1162 9.3005
R5573 vdd.n1972 vdd.n1971 9.3005
R5574 vdd.n1970 vdd.n1163 9.3005
R5575 vdd.n1969 vdd.n1152 9.3005
R5576 vdd.n1267 vdd.n1266 9.3005
R5577 vdd.n1403 vdd.n1402 9.3005
R5578 vdd.n1404 vdd.n1393 9.3005
R5579 vdd.n1406 vdd.n1405 9.3005
R5580 vdd.n1407 vdd.n1392 9.3005
R5581 vdd.n1409 vdd.n1408 9.3005
R5582 vdd.n1410 vdd.n1387 9.3005
R5583 vdd.n1412 vdd.n1411 9.3005
R5584 vdd.n1413 vdd.n1386 9.3005
R5585 vdd.n1415 vdd.n1414 9.3005
R5586 vdd.n1416 vdd.n1381 9.3005
R5587 vdd.n1418 vdd.n1417 9.3005
R5588 vdd.n1419 vdd.n1380 9.3005
R5589 vdd.n1421 vdd.n1420 9.3005
R5590 vdd.n1422 vdd.n1375 9.3005
R5591 vdd.n1424 vdd.n1423 9.3005
R5592 vdd.n1425 vdd.n1374 9.3005
R5593 vdd.n1427 vdd.n1426 9.3005
R5594 vdd.n1428 vdd.n1369 9.3005
R5595 vdd.n1430 vdd.n1429 9.3005
R5596 vdd.n1431 vdd.n1368 9.3005
R5597 vdd.n1433 vdd.n1432 9.3005
R5598 vdd.n1437 vdd.n1364 9.3005
R5599 vdd.n1439 vdd.n1438 9.3005
R5600 vdd.n1440 vdd.n1363 9.3005
R5601 vdd.n1442 vdd.n1441 9.3005
R5602 vdd.n1443 vdd.n1358 9.3005
R5603 vdd.n1445 vdd.n1444 9.3005
R5604 vdd.n1446 vdd.n1357 9.3005
R5605 vdd.n1448 vdd.n1447 9.3005
R5606 vdd.n1449 vdd.n1352 9.3005
R5607 vdd.n1451 vdd.n1450 9.3005
R5608 vdd.n1452 vdd.n1351 9.3005
R5609 vdd.n1454 vdd.n1453 9.3005
R5610 vdd.n1455 vdd.n1346 9.3005
R5611 vdd.n1457 vdd.n1456 9.3005
R5612 vdd.n1458 vdd.n1345 9.3005
R5613 vdd.n1460 vdd.n1459 9.3005
R5614 vdd.n1461 vdd.n1340 9.3005
R5615 vdd.n1463 vdd.n1462 9.3005
R5616 vdd.n1464 vdd.n1339 9.3005
R5617 vdd.n1466 vdd.n1465 9.3005
R5618 vdd.n1467 vdd.n1334 9.3005
R5619 vdd.n1469 vdd.n1468 9.3005
R5620 vdd.n1470 vdd.n1333 9.3005
R5621 vdd.n1472 vdd.n1471 9.3005
R5622 vdd.n1473 vdd.n1326 9.3005
R5623 vdd.n1475 vdd.n1474 9.3005
R5624 vdd.n1476 vdd.n1325 9.3005
R5625 vdd.n1478 vdd.n1477 9.3005
R5626 vdd.n1479 vdd.n1320 9.3005
R5627 vdd.n1481 vdd.n1480 9.3005
R5628 vdd.n1482 vdd.n1319 9.3005
R5629 vdd.n1484 vdd.n1483 9.3005
R5630 vdd.n1485 vdd.n1314 9.3005
R5631 vdd.n1487 vdd.n1486 9.3005
R5632 vdd.n1488 vdd.n1313 9.3005
R5633 vdd.n1490 vdd.n1489 9.3005
R5634 vdd.n1491 vdd.n1308 9.3005
R5635 vdd.n1493 vdd.n1492 9.3005
R5636 vdd.n1494 vdd.n1307 9.3005
R5637 vdd.n1496 vdd.n1495 9.3005
R5638 vdd.n1272 vdd.n1271 9.3005
R5639 vdd.n1502 vdd.n1501 9.3005
R5640 vdd.n1401 vdd.n1400 9.3005
R5641 vdd.n1505 vdd.n1504 9.3005
R5642 vdd.n1261 vdd.n1260 9.3005
R5643 vdd.n1519 vdd.n1518 9.3005
R5644 vdd.n1520 vdd.n1259 9.3005
R5645 vdd.n1522 vdd.n1521 9.3005
R5646 vdd.n1250 vdd.n1249 9.3005
R5647 vdd.n1536 vdd.n1535 9.3005
R5648 vdd.n1537 vdd.n1248 9.3005
R5649 vdd.n1539 vdd.n1538 9.3005
R5650 vdd.n1239 vdd.n1238 9.3005
R5651 vdd.n1552 vdd.n1551 9.3005
R5652 vdd.n1553 vdd.n1237 9.3005
R5653 vdd.n1555 vdd.n1554 9.3005
R5654 vdd.n1227 vdd.n1226 9.3005
R5655 vdd.n1569 vdd.n1568 9.3005
R5656 vdd.n1570 vdd.n1225 9.3005
R5657 vdd.n1572 vdd.n1571 9.3005
R5658 vdd.n1216 vdd.n1215 9.3005
R5659 vdd.n1585 vdd.n1584 9.3005
R5660 vdd.n1586 vdd.n1214 9.3005
R5661 vdd.n1503 vdd.n1270 9.3005
R5662 vdd.n1806 vdd.n1805 9.3005
R5663 vdd.n1801 vdd.n1800 9.3005
R5664 vdd.n1812 vdd.n1811 9.3005
R5665 vdd.n1814 vdd.n1813 9.3005
R5666 vdd.n1797 vdd.n1796 9.3005
R5667 vdd.n1820 vdd.n1819 9.3005
R5668 vdd.n1822 vdd.n1821 9.3005
R5669 vdd.n1794 vdd.n1791 9.3005
R5670 vdd.n1829 vdd.n1828 9.3005
R5671 vdd.n1865 vdd.n1864 9.3005
R5672 vdd.n1860 vdd.n1859 9.3005
R5673 vdd.n1871 vdd.n1870 9.3005
R5674 vdd.n1873 vdd.n1872 9.3005
R5675 vdd.n1856 vdd.n1855 9.3005
R5676 vdd.n1879 vdd.n1878 9.3005
R5677 vdd.n1881 vdd.n1880 9.3005
R5678 vdd.n1853 vdd.n1850 9.3005
R5679 vdd.n1888 vdd.n1887 9.3005
R5680 vdd.n1704 vdd.n1703 9.3005
R5681 vdd.n1699 vdd.n1698 9.3005
R5682 vdd.n1710 vdd.n1709 9.3005
R5683 vdd.n1712 vdd.n1711 9.3005
R5684 vdd.n1695 vdd.n1694 9.3005
R5685 vdd.n1718 vdd.n1717 9.3005
R5686 vdd.n1720 vdd.n1719 9.3005
R5687 vdd.n1692 vdd.n1689 9.3005
R5688 vdd.n1727 vdd.n1726 9.3005
R5689 vdd.n1763 vdd.n1762 9.3005
R5690 vdd.n1758 vdd.n1757 9.3005
R5691 vdd.n1769 vdd.n1768 9.3005
R5692 vdd.n1771 vdd.n1770 9.3005
R5693 vdd.n1754 vdd.n1753 9.3005
R5694 vdd.n1777 vdd.n1776 9.3005
R5695 vdd.n1779 vdd.n1778 9.3005
R5696 vdd.n1751 vdd.n1748 9.3005
R5697 vdd.n1786 vdd.n1785 9.3005
R5698 vdd.n1603 vdd.n1602 9.3005
R5699 vdd.n1598 vdd.n1597 9.3005
R5700 vdd.n1609 vdd.n1608 9.3005
R5701 vdd.n1611 vdd.n1610 9.3005
R5702 vdd.n1594 vdd.n1593 9.3005
R5703 vdd.n1617 vdd.n1616 9.3005
R5704 vdd.n1619 vdd.n1618 9.3005
R5705 vdd.n1591 vdd.n1588 9.3005
R5706 vdd.n1626 vdd.n1625 9.3005
R5707 vdd.n1662 vdd.n1661 9.3005
R5708 vdd.n1657 vdd.n1656 9.3005
R5709 vdd.n1668 vdd.n1667 9.3005
R5710 vdd.n1670 vdd.n1669 9.3005
R5711 vdd.n1653 vdd.n1652 9.3005
R5712 vdd.n1676 vdd.n1675 9.3005
R5713 vdd.n1678 vdd.n1677 9.3005
R5714 vdd.n1650 vdd.n1647 9.3005
R5715 vdd.n1685 vdd.n1684 9.3005
R5716 vdd.n1541 vdd.t253 9.18308
R5717 vdd.n3513 vdd.t189 9.18308
R5718 vdd.n1235 vdd.t232 8.95635
R5719 vdd.n2196 vdd.t48 8.95635
R5720 vdd.n723 vdd.t22 8.95635
R5721 vdd.t198 vdd.n3567 8.95635
R5722 vdd.n312 vdd.n311 8.92171
R5723 vdd.n253 vdd.n252 8.92171
R5724 vdd.n210 vdd.n209 8.92171
R5725 vdd.n151 vdd.n150 8.92171
R5726 vdd.n109 vdd.n108 8.92171
R5727 vdd.n50 vdd.n49 8.92171
R5728 vdd.n1811 vdd.n1810 8.92171
R5729 vdd.n1870 vdd.n1869 8.92171
R5730 vdd.n1709 vdd.n1708 8.92171
R5731 vdd.n1768 vdd.n1767 8.92171
R5732 vdd.n1608 vdd.n1607 8.92171
R5733 vdd.n1667 vdd.n1666 8.92171
R5734 vdd.n231 vdd.n129 8.81535
R5735 vdd.n1789 vdd.n1687 8.81535
R5736 vdd.n1582 vdd.t143 8.72962
R5737 vdd.t225 vdd.n3576 8.72962
R5738 vdd.n1905 vdd.t151 8.50289
R5739 vdd.n3482 vdd.t168 8.50289
R5740 vdd.n28 vdd.n14 8.42249
R5741 vdd.n1931 vdd.t181 8.27616
R5742 vdd.t227 vdd.n656 8.27616
R5743 vdd.n3582 vdd.n3581 8.16225
R5744 vdd.n1893 vdd.n1892 8.16225
R5745 vdd.n308 vdd.n302 8.14595
R5746 vdd.n249 vdd.n243 8.14595
R5747 vdd.n206 vdd.n200 8.14595
R5748 vdd.n147 vdd.n141 8.14595
R5749 vdd.n105 vdd.n99 8.14595
R5750 vdd.n46 vdd.n40 8.14595
R5751 vdd.n1807 vdd.n1801 8.14595
R5752 vdd.n1866 vdd.n1860 8.14595
R5753 vdd.n1705 vdd.n1699 8.14595
R5754 vdd.n1764 vdd.n1758 8.14595
R5755 vdd.n1604 vdd.n1598 8.14595
R5756 vdd.n1663 vdd.n1657 8.14595
R5757 vdd.n1178 vdd.t153 8.04943
R5758 vdd.n3438 vdd.t149 8.04943
R5759 vdd.n2467 vdd.n1104 7.70933
R5760 vdd.n2473 vdd.n1104 7.70933
R5761 vdd.n2479 vdd.n1098 7.70933
R5762 vdd.n2479 vdd.n1092 7.70933
R5763 vdd.n2485 vdd.n1092 7.70933
R5764 vdd.n2485 vdd.n1086 7.70933
R5765 vdd.n2491 vdd.n1086 7.70933
R5766 vdd.n2497 vdd.n1080 7.70933
R5767 vdd.n2503 vdd.n1074 7.70933
R5768 vdd.n2509 vdd.n1067 7.70933
R5769 vdd.n2509 vdd.n1070 7.70933
R5770 vdd.n2515 vdd.n1063 7.70933
R5771 vdd.n2522 vdd.n1049 7.70933
R5772 vdd.n2528 vdd.n1049 7.70933
R5773 vdd.n2534 vdd.n1043 7.70933
R5774 vdd.n2540 vdd.n1039 7.70933
R5775 vdd.n2546 vdd.n1033 7.70933
R5776 vdd.n2564 vdd.n1015 7.70933
R5777 vdd.n2564 vdd.n1008 7.70933
R5778 vdd.n2572 vdd.n1008 7.70933
R5779 vdd.n2654 vdd.n992 7.70933
R5780 vdd.n3017 vdd.n946 7.70933
R5781 vdd.n3029 vdd.n927 7.70933
R5782 vdd.n3035 vdd.n927 7.70933
R5783 vdd.n3035 vdd.n930 7.70933
R5784 vdd.n3053 vdd.n911 7.70933
R5785 vdd.n3059 vdd.n905 7.70933
R5786 vdd.n3065 vdd.n901 7.70933
R5787 vdd.n3071 vdd.n888 7.70933
R5788 vdd.n3077 vdd.n888 7.70933
R5789 vdd.n3084 vdd.n881 7.70933
R5790 vdd.n3090 vdd.n874 7.70933
R5791 vdd.n3090 vdd.n877 7.70933
R5792 vdd.n3096 vdd.n870 7.70933
R5793 vdd.n3102 vdd.n864 7.70933
R5794 vdd.n3108 vdd.n851 7.70933
R5795 vdd.n3114 vdd.n851 7.70933
R5796 vdd.n3114 vdd.n843 7.70933
R5797 vdd.n3165 vdd.n843 7.70933
R5798 vdd.n3165 vdd.n846 7.70933
R5799 vdd.n3171 vdd.n805 7.70933
R5800 vdd.n3241 vdd.n805 7.70933
R5801 vdd.t117 vdd.n1080 7.59597
R5802 vdd.n2346 vdd.t131 7.59597
R5803 vdd.n2989 vdd.t0 7.59597
R5804 vdd.n864 vdd.t9 7.59597
R5805 vdd.n307 vdd.n304 7.3702
R5806 vdd.n248 vdd.n245 7.3702
R5807 vdd.n205 vdd.n202 7.3702
R5808 vdd.n146 vdd.n143 7.3702
R5809 vdd.n104 vdd.n101 7.3702
R5810 vdd.n45 vdd.n42 7.3702
R5811 vdd.n1806 vdd.n1803 7.3702
R5812 vdd.n1865 vdd.n1862 7.3702
R5813 vdd.n1704 vdd.n1701 7.3702
R5814 vdd.n1763 vdd.n1760 7.3702
R5815 vdd.n1603 vdd.n1600 7.3702
R5816 vdd.n1662 vdd.n1659 7.3702
R5817 vdd.n1964 vdd.t240 7.1425
R5818 vdd.n679 vdd.t200 7.1425
R5819 vdd.n1438 vdd.n1437 6.98232
R5820 vdd.n2119 vdd.n2118 6.98232
R5821 vdd.n566 vdd.n565 6.98232
R5822 vdd.n3323 vdd.n3320 6.98232
R5823 vdd.t166 vdd.n1177 6.91577
R5824 vdd.n2503 vdd.t130 6.91577
R5825 vdd.n3096 vdd.t7 6.91577
R5826 vdd.n3446 vdd.t163 6.91577
R5827 vdd.n3081 vdd.n3080 6.86879
R5828 vdd.n2519 vdd.n2518 6.86879
R5829 vdd.n2579 vdd.t137 6.80241
R5830 vdd.n3023 vdd.t3 6.80241
R5831 vdd.n1923 vdd.t238 6.68904
R5832 vdd.n3462 vdd.t161 6.68904
R5833 vdd.t178 vdd.n1206 6.46231
R5834 vdd.n3490 vdd.t155 6.46231
R5835 vdd.n3582 vdd.n333 6.38151
R5836 vdd.n1892 vdd.n1891 6.38151
R5837 vdd.n2346 vdd.t1 6.34895
R5838 vdd.n2989 vdd.t107 6.34895
R5839 vdd.n1574 vdd.t206 6.23558
R5840 vdd.t145 vdd.n344 6.23558
R5841 vdd.t194 vdd.n1234 6.00885
R5842 vdd.t11 vdd.n1043 6.00885
R5843 vdd.n901 vdd.t14 6.00885
R5844 vdd.n3561 vdd.t157 6.00885
R5845 vdd.n308 vdd.n307 5.81868
R5846 vdd.n249 vdd.n248 5.81868
R5847 vdd.n206 vdd.n205 5.81868
R5848 vdd.n147 vdd.n146 5.81868
R5849 vdd.n105 vdd.n104 5.81868
R5850 vdd.n46 vdd.n45 5.81868
R5851 vdd.n1807 vdd.n1806 5.81868
R5852 vdd.n1866 vdd.n1865 5.81868
R5853 vdd.n1705 vdd.n1704 5.81868
R5854 vdd.n1764 vdd.n1763 5.81868
R5855 vdd.n1604 vdd.n1603 5.81868
R5856 vdd.n1663 vdd.n1662 5.81868
R5857 vdd.n1533 vdd.t183 5.78212
R5858 vdd.n3552 vdd.t280 5.78212
R5859 vdd.n2662 vdd.n2661 5.77611
R5860 vdd.n2402 vdd.n2401 5.77611
R5861 vdd.n2891 vdd.n2890 5.77611
R5862 vdd.n3182 vdd.n3181 5.77611
R5863 vdd.n3246 vdd.n801 5.77611
R5864 vdd.n2827 vdd.n2763 5.77611
R5865 vdd.n2587 vdd.n999 5.77611
R5866 vdd.n2278 vdd.n2277 5.77611
R5867 vdd.n1400 vdd.n1399 5.62474
R5868 vdd.n2202 vdd.n2199 5.62474
R5869 vdd.n3533 vdd.n428 5.62474
R5870 vdd.n3407 vdd.n690 5.62474
R5871 vdd.n1257 vdd.t183 5.55539
R5872 vdd.t280 vdd.n3551 5.55539
R5873 vdd.n2540 vdd.t109 5.44203
R5874 vdd.n3059 vdd.t120 5.44203
R5875 vdd.n1549 vdd.t194 5.32866
R5876 vdd.t157 vdd.n3560 5.32866
R5877 vdd.n1565 vdd.t206 5.10193
R5878 vdd.n2515 vdd.t8 5.10193
R5879 vdd.n2534 vdd.t124 5.10193
R5880 vdd.n3065 vdd.t15 5.10193
R5881 vdd.n3084 vdd.t114 5.10193
R5882 vdd.n3569 vdd.t145 5.10193
R5883 vdd.n311 vdd.n302 5.04292
R5884 vdd.n252 vdd.n243 5.04292
R5885 vdd.n209 vdd.n200 5.04292
R5886 vdd.n150 vdd.n141 5.04292
R5887 vdd.n108 vdd.n99 5.04292
R5888 vdd.n49 vdd.n40 5.04292
R5889 vdd.n1810 vdd.n1801 5.04292
R5890 vdd.n1869 vdd.n1860 5.04292
R5891 vdd.n1708 vdd.n1699 5.04292
R5892 vdd.n1767 vdd.n1758 5.04292
R5893 vdd.n1607 vdd.n1598 5.04292
R5894 vdd.n1666 vdd.n1657 5.04292
R5895 vdd.n1063 vdd.t82 4.98857
R5896 vdd.t41 vdd.n881 4.98857
R5897 vdd.n1897 vdd.t178 4.8752
R5898 vdd.t30 vdd.n1098 4.8752
R5899 vdd.t105 vdd.t103 4.8752
R5900 vdd.n2334 vdd.t68 4.8752
R5901 vdd.n3001 vdd.t72 4.8752
R5902 vdd.t122 vdd.t127 4.8752
R5903 vdd.n846 vdd.t26 4.8752
R5904 vdd.t155 vdd.n340 4.8752
R5905 vdd.n2663 vdd.n2662 4.83952
R5906 vdd.n2403 vdd.n2402 4.83952
R5907 vdd.n2890 vdd.n2889 4.83952
R5908 vdd.n3183 vdd.n3182 4.83952
R5909 vdd.n801 vdd.n796 4.83952
R5910 vdd.n2824 vdd.n2763 4.83952
R5911 vdd.n2590 vdd.n999 4.83952
R5912 vdd.n2277 vdd.n2276 4.83952
R5913 vdd.n2558 vdd.t302 4.76184
R5914 vdd.n3041 vdd.t101 4.76184
R5915 vdd.n2087 vdd.n1145 4.74817
R5916 vdd.n2082 vdd.n1146 4.74817
R5917 vdd.n1984 vdd.n1981 4.74817
R5918 vdd.n2183 vdd.n1985 4.74817
R5919 vdd.n2185 vdd.n1984 4.74817
R5920 vdd.n2184 vdd.n2183 4.74817
R5921 vdd.n3400 vdd.n3399 4.74817
R5922 vdd.n3397 vdd.n3396 4.74817
R5923 vdd.n3397 vdd.n732 4.74817
R5924 vdd.n3399 vdd.n729 4.74817
R5925 vdd.n3282 vdd.n784 4.74817
R5926 vdd.n3278 vdd.n3276 4.74817
R5927 vdd.n3281 vdd.n3276 4.74817
R5928 vdd.n3285 vdd.n784 4.74817
R5929 vdd.n2083 vdd.n1145 4.74817
R5930 vdd.n1148 vdd.n1146 4.74817
R5931 vdd.n333 vdd.n332 4.7074
R5932 vdd.n231 vdd.n230 4.7074
R5933 vdd.n1891 vdd.n1890 4.7074
R5934 vdd.n1789 vdd.n1788 4.7074
R5935 vdd.n1200 vdd.t238 4.64847
R5936 vdd.n3471 vdd.t161 4.64847
R5937 vdd.n1939 vdd.t166 4.42174
R5938 vdd.t163 vdd.n655 4.42174
R5939 vdd.n2334 vdd.t118 4.30838
R5940 vdd.n3001 vdd.t132 4.30838
R5941 vdd.n312 vdd.n300 4.26717
R5942 vdd.n253 vdd.n241 4.26717
R5943 vdd.n210 vdd.n198 4.26717
R5944 vdd.n151 vdd.n139 4.26717
R5945 vdd.n109 vdd.n97 4.26717
R5946 vdd.n50 vdd.n38 4.26717
R5947 vdd.n1811 vdd.n1799 4.26717
R5948 vdd.n1870 vdd.n1858 4.26717
R5949 vdd.n1709 vdd.n1697 4.26717
R5950 vdd.n1768 vdd.n1756 4.26717
R5951 vdd.n1608 vdd.n1596 4.26717
R5952 vdd.n1667 vdd.n1655 4.26717
R5953 vdd.n1955 vdd.t240 4.19501
R5954 vdd.t19 vdd.n1074 4.19501
R5955 vdd.n1033 vdd.t20 4.19501
R5956 vdd.t106 vdd.n911 4.19501
R5957 vdd.n870 vdd.t111 4.19501
R5958 vdd.n3430 vdd.t200 4.19501
R5959 vdd.n333 vdd.n231 4.10845
R5960 vdd.n1891 vdd.n1789 4.10845
R5961 vdd.n289 vdd.t251 4.06363
R5962 vdd.n289 vdd.t292 4.06363
R5963 vdd.n287 vdd.t158 4.06363
R5964 vdd.n287 vdd.t215 4.06363
R5965 vdd.n285 vdd.t218 4.06363
R5966 vdd.n285 vdd.t271 4.06363
R5967 vdd.n283 vdd.t273 4.06363
R5968 vdd.n283 vdd.t146 4.06363
R5969 vdd.n281 vdd.t175 4.06363
R5970 vdd.n281 vdd.t245 4.06363
R5971 vdd.n279 vdd.t274 4.06363
R5972 vdd.n279 vdd.t289 4.06363
R5973 vdd.n277 vdd.t293 4.06363
R5974 vdd.n277 vdd.t185 4.06363
R5975 vdd.n275 vdd.t216 4.06363
R5976 vdd.n275 vdd.t291 4.06363
R5977 vdd.n273 vdd.t297 4.06363
R5978 vdd.n273 vdd.t214 4.06363
R5979 vdd.n187 vdd.t242 4.06363
R5980 vdd.n187 vdd.t281 4.06363
R5981 vdd.n185 vdd.t298 4.06363
R5982 vdd.n185 vdd.t190 4.06363
R5983 vdd.n183 vdd.t199 4.06363
R5984 vdd.n183 vdd.t261 4.06363
R5985 vdd.n181 vdd.t262 4.06363
R5986 vdd.n181 vdd.t290 4.06363
R5987 vdd.n179 vdd.t156 4.06363
R5988 vdd.n179 vdd.t226 4.06363
R5989 vdd.n177 vdd.t265 4.06363
R5990 vdd.n177 vdd.t275 4.06363
R5991 vdd.n175 vdd.t283 4.06363
R5992 vdd.n175 vdd.t162 4.06363
R5993 vdd.n173 vdd.t191 4.06363
R5994 vdd.n173 vdd.t282 4.06363
R5995 vdd.n171 vdd.t286 4.06363
R5996 vdd.n171 vdd.t188 4.06363
R5997 vdd.n86 vdd.t220 4.06363
R5998 vdd.n86 vdd.t294 4.06363
R5999 vdd.n84 vdd.t196 4.06363
R6000 vdd.n84 vdd.t278 4.06363
R6001 vdd.n82 vdd.t231 4.06363
R6002 vdd.n82 vdd.t263 4.06363
R6003 vdd.n80 vdd.t211 4.06363
R6004 vdd.n80 vdd.t284 4.06363
R6005 vdd.n78 vdd.t174 4.06363
R6006 vdd.n78 vdd.t272 4.06363
R6007 vdd.n76 vdd.t169 4.06363
R6008 vdd.n76 vdd.t257 4.06363
R6009 vdd.n74 vdd.t193 4.06363
R6010 vdd.n74 vdd.t276 4.06363
R6011 vdd.n72 vdd.t164 4.06363
R6012 vdd.n72 vdd.t228 4.06363
R6013 vdd.n70 vdd.t150 4.06363
R6014 vdd.n70 vdd.t202 4.06363
R6015 vdd.n1831 vdd.t266 4.06363
R6016 vdd.n1831 vdd.t213 4.06363
R6017 vdd.n1833 vdd.t208 4.06363
R6018 vdd.n1833 vdd.t268 4.06363
R6019 vdd.n1835 vdd.t250 4.06363
R6020 vdd.n1835 vdd.t248 4.06363
R6021 vdd.n1837 vdd.t203 4.06363
R6022 vdd.n1837 vdd.t173 4.06363
R6023 vdd.n1839 vdd.t171 4.06363
R6024 vdd.n1839 vdd.t247 4.06363
R6025 vdd.n1841 vdd.t224 4.06363
R6026 vdd.n1841 vdd.t172 4.06363
R6027 vdd.n1843 vdd.t165 4.06363
R6028 vdd.n1843 vdd.t269 4.06363
R6029 vdd.n1845 vdd.t267 4.06363
R6030 vdd.n1845 vdd.t217 4.06363
R6031 vdd.n1847 vdd.t209 4.06363
R6032 vdd.n1847 vdd.t296 4.06363
R6033 vdd.n1729 vdd.t252 4.06363
R6034 vdd.n1729 vdd.t186 4.06363
R6035 vdd.n1731 vdd.t182 4.06363
R6036 vdd.n1731 vdd.t255 4.06363
R6037 vdd.n1733 vdd.t239 4.06363
R6038 vdd.n1733 vdd.t235 4.06363
R6039 vdd.n1735 vdd.t177 4.06363
R6040 vdd.n1735 vdd.t152 4.06363
R6041 vdd.n1737 vdd.t144 4.06363
R6042 vdd.n1737 vdd.t230 4.06363
R6043 vdd.n1739 vdd.t207 4.06363
R6044 vdd.n1739 vdd.t148 4.06363
R6045 vdd.n1741 vdd.t142 4.06363
R6046 vdd.n1741 vdd.t259 4.06363
R6047 vdd.n1743 vdd.t254 4.06363
R6048 vdd.n1743 vdd.t197 4.06363
R6049 vdd.n1745 vdd.t184 4.06363
R6050 vdd.n1745 vdd.t285 4.06363
R6051 vdd.n1628 vdd.t205 4.06363
R6052 vdd.n1628 vdd.t154 4.06363
R6053 vdd.n1630 vdd.t229 4.06363
R6054 vdd.n1630 vdd.t167 4.06363
R6055 vdd.n1632 vdd.t277 4.06363
R6056 vdd.n1632 vdd.t299 4.06363
R6057 vdd.n1634 vdd.t258 4.06363
R6058 vdd.n1634 vdd.t170 4.06363
R6059 vdd.n1636 vdd.t243 4.06363
R6060 vdd.n1636 vdd.t179 4.06363
R6061 vdd.n1638 vdd.t287 4.06363
R6062 vdd.n1638 vdd.t212 4.06363
R6063 vdd.n1640 vdd.t264 4.06363
R6064 vdd.n1640 vdd.t233 4.06363
R6065 vdd.n1642 vdd.t279 4.06363
R6066 vdd.n1642 vdd.t195 4.06363
R6067 vdd.n1644 vdd.t295 4.06363
R6068 vdd.n1644 vdd.t223 4.06363
R6069 vdd.n26 vdd.t136 3.9605
R6070 vdd.n26 vdd.t134 3.9605
R6071 vdd.n23 vdd.t18 3.9605
R6072 vdd.n23 vdd.t112 3.9605
R6073 vdd.n21 vdd.t115 3.9605
R6074 vdd.n21 vdd.t100 3.9605
R6075 vdd.n20 vdd.t13 3.9605
R6076 vdd.n20 vdd.t17 3.9605
R6077 vdd.n15 vdd.t301 3.9605
R6078 vdd.n15 vdd.t16 3.9605
R6079 vdd.n16 vdd.t12 3.9605
R6080 vdd.n16 vdd.t113 3.9605
R6081 vdd.n18 vdd.t116 3.9605
R6082 vdd.n18 vdd.t98 3.9605
R6083 vdd.n25 vdd.t135 3.9605
R6084 vdd.n25 vdd.t99 3.9605
R6085 vdd.n3080 vdd.n3079 3.74684
R6086 vdd.n2520 vdd.n2519 3.74684
R6087 vdd.n7 vdd.t123 3.61217
R6088 vdd.n7 vdd.t121 3.61217
R6089 vdd.n8 vdd.t102 3.61217
R6090 vdd.n8 vdd.t108 3.61217
R6091 vdd.n10 vdd.t4 3.61217
R6092 vdd.n10 vdd.t133 3.61217
R6093 vdd.n12 vdd.t126 3.61217
R6094 vdd.n12 vdd.t6 3.61217
R6095 vdd.n5 vdd.t140 3.61217
R6096 vdd.n5 vdd.t129 3.61217
R6097 vdd.n3 vdd.t119 3.61217
R6098 vdd.n3 vdd.t138 3.61217
R6099 vdd.n1 vdd.t2 3.61217
R6100 vdd.n1 vdd.t303 3.61217
R6101 vdd.n0 vdd.t110 3.61217
R6102 vdd.n0 vdd.t104 3.61217
R6103 vdd.n2497 vdd.t19 3.51482
R6104 vdd.n2552 vdd.t20 3.51482
R6105 vdd.n3047 vdd.t106 3.51482
R6106 vdd.n3102 vdd.t111 3.51482
R6107 vdd.n316 vdd.n315 3.49141
R6108 vdd.n257 vdd.n256 3.49141
R6109 vdd.n214 vdd.n213 3.49141
R6110 vdd.n155 vdd.n154 3.49141
R6111 vdd.n113 vdd.n112 3.49141
R6112 vdd.n54 vdd.n53 3.49141
R6113 vdd.n1815 vdd.n1814 3.49141
R6114 vdd.n1874 vdd.n1873 3.49141
R6115 vdd.n1713 vdd.n1712 3.49141
R6116 vdd.n1772 vdd.n1771 3.49141
R6117 vdd.n1612 vdd.n1611 3.49141
R6118 vdd.n1671 vdd.n1670 3.49141
R6119 vdd.n2572 vdd.t118 3.40145
R6120 vdd.n2726 vdd.t139 3.40145
R6121 vdd.n3010 vdd.t5 3.40145
R6122 vdd.n3029 vdd.t132 3.40145
R6123 vdd.n1956 vdd.t153 3.28809
R6124 vdd.n3429 vdd.t149 3.28809
R6125 vdd.t181 vdd.n1184 3.06136
R6126 vdd.n3454 vdd.t227 3.06136
R6127 vdd.t302 vdd.n1015 2.94799
R6128 vdd.n930 vdd.t101 2.94799
R6129 vdd.n1914 vdd.t151 2.83463
R6130 vdd.n2473 vdd.t30 2.83463
R6131 vdd.n2579 vdd.t68 2.83463
R6132 vdd.n3023 vdd.t72 2.83463
R6133 vdd.n3171 vdd.t26 2.83463
R6134 vdd.n644 vdd.t168 2.83463
R6135 vdd.n319 vdd.n298 2.71565
R6136 vdd.n260 vdd.n239 2.71565
R6137 vdd.n217 vdd.n196 2.71565
R6138 vdd.n158 vdd.n137 2.71565
R6139 vdd.n116 vdd.n95 2.71565
R6140 vdd.n57 vdd.n36 2.71565
R6141 vdd.n1818 vdd.n1797 2.71565
R6142 vdd.n1877 vdd.n1856 2.71565
R6143 vdd.n1716 vdd.n1695 2.71565
R6144 vdd.n1775 vdd.n1754 2.71565
R6145 vdd.n1615 vdd.n1594 2.71565
R6146 vdd.n1674 vdd.n1653 2.71565
R6147 vdd.t143 vdd.n1212 2.6079
R6148 vdd.n1070 vdd.t8 2.6079
R6149 vdd.n2358 vdd.t124 2.6079
R6150 vdd.n2977 vdd.t15 2.6079
R6151 vdd.t114 vdd.n874 2.6079
R6152 vdd.n3577 vdd.t225 2.6079
R6153 vdd.n306 vdd.n305 2.4129
R6154 vdd.n247 vdd.n246 2.4129
R6155 vdd.n204 vdd.n203 2.4129
R6156 vdd.n145 vdd.n144 2.4129
R6157 vdd.n103 vdd.n102 2.4129
R6158 vdd.n44 vdd.n43 2.4129
R6159 vdd.n1805 vdd.n1804 2.4129
R6160 vdd.n1864 vdd.n1863 2.4129
R6161 vdd.n1703 vdd.n1702 2.4129
R6162 vdd.n1762 vdd.n1761 2.4129
R6163 vdd.n1602 vdd.n1601 2.4129
R6164 vdd.n1661 vdd.n1660 2.4129
R6165 vdd.n1566 vdd.t232 2.38117
R6166 vdd.n1974 vdd.t48 2.38117
R6167 vdd.n3413 vdd.t22 2.38117
R6168 vdd.n3568 vdd.t198 2.38117
R6169 vdd.n2182 vdd.n1984 2.27742
R6170 vdd.n2183 vdd.n2182 2.27742
R6171 vdd.n3398 vdd.n3397 2.27742
R6172 vdd.n3399 vdd.n3398 2.27742
R6173 vdd.n3276 vdd.n3275 2.27742
R6174 vdd.n3275 vdd.n784 2.27742
R6175 vdd.n2205 vdd.n1145 2.27742
R6176 vdd.n2205 vdd.n1146 2.27742
R6177 vdd.n2358 vdd.t109 2.2678
R6178 vdd.n2977 vdd.t120 2.2678
R6179 vdd.t253 vdd.n1241 2.15444
R6180 vdd.n3559 vdd.t189 2.15444
R6181 vdd.n2546 vdd.t103 2.04107
R6182 vdd.n3053 vdd.t122 2.04107
R6183 vdd.n320 vdd.n296 1.93989
R6184 vdd.n261 vdd.n237 1.93989
R6185 vdd.n218 vdd.n194 1.93989
R6186 vdd.n159 vdd.n135 1.93989
R6187 vdd.n117 vdd.n93 1.93989
R6188 vdd.n58 vdd.n34 1.93989
R6189 vdd.n1819 vdd.n1795 1.93989
R6190 vdd.n1878 vdd.n1854 1.93989
R6191 vdd.n1717 vdd.n1693 1.93989
R6192 vdd.n1776 vdd.n1752 1.93989
R6193 vdd.n1616 vdd.n1592 1.93989
R6194 vdd.n1675 vdd.n1651 1.93989
R6195 vdd.n1524 vdd.t236 1.92771
R6196 vdd.t159 vdd.n375 1.92771
R6197 vdd.n1532 vdd.t222 1.70098
R6198 vdd.n2522 vdd.t10 1.70098
R6199 vdd.n2528 vdd.t11 1.70098
R6200 vdd.n3071 vdd.t14 1.70098
R6201 vdd.n3077 vdd.t97 1.70098
R6202 vdd.n3553 vdd.t219 1.70098
R6203 vdd.n1557 vdd.t141 1.47425
R6204 vdd.n361 vdd.t260 1.47425
R6205 vdd.n2552 vdd.t1 1.36088
R6206 vdd.n3047 vdd.t107 1.36088
R6207 vdd.n1223 vdd.t147 1.24752
R6208 vdd.t210 vdd.n3575 1.24752
R6209 vdd.n331 vdd.n291 1.16414
R6210 vdd.n324 vdd.n323 1.16414
R6211 vdd.n272 vdd.n232 1.16414
R6212 vdd.n265 vdd.n264 1.16414
R6213 vdd.n229 vdd.n189 1.16414
R6214 vdd.n222 vdd.n221 1.16414
R6215 vdd.n170 vdd.n130 1.16414
R6216 vdd.n163 vdd.n162 1.16414
R6217 vdd.n128 vdd.n88 1.16414
R6218 vdd.n121 vdd.n120 1.16414
R6219 vdd.n69 vdd.n29 1.16414
R6220 vdd.n62 vdd.n61 1.16414
R6221 vdd.n1830 vdd.n1790 1.16414
R6222 vdd.n1823 vdd.n1822 1.16414
R6223 vdd.n1889 vdd.n1849 1.16414
R6224 vdd.n1882 vdd.n1881 1.16414
R6225 vdd.n1728 vdd.n1688 1.16414
R6226 vdd.n1721 vdd.n1720 1.16414
R6227 vdd.n1787 vdd.n1747 1.16414
R6228 vdd.n1780 vdd.n1779 1.16414
R6229 vdd.n1627 vdd.n1587 1.16414
R6230 vdd.n1620 vdd.n1619 1.16414
R6231 vdd.n1686 vdd.n1646 1.16414
R6232 vdd.n1679 vdd.n1678 1.16414
R6233 vdd.n1892 vdd.n28 1.11236
R6234 vdd vdd.n3582 1.10453
R6235 vdd.n1906 vdd.t176 1.02079
R6236 vdd.t82 vdd.t10 1.02079
R6237 vdd.t97 vdd.t41 1.02079
R6238 vdd.t256 vdd.n633 1.02079
R6239 vdd.n1403 vdd.n1399 0.970197
R6240 vdd.n2203 vdd.n2202 0.970197
R6241 vdd.n618 vdd.n428 0.970197
R6242 vdd.n3277 vdd.n690 0.970197
R6243 vdd.t137 vdd.n992 0.907421
R6244 vdd.n946 vdd.t3 0.907421
R6245 vdd.n1922 vdd.t234 0.794056
R6246 vdd.t130 vdd.n1067 0.794056
R6247 vdd.n1039 vdd.t105 0.794056
R6248 vdd.t127 vdd.n905 0.794056
R6249 vdd.n877 vdd.t7 0.794056
R6250 vdd.n3463 vdd.t192 0.794056
R6251 vdd.n1947 vdd.t204 0.567326
R6252 vdd.t187 vdd.n662 0.567326
R6253 vdd.n2193 vdd.n2192 0.530988
R6254 vdd.n726 vdd.n682 0.530988
R6255 vdd.n464 vdd.n391 0.530988
R6256 vdd.n3532 vdd.n3531 0.530988
R6257 vdd.n3409 vdd.n3408 0.530988
R6258 vdd.n1969 vdd.n1147 0.530988
R6259 vdd.n1401 vdd.n1266 0.530988
R6260 vdd.n1503 vdd.n1502 0.530988
R6261 vdd.n4 vdd.n2 0.459552
R6262 vdd.n11 vdd.n9 0.459552
R6263 vdd.n329 vdd.n328 0.388379
R6264 vdd.n295 vdd.n293 0.388379
R6265 vdd.n270 vdd.n269 0.388379
R6266 vdd.n236 vdd.n234 0.388379
R6267 vdd.n227 vdd.n226 0.388379
R6268 vdd.n193 vdd.n191 0.388379
R6269 vdd.n168 vdd.n167 0.388379
R6270 vdd.n134 vdd.n132 0.388379
R6271 vdd.n126 vdd.n125 0.388379
R6272 vdd.n92 vdd.n90 0.388379
R6273 vdd.n67 vdd.n66 0.388379
R6274 vdd.n33 vdd.n31 0.388379
R6275 vdd.n1828 vdd.n1827 0.388379
R6276 vdd.n1794 vdd.n1792 0.388379
R6277 vdd.n1887 vdd.n1886 0.388379
R6278 vdd.n1853 vdd.n1851 0.388379
R6279 vdd.n1726 vdd.n1725 0.388379
R6280 vdd.n1692 vdd.n1690 0.388379
R6281 vdd.n1785 vdd.n1784 0.388379
R6282 vdd.n1751 vdd.n1749 0.388379
R6283 vdd.n1625 vdd.n1624 0.388379
R6284 vdd.n1591 vdd.n1589 0.388379
R6285 vdd.n1684 vdd.n1683 0.388379
R6286 vdd.n1650 vdd.n1648 0.388379
R6287 vdd.n19 vdd.n17 0.387128
R6288 vdd.n24 vdd.n22 0.387128
R6289 vdd.n6 vdd.n4 0.358259
R6290 vdd.n13 vdd.n11 0.358259
R6291 vdd.n276 vdd.n274 0.358259
R6292 vdd.n278 vdd.n276 0.358259
R6293 vdd.n280 vdd.n278 0.358259
R6294 vdd.n282 vdd.n280 0.358259
R6295 vdd.n284 vdd.n282 0.358259
R6296 vdd.n286 vdd.n284 0.358259
R6297 vdd.n288 vdd.n286 0.358259
R6298 vdd.n290 vdd.n288 0.358259
R6299 vdd.n332 vdd.n290 0.358259
R6300 vdd.n174 vdd.n172 0.358259
R6301 vdd.n176 vdd.n174 0.358259
R6302 vdd.n178 vdd.n176 0.358259
R6303 vdd.n180 vdd.n178 0.358259
R6304 vdd.n182 vdd.n180 0.358259
R6305 vdd.n184 vdd.n182 0.358259
R6306 vdd.n186 vdd.n184 0.358259
R6307 vdd.n188 vdd.n186 0.358259
R6308 vdd.n230 vdd.n188 0.358259
R6309 vdd.n73 vdd.n71 0.358259
R6310 vdd.n75 vdd.n73 0.358259
R6311 vdd.n77 vdd.n75 0.358259
R6312 vdd.n79 vdd.n77 0.358259
R6313 vdd.n81 vdd.n79 0.358259
R6314 vdd.n83 vdd.n81 0.358259
R6315 vdd.n85 vdd.n83 0.358259
R6316 vdd.n87 vdd.n85 0.358259
R6317 vdd.n129 vdd.n87 0.358259
R6318 vdd.n1890 vdd.n1848 0.358259
R6319 vdd.n1848 vdd.n1846 0.358259
R6320 vdd.n1846 vdd.n1844 0.358259
R6321 vdd.n1844 vdd.n1842 0.358259
R6322 vdd.n1842 vdd.n1840 0.358259
R6323 vdd.n1840 vdd.n1838 0.358259
R6324 vdd.n1838 vdd.n1836 0.358259
R6325 vdd.n1836 vdd.n1834 0.358259
R6326 vdd.n1834 vdd.n1832 0.358259
R6327 vdd.n1788 vdd.n1746 0.358259
R6328 vdd.n1746 vdd.n1744 0.358259
R6329 vdd.n1744 vdd.n1742 0.358259
R6330 vdd.n1742 vdd.n1740 0.358259
R6331 vdd.n1740 vdd.n1738 0.358259
R6332 vdd.n1738 vdd.n1736 0.358259
R6333 vdd.n1736 vdd.n1734 0.358259
R6334 vdd.n1734 vdd.n1732 0.358259
R6335 vdd.n1732 vdd.n1730 0.358259
R6336 vdd.n1687 vdd.n1645 0.358259
R6337 vdd.n1645 vdd.n1643 0.358259
R6338 vdd.n1643 vdd.n1641 0.358259
R6339 vdd.n1641 vdd.n1639 0.358259
R6340 vdd.n1639 vdd.n1637 0.358259
R6341 vdd.n1637 vdd.n1635 0.358259
R6342 vdd.n1635 vdd.n1633 0.358259
R6343 vdd.n1633 vdd.n1631 0.358259
R6344 vdd.n1631 vdd.n1629 0.358259
R6345 vdd.n14 vdd.n6 0.334552
R6346 vdd.n14 vdd.n13 0.334552
R6347 vdd.n27 vdd.n19 0.21707
R6348 vdd.n27 vdd.n24 0.21707
R6349 vdd.n330 vdd.n292 0.155672
R6350 vdd.n322 vdd.n292 0.155672
R6351 vdd.n322 vdd.n321 0.155672
R6352 vdd.n321 vdd.n297 0.155672
R6353 vdd.n314 vdd.n297 0.155672
R6354 vdd.n314 vdd.n313 0.155672
R6355 vdd.n313 vdd.n301 0.155672
R6356 vdd.n306 vdd.n301 0.155672
R6357 vdd.n271 vdd.n233 0.155672
R6358 vdd.n263 vdd.n233 0.155672
R6359 vdd.n263 vdd.n262 0.155672
R6360 vdd.n262 vdd.n238 0.155672
R6361 vdd.n255 vdd.n238 0.155672
R6362 vdd.n255 vdd.n254 0.155672
R6363 vdd.n254 vdd.n242 0.155672
R6364 vdd.n247 vdd.n242 0.155672
R6365 vdd.n228 vdd.n190 0.155672
R6366 vdd.n220 vdd.n190 0.155672
R6367 vdd.n220 vdd.n219 0.155672
R6368 vdd.n219 vdd.n195 0.155672
R6369 vdd.n212 vdd.n195 0.155672
R6370 vdd.n212 vdd.n211 0.155672
R6371 vdd.n211 vdd.n199 0.155672
R6372 vdd.n204 vdd.n199 0.155672
R6373 vdd.n169 vdd.n131 0.155672
R6374 vdd.n161 vdd.n131 0.155672
R6375 vdd.n161 vdd.n160 0.155672
R6376 vdd.n160 vdd.n136 0.155672
R6377 vdd.n153 vdd.n136 0.155672
R6378 vdd.n153 vdd.n152 0.155672
R6379 vdd.n152 vdd.n140 0.155672
R6380 vdd.n145 vdd.n140 0.155672
R6381 vdd.n127 vdd.n89 0.155672
R6382 vdd.n119 vdd.n89 0.155672
R6383 vdd.n119 vdd.n118 0.155672
R6384 vdd.n118 vdd.n94 0.155672
R6385 vdd.n111 vdd.n94 0.155672
R6386 vdd.n111 vdd.n110 0.155672
R6387 vdd.n110 vdd.n98 0.155672
R6388 vdd.n103 vdd.n98 0.155672
R6389 vdd.n68 vdd.n30 0.155672
R6390 vdd.n60 vdd.n30 0.155672
R6391 vdd.n60 vdd.n59 0.155672
R6392 vdd.n59 vdd.n35 0.155672
R6393 vdd.n52 vdd.n35 0.155672
R6394 vdd.n52 vdd.n51 0.155672
R6395 vdd.n51 vdd.n39 0.155672
R6396 vdd.n44 vdd.n39 0.155672
R6397 vdd.n1829 vdd.n1791 0.155672
R6398 vdd.n1821 vdd.n1791 0.155672
R6399 vdd.n1821 vdd.n1820 0.155672
R6400 vdd.n1820 vdd.n1796 0.155672
R6401 vdd.n1813 vdd.n1796 0.155672
R6402 vdd.n1813 vdd.n1812 0.155672
R6403 vdd.n1812 vdd.n1800 0.155672
R6404 vdd.n1805 vdd.n1800 0.155672
R6405 vdd.n1888 vdd.n1850 0.155672
R6406 vdd.n1880 vdd.n1850 0.155672
R6407 vdd.n1880 vdd.n1879 0.155672
R6408 vdd.n1879 vdd.n1855 0.155672
R6409 vdd.n1872 vdd.n1855 0.155672
R6410 vdd.n1872 vdd.n1871 0.155672
R6411 vdd.n1871 vdd.n1859 0.155672
R6412 vdd.n1864 vdd.n1859 0.155672
R6413 vdd.n1727 vdd.n1689 0.155672
R6414 vdd.n1719 vdd.n1689 0.155672
R6415 vdd.n1719 vdd.n1718 0.155672
R6416 vdd.n1718 vdd.n1694 0.155672
R6417 vdd.n1711 vdd.n1694 0.155672
R6418 vdd.n1711 vdd.n1710 0.155672
R6419 vdd.n1710 vdd.n1698 0.155672
R6420 vdd.n1703 vdd.n1698 0.155672
R6421 vdd.n1786 vdd.n1748 0.155672
R6422 vdd.n1778 vdd.n1748 0.155672
R6423 vdd.n1778 vdd.n1777 0.155672
R6424 vdd.n1777 vdd.n1753 0.155672
R6425 vdd.n1770 vdd.n1753 0.155672
R6426 vdd.n1770 vdd.n1769 0.155672
R6427 vdd.n1769 vdd.n1757 0.155672
R6428 vdd.n1762 vdd.n1757 0.155672
R6429 vdd.n1626 vdd.n1588 0.155672
R6430 vdd.n1618 vdd.n1588 0.155672
R6431 vdd.n1618 vdd.n1617 0.155672
R6432 vdd.n1617 vdd.n1593 0.155672
R6433 vdd.n1610 vdd.n1593 0.155672
R6434 vdd.n1610 vdd.n1609 0.155672
R6435 vdd.n1609 vdd.n1597 0.155672
R6436 vdd.n1602 vdd.n1597 0.155672
R6437 vdd.n1685 vdd.n1647 0.155672
R6438 vdd.n1677 vdd.n1647 0.155672
R6439 vdd.n1677 vdd.n1676 0.155672
R6440 vdd.n1676 vdd.n1652 0.155672
R6441 vdd.n1669 vdd.n1652 0.155672
R6442 vdd.n1669 vdd.n1668 0.155672
R6443 vdd.n1668 vdd.n1656 0.155672
R6444 vdd.n1661 vdd.n1656 0.155672
R6445 vdd.n2181 vdd.n1986 0.152939
R6446 vdd.n1992 vdd.n1986 0.152939
R6447 vdd.n1993 vdd.n1992 0.152939
R6448 vdd.n1994 vdd.n1993 0.152939
R6449 vdd.n1995 vdd.n1994 0.152939
R6450 vdd.n1999 vdd.n1995 0.152939
R6451 vdd.n2000 vdd.n1999 0.152939
R6452 vdd.n2001 vdd.n2000 0.152939
R6453 vdd.n2002 vdd.n2001 0.152939
R6454 vdd.n2006 vdd.n2002 0.152939
R6455 vdd.n2007 vdd.n2006 0.152939
R6456 vdd.n2008 vdd.n2007 0.152939
R6457 vdd.n2156 vdd.n2008 0.152939
R6458 vdd.n2156 vdd.n2155 0.152939
R6459 vdd.n2155 vdd.n2154 0.152939
R6460 vdd.n2154 vdd.n2014 0.152939
R6461 vdd.n2019 vdd.n2014 0.152939
R6462 vdd.n2020 vdd.n2019 0.152939
R6463 vdd.n2021 vdd.n2020 0.152939
R6464 vdd.n2025 vdd.n2021 0.152939
R6465 vdd.n2026 vdd.n2025 0.152939
R6466 vdd.n2027 vdd.n2026 0.152939
R6467 vdd.n2028 vdd.n2027 0.152939
R6468 vdd.n2032 vdd.n2028 0.152939
R6469 vdd.n2033 vdd.n2032 0.152939
R6470 vdd.n2034 vdd.n2033 0.152939
R6471 vdd.n2035 vdd.n2034 0.152939
R6472 vdd.n2039 vdd.n2035 0.152939
R6473 vdd.n2040 vdd.n2039 0.152939
R6474 vdd.n2041 vdd.n2040 0.152939
R6475 vdd.n2042 vdd.n2041 0.152939
R6476 vdd.n2046 vdd.n2042 0.152939
R6477 vdd.n2047 vdd.n2046 0.152939
R6478 vdd.n2048 vdd.n2047 0.152939
R6479 vdd.n2117 vdd.n2048 0.152939
R6480 vdd.n2117 vdd.n2116 0.152939
R6481 vdd.n2116 vdd.n2115 0.152939
R6482 vdd.n2115 vdd.n2054 0.152939
R6483 vdd.n2059 vdd.n2054 0.152939
R6484 vdd.n2060 vdd.n2059 0.152939
R6485 vdd.n2061 vdd.n2060 0.152939
R6486 vdd.n2065 vdd.n2061 0.152939
R6487 vdd.n2066 vdd.n2065 0.152939
R6488 vdd.n2067 vdd.n2066 0.152939
R6489 vdd.n2068 vdd.n2067 0.152939
R6490 vdd.n2072 vdd.n2068 0.152939
R6491 vdd.n2073 vdd.n2072 0.152939
R6492 vdd.n2074 vdd.n2073 0.152939
R6493 vdd.n2075 vdd.n2074 0.152939
R6494 vdd.n2076 vdd.n2075 0.152939
R6495 vdd.n2076 vdd.n1144 0.152939
R6496 vdd.n2192 vdd.n1980 0.152939
R6497 vdd.n1894 vdd.n1203 0.152939
R6498 vdd.n1909 vdd.n1203 0.152939
R6499 vdd.n1910 vdd.n1909 0.152939
R6500 vdd.n1911 vdd.n1910 0.152939
R6501 vdd.n1911 vdd.n1192 0.152939
R6502 vdd.n1926 vdd.n1192 0.152939
R6503 vdd.n1927 vdd.n1926 0.152939
R6504 vdd.n1928 vdd.n1927 0.152939
R6505 vdd.n1928 vdd.n1181 0.152939
R6506 vdd.n1942 vdd.n1181 0.152939
R6507 vdd.n1943 vdd.n1942 0.152939
R6508 vdd.n1944 vdd.n1943 0.152939
R6509 vdd.n1944 vdd.n1169 0.152939
R6510 vdd.n1959 vdd.n1169 0.152939
R6511 vdd.n1960 vdd.n1959 0.152939
R6512 vdd.n1961 vdd.n1960 0.152939
R6513 vdd.n1961 vdd.n1157 0.152939
R6514 vdd.n1978 vdd.n1157 0.152939
R6515 vdd.n1979 vdd.n1978 0.152939
R6516 vdd.n2193 vdd.n1979 0.152939
R6517 vdd.n735 vdd.n730 0.152939
R6518 vdd.n736 vdd.n735 0.152939
R6519 vdd.n737 vdd.n736 0.152939
R6520 vdd.n738 vdd.n737 0.152939
R6521 vdd.n739 vdd.n738 0.152939
R6522 vdd.n740 vdd.n739 0.152939
R6523 vdd.n741 vdd.n740 0.152939
R6524 vdd.n742 vdd.n741 0.152939
R6525 vdd.n743 vdd.n742 0.152939
R6526 vdd.n744 vdd.n743 0.152939
R6527 vdd.n745 vdd.n744 0.152939
R6528 vdd.n746 vdd.n745 0.152939
R6529 vdd.n3365 vdd.n746 0.152939
R6530 vdd.n3365 vdd.n3364 0.152939
R6531 vdd.n3364 vdd.n3363 0.152939
R6532 vdd.n3363 vdd.n748 0.152939
R6533 vdd.n749 vdd.n748 0.152939
R6534 vdd.n750 vdd.n749 0.152939
R6535 vdd.n751 vdd.n750 0.152939
R6536 vdd.n752 vdd.n751 0.152939
R6537 vdd.n753 vdd.n752 0.152939
R6538 vdd.n754 vdd.n753 0.152939
R6539 vdd.n755 vdd.n754 0.152939
R6540 vdd.n756 vdd.n755 0.152939
R6541 vdd.n757 vdd.n756 0.152939
R6542 vdd.n758 vdd.n757 0.152939
R6543 vdd.n759 vdd.n758 0.152939
R6544 vdd.n760 vdd.n759 0.152939
R6545 vdd.n761 vdd.n760 0.152939
R6546 vdd.n762 vdd.n761 0.152939
R6547 vdd.n763 vdd.n762 0.152939
R6548 vdd.n764 vdd.n763 0.152939
R6549 vdd.n765 vdd.n764 0.152939
R6550 vdd.n766 vdd.n765 0.152939
R6551 vdd.n3319 vdd.n766 0.152939
R6552 vdd.n3319 vdd.n3318 0.152939
R6553 vdd.n3318 vdd.n3317 0.152939
R6554 vdd.n3317 vdd.n770 0.152939
R6555 vdd.n771 vdd.n770 0.152939
R6556 vdd.n772 vdd.n771 0.152939
R6557 vdd.n773 vdd.n772 0.152939
R6558 vdd.n774 vdd.n773 0.152939
R6559 vdd.n775 vdd.n774 0.152939
R6560 vdd.n776 vdd.n775 0.152939
R6561 vdd.n777 vdd.n776 0.152939
R6562 vdd.n778 vdd.n777 0.152939
R6563 vdd.n779 vdd.n778 0.152939
R6564 vdd.n780 vdd.n779 0.152939
R6565 vdd.n781 vdd.n780 0.152939
R6566 vdd.n782 vdd.n781 0.152939
R6567 vdd.n783 vdd.n782 0.152939
R6568 vdd.n727 vdd.n726 0.152939
R6569 vdd.n3416 vdd.n682 0.152939
R6570 vdd.n3417 vdd.n3416 0.152939
R6571 vdd.n3418 vdd.n3417 0.152939
R6572 vdd.n3418 vdd.n670 0.152939
R6573 vdd.n3433 vdd.n670 0.152939
R6574 vdd.n3434 vdd.n3433 0.152939
R6575 vdd.n3435 vdd.n3434 0.152939
R6576 vdd.n3435 vdd.n659 0.152939
R6577 vdd.n3449 vdd.n659 0.152939
R6578 vdd.n3450 vdd.n3449 0.152939
R6579 vdd.n3451 vdd.n3450 0.152939
R6580 vdd.n3451 vdd.n647 0.152939
R6581 vdd.n3466 vdd.n647 0.152939
R6582 vdd.n3467 vdd.n3466 0.152939
R6583 vdd.n3468 vdd.n3467 0.152939
R6584 vdd.n3468 vdd.n636 0.152939
R6585 vdd.n3485 vdd.n636 0.152939
R6586 vdd.n3486 vdd.n3485 0.152939
R6587 vdd.n3487 vdd.n3486 0.152939
R6588 vdd.n3487 vdd.n334 0.152939
R6589 vdd.n3580 vdd.n335 0.152939
R6590 vdd.n346 vdd.n335 0.152939
R6591 vdd.n347 vdd.n346 0.152939
R6592 vdd.n348 vdd.n347 0.152939
R6593 vdd.n355 vdd.n348 0.152939
R6594 vdd.n356 vdd.n355 0.152939
R6595 vdd.n357 vdd.n356 0.152939
R6596 vdd.n358 vdd.n357 0.152939
R6597 vdd.n366 vdd.n358 0.152939
R6598 vdd.n367 vdd.n366 0.152939
R6599 vdd.n368 vdd.n367 0.152939
R6600 vdd.n369 vdd.n368 0.152939
R6601 vdd.n377 vdd.n369 0.152939
R6602 vdd.n378 vdd.n377 0.152939
R6603 vdd.n379 vdd.n378 0.152939
R6604 vdd.n380 vdd.n379 0.152939
R6605 vdd.n388 vdd.n380 0.152939
R6606 vdd.n389 vdd.n388 0.152939
R6607 vdd.n390 vdd.n389 0.152939
R6608 vdd.n391 vdd.n390 0.152939
R6609 vdd.n464 vdd.n463 0.152939
R6610 vdd.n470 vdd.n463 0.152939
R6611 vdd.n471 vdd.n470 0.152939
R6612 vdd.n472 vdd.n471 0.152939
R6613 vdd.n472 vdd.n461 0.152939
R6614 vdd.n480 vdd.n461 0.152939
R6615 vdd.n481 vdd.n480 0.152939
R6616 vdd.n482 vdd.n481 0.152939
R6617 vdd.n482 vdd.n459 0.152939
R6618 vdd.n490 vdd.n459 0.152939
R6619 vdd.n491 vdd.n490 0.152939
R6620 vdd.n492 vdd.n491 0.152939
R6621 vdd.n492 vdd.n457 0.152939
R6622 vdd.n500 vdd.n457 0.152939
R6623 vdd.n501 vdd.n500 0.152939
R6624 vdd.n502 vdd.n501 0.152939
R6625 vdd.n502 vdd.n455 0.152939
R6626 vdd.n510 vdd.n455 0.152939
R6627 vdd.n511 vdd.n510 0.152939
R6628 vdd.n512 vdd.n511 0.152939
R6629 vdd.n512 vdd.n451 0.152939
R6630 vdd.n520 vdd.n451 0.152939
R6631 vdd.n521 vdd.n520 0.152939
R6632 vdd.n522 vdd.n521 0.152939
R6633 vdd.n522 vdd.n449 0.152939
R6634 vdd.n530 vdd.n449 0.152939
R6635 vdd.n531 vdd.n530 0.152939
R6636 vdd.n532 vdd.n531 0.152939
R6637 vdd.n532 vdd.n447 0.152939
R6638 vdd.n540 vdd.n447 0.152939
R6639 vdd.n541 vdd.n540 0.152939
R6640 vdd.n542 vdd.n541 0.152939
R6641 vdd.n542 vdd.n445 0.152939
R6642 vdd.n550 vdd.n445 0.152939
R6643 vdd.n551 vdd.n550 0.152939
R6644 vdd.n552 vdd.n551 0.152939
R6645 vdd.n552 vdd.n443 0.152939
R6646 vdd.n560 vdd.n443 0.152939
R6647 vdd.n561 vdd.n560 0.152939
R6648 vdd.n562 vdd.n561 0.152939
R6649 vdd.n562 vdd.n439 0.152939
R6650 vdd.n570 vdd.n439 0.152939
R6651 vdd.n571 vdd.n570 0.152939
R6652 vdd.n572 vdd.n571 0.152939
R6653 vdd.n572 vdd.n437 0.152939
R6654 vdd.n580 vdd.n437 0.152939
R6655 vdd.n581 vdd.n580 0.152939
R6656 vdd.n582 vdd.n581 0.152939
R6657 vdd.n582 vdd.n435 0.152939
R6658 vdd.n590 vdd.n435 0.152939
R6659 vdd.n591 vdd.n590 0.152939
R6660 vdd.n592 vdd.n591 0.152939
R6661 vdd.n592 vdd.n433 0.152939
R6662 vdd.n600 vdd.n433 0.152939
R6663 vdd.n601 vdd.n600 0.152939
R6664 vdd.n602 vdd.n601 0.152939
R6665 vdd.n602 vdd.n431 0.152939
R6666 vdd.n610 vdd.n431 0.152939
R6667 vdd.n611 vdd.n610 0.152939
R6668 vdd.n612 vdd.n611 0.152939
R6669 vdd.n612 vdd.n429 0.152939
R6670 vdd.n619 vdd.n429 0.152939
R6671 vdd.n3532 vdd.n619 0.152939
R6672 vdd.n3410 vdd.n3409 0.152939
R6673 vdd.n3410 vdd.n675 0.152939
R6674 vdd.n3424 vdd.n675 0.152939
R6675 vdd.n3425 vdd.n3424 0.152939
R6676 vdd.n3426 vdd.n3425 0.152939
R6677 vdd.n3426 vdd.n665 0.152939
R6678 vdd.n3441 vdd.n665 0.152939
R6679 vdd.n3442 vdd.n3441 0.152939
R6680 vdd.n3443 vdd.n3442 0.152939
R6681 vdd.n3443 vdd.n652 0.152939
R6682 vdd.n3457 vdd.n652 0.152939
R6683 vdd.n3458 vdd.n3457 0.152939
R6684 vdd.n3459 vdd.n3458 0.152939
R6685 vdd.n3459 vdd.n641 0.152939
R6686 vdd.n3474 vdd.n641 0.152939
R6687 vdd.n3475 vdd.n3474 0.152939
R6688 vdd.n3476 vdd.n3475 0.152939
R6689 vdd.n3478 vdd.n3476 0.152939
R6690 vdd.n3478 vdd.n3477 0.152939
R6691 vdd.n3477 vdd.n630 0.152939
R6692 vdd.n3495 vdd.n630 0.152939
R6693 vdd.n3496 vdd.n3495 0.152939
R6694 vdd.n3497 vdd.n3496 0.152939
R6695 vdd.n3497 vdd.n628 0.152939
R6696 vdd.n3502 vdd.n628 0.152939
R6697 vdd.n3503 vdd.n3502 0.152939
R6698 vdd.n3504 vdd.n3503 0.152939
R6699 vdd.n3504 vdd.n626 0.152939
R6700 vdd.n3509 vdd.n626 0.152939
R6701 vdd.n3510 vdd.n3509 0.152939
R6702 vdd.n3511 vdd.n3510 0.152939
R6703 vdd.n3511 vdd.n624 0.152939
R6704 vdd.n3517 vdd.n624 0.152939
R6705 vdd.n3518 vdd.n3517 0.152939
R6706 vdd.n3519 vdd.n3518 0.152939
R6707 vdd.n3519 vdd.n622 0.152939
R6708 vdd.n3524 vdd.n622 0.152939
R6709 vdd.n3525 vdd.n3524 0.152939
R6710 vdd.n3526 vdd.n3525 0.152939
R6711 vdd.n3526 vdd.n620 0.152939
R6712 vdd.n3531 vdd.n620 0.152939
R6713 vdd.n3408 vdd.n687 0.152939
R6714 vdd.n2204 vdd.n1147 0.152939
R6715 vdd.n1510 vdd.n1266 0.152939
R6716 vdd.n1511 vdd.n1510 0.152939
R6717 vdd.n1512 vdd.n1511 0.152939
R6718 vdd.n1512 vdd.n1254 0.152939
R6719 vdd.n1527 vdd.n1254 0.152939
R6720 vdd.n1528 vdd.n1527 0.152939
R6721 vdd.n1529 vdd.n1528 0.152939
R6722 vdd.n1529 vdd.n1244 0.152939
R6723 vdd.n1544 vdd.n1244 0.152939
R6724 vdd.n1545 vdd.n1544 0.152939
R6725 vdd.n1546 vdd.n1545 0.152939
R6726 vdd.n1546 vdd.n1231 0.152939
R6727 vdd.n1560 vdd.n1231 0.152939
R6728 vdd.n1561 vdd.n1560 0.152939
R6729 vdd.n1562 vdd.n1561 0.152939
R6730 vdd.n1562 vdd.n1220 0.152939
R6731 vdd.n1577 vdd.n1220 0.152939
R6732 vdd.n1578 vdd.n1577 0.152939
R6733 vdd.n1579 vdd.n1578 0.152939
R6734 vdd.n1579 vdd.n1209 0.152939
R6735 vdd.n1900 vdd.n1209 0.152939
R6736 vdd.n1901 vdd.n1900 0.152939
R6737 vdd.n1902 vdd.n1901 0.152939
R6738 vdd.n1902 vdd.n1197 0.152939
R6739 vdd.n1917 vdd.n1197 0.152939
R6740 vdd.n1918 vdd.n1917 0.152939
R6741 vdd.n1919 vdd.n1918 0.152939
R6742 vdd.n1919 vdd.n1187 0.152939
R6743 vdd.n1934 vdd.n1187 0.152939
R6744 vdd.n1935 vdd.n1934 0.152939
R6745 vdd.n1936 vdd.n1935 0.152939
R6746 vdd.n1936 vdd.n1174 0.152939
R6747 vdd.n1950 vdd.n1174 0.152939
R6748 vdd.n1951 vdd.n1950 0.152939
R6749 vdd.n1952 vdd.n1951 0.152939
R6750 vdd.n1952 vdd.n1164 0.152939
R6751 vdd.n1967 vdd.n1164 0.152939
R6752 vdd.n1968 vdd.n1967 0.152939
R6753 vdd.n1971 vdd.n1968 0.152939
R6754 vdd.n1971 vdd.n1970 0.152939
R6755 vdd.n1970 vdd.n1969 0.152939
R6756 vdd.n1502 vdd.n1271 0.152939
R6757 vdd.n1495 vdd.n1271 0.152939
R6758 vdd.n1495 vdd.n1494 0.152939
R6759 vdd.n1494 vdd.n1493 0.152939
R6760 vdd.n1493 vdd.n1308 0.152939
R6761 vdd.n1489 vdd.n1308 0.152939
R6762 vdd.n1489 vdd.n1488 0.152939
R6763 vdd.n1488 vdd.n1487 0.152939
R6764 vdd.n1487 vdd.n1314 0.152939
R6765 vdd.n1483 vdd.n1314 0.152939
R6766 vdd.n1483 vdd.n1482 0.152939
R6767 vdd.n1482 vdd.n1481 0.152939
R6768 vdd.n1481 vdd.n1320 0.152939
R6769 vdd.n1477 vdd.n1320 0.152939
R6770 vdd.n1477 vdd.n1476 0.152939
R6771 vdd.n1476 vdd.n1475 0.152939
R6772 vdd.n1475 vdd.n1326 0.152939
R6773 vdd.n1471 vdd.n1326 0.152939
R6774 vdd.n1471 vdd.n1470 0.152939
R6775 vdd.n1470 vdd.n1469 0.152939
R6776 vdd.n1469 vdd.n1334 0.152939
R6777 vdd.n1465 vdd.n1334 0.152939
R6778 vdd.n1465 vdd.n1464 0.152939
R6779 vdd.n1464 vdd.n1463 0.152939
R6780 vdd.n1463 vdd.n1340 0.152939
R6781 vdd.n1459 vdd.n1340 0.152939
R6782 vdd.n1459 vdd.n1458 0.152939
R6783 vdd.n1458 vdd.n1457 0.152939
R6784 vdd.n1457 vdd.n1346 0.152939
R6785 vdd.n1453 vdd.n1346 0.152939
R6786 vdd.n1453 vdd.n1452 0.152939
R6787 vdd.n1452 vdd.n1451 0.152939
R6788 vdd.n1451 vdd.n1352 0.152939
R6789 vdd.n1447 vdd.n1352 0.152939
R6790 vdd.n1447 vdd.n1446 0.152939
R6791 vdd.n1446 vdd.n1445 0.152939
R6792 vdd.n1445 vdd.n1358 0.152939
R6793 vdd.n1441 vdd.n1358 0.152939
R6794 vdd.n1441 vdd.n1440 0.152939
R6795 vdd.n1440 vdd.n1439 0.152939
R6796 vdd.n1439 vdd.n1364 0.152939
R6797 vdd.n1432 vdd.n1364 0.152939
R6798 vdd.n1432 vdd.n1431 0.152939
R6799 vdd.n1431 vdd.n1430 0.152939
R6800 vdd.n1430 vdd.n1369 0.152939
R6801 vdd.n1426 vdd.n1369 0.152939
R6802 vdd.n1426 vdd.n1425 0.152939
R6803 vdd.n1425 vdd.n1424 0.152939
R6804 vdd.n1424 vdd.n1375 0.152939
R6805 vdd.n1420 vdd.n1375 0.152939
R6806 vdd.n1420 vdd.n1419 0.152939
R6807 vdd.n1419 vdd.n1418 0.152939
R6808 vdd.n1418 vdd.n1381 0.152939
R6809 vdd.n1414 vdd.n1381 0.152939
R6810 vdd.n1414 vdd.n1413 0.152939
R6811 vdd.n1413 vdd.n1412 0.152939
R6812 vdd.n1412 vdd.n1387 0.152939
R6813 vdd.n1408 vdd.n1387 0.152939
R6814 vdd.n1408 vdd.n1407 0.152939
R6815 vdd.n1407 vdd.n1406 0.152939
R6816 vdd.n1406 vdd.n1393 0.152939
R6817 vdd.n1402 vdd.n1393 0.152939
R6818 vdd.n1402 vdd.n1401 0.152939
R6819 vdd.n1504 vdd.n1503 0.152939
R6820 vdd.n1504 vdd.n1260 0.152939
R6821 vdd.n1519 vdd.n1260 0.152939
R6822 vdd.n1520 vdd.n1519 0.152939
R6823 vdd.n1521 vdd.n1520 0.152939
R6824 vdd.n1521 vdd.n1249 0.152939
R6825 vdd.n1536 vdd.n1249 0.152939
R6826 vdd.n1537 vdd.n1536 0.152939
R6827 vdd.n1538 vdd.n1537 0.152939
R6828 vdd.n1538 vdd.n1238 0.152939
R6829 vdd.n1552 vdd.n1238 0.152939
R6830 vdd.n1553 vdd.n1552 0.152939
R6831 vdd.n1554 vdd.n1553 0.152939
R6832 vdd.n1554 vdd.n1226 0.152939
R6833 vdd.n1569 vdd.n1226 0.152939
R6834 vdd.n1570 vdd.n1569 0.152939
R6835 vdd.n1571 vdd.n1570 0.152939
R6836 vdd.n1571 vdd.n1215 0.152939
R6837 vdd.n1585 vdd.n1215 0.152939
R6838 vdd.n1586 vdd.n1585 0.152939
R6839 vdd.n1507 vdd.t64 0.113865
R6840 vdd.n2491 vdd.t117 0.113865
R6841 vdd.n2558 vdd.t131 0.113865
R6842 vdd.n3041 vdd.t0 0.113865
R6843 vdd.n3108 vdd.t9 0.113865
R6844 vdd.t34 vdd.n386 0.113865
R6845 vdd.n2182 vdd.n1980 0.110256
R6846 vdd.n3398 vdd.n727 0.110256
R6847 vdd.n3275 vdd.n687 0.110256
R6848 vdd.n2205 vdd.n2204 0.110256
R6849 vdd.n1894 vdd.n1893 0.0695946
R6850 vdd.n3581 vdd.n334 0.0695946
R6851 vdd.n3581 vdd.n3580 0.0695946
R6852 vdd.n1893 vdd.n1586 0.0695946
R6853 vdd.n2182 vdd.n2181 0.0431829
R6854 vdd.n2205 vdd.n1144 0.0431829
R6855 vdd.n3398 vdd.n730 0.0431829
R6856 vdd.n3275 vdd.n783 0.0431829
R6857 vdd vdd.n28 0.00833333
R6858 CSoutput.n19 CSoutput.t188 184.661
R6859 CSoutput.n78 CSoutput.n77 165.8
R6860 CSoutput.n76 CSoutput.n0 165.8
R6861 CSoutput.n75 CSoutput.n74 165.8
R6862 CSoutput.n73 CSoutput.n72 165.8
R6863 CSoutput.n71 CSoutput.n2 165.8
R6864 CSoutput.n69 CSoutput.n68 165.8
R6865 CSoutput.n67 CSoutput.n3 165.8
R6866 CSoutput.n66 CSoutput.n65 165.8
R6867 CSoutput.n63 CSoutput.n4 165.8
R6868 CSoutput.n61 CSoutput.n60 165.8
R6869 CSoutput.n59 CSoutput.n5 165.8
R6870 CSoutput.n58 CSoutput.n57 165.8
R6871 CSoutput.n55 CSoutput.n6 165.8
R6872 CSoutput.n54 CSoutput.n53 165.8
R6873 CSoutput.n52 CSoutput.n51 165.8
R6874 CSoutput.n50 CSoutput.n8 165.8
R6875 CSoutput.n48 CSoutput.n47 165.8
R6876 CSoutput.n46 CSoutput.n9 165.8
R6877 CSoutput.n45 CSoutput.n44 165.8
R6878 CSoutput.n42 CSoutput.n10 165.8
R6879 CSoutput.n41 CSoutput.n40 165.8
R6880 CSoutput.n39 CSoutput.n38 165.8
R6881 CSoutput.n37 CSoutput.n12 165.8
R6882 CSoutput.n35 CSoutput.n34 165.8
R6883 CSoutput.n33 CSoutput.n13 165.8
R6884 CSoutput.n32 CSoutput.n31 165.8
R6885 CSoutput.n29 CSoutput.n14 165.8
R6886 CSoutput.n28 CSoutput.n27 165.8
R6887 CSoutput.n26 CSoutput.n25 165.8
R6888 CSoutput.n24 CSoutput.n16 165.8
R6889 CSoutput.n22 CSoutput.n21 165.8
R6890 CSoutput.n20 CSoutput.n17 165.8
R6891 CSoutput.n77 CSoutput.t189 162.194
R6892 CSoutput.n18 CSoutput.t190 120.501
R6893 CSoutput.n23 CSoutput.t198 120.501
R6894 CSoutput.n15 CSoutput.t194 120.501
R6895 CSoutput.n30 CSoutput.t191 120.501
R6896 CSoutput.n36 CSoutput.t201 120.501
R6897 CSoutput.n11 CSoutput.t204 120.501
R6898 CSoutput.n43 CSoutput.t193 120.501
R6899 CSoutput.n49 CSoutput.t205 120.501
R6900 CSoutput.n7 CSoutput.t184 120.501
R6901 CSoutput.n56 CSoutput.t200 120.501
R6902 CSoutput.n62 CSoutput.t192 120.501
R6903 CSoutput.n64 CSoutput.t186 120.501
R6904 CSoutput.n70 CSoutput.t203 120.501
R6905 CSoutput.n1 CSoutput.t197 120.501
R6906 CSoutput.n330 CSoutput.n328 103.469
R6907 CSoutput.n310 CSoutput.n308 103.469
R6908 CSoutput.n291 CSoutput.n289 103.469
R6909 CSoutput.n120 CSoutput.n118 103.469
R6910 CSoutput.n100 CSoutput.n98 103.469
R6911 CSoutput.n81 CSoutput.n79 103.469
R6912 CSoutput.n344 CSoutput.n343 103.111
R6913 CSoutput.n342 CSoutput.n341 103.111
R6914 CSoutput.n340 CSoutput.n339 103.111
R6915 CSoutput.n338 CSoutput.n337 103.111
R6916 CSoutput.n336 CSoutput.n335 103.111
R6917 CSoutput.n334 CSoutput.n333 103.111
R6918 CSoutput.n332 CSoutput.n331 103.111
R6919 CSoutput.n330 CSoutput.n329 103.111
R6920 CSoutput.n326 CSoutput.n325 103.111
R6921 CSoutput.n324 CSoutput.n323 103.111
R6922 CSoutput.n322 CSoutput.n321 103.111
R6923 CSoutput.n320 CSoutput.n319 103.111
R6924 CSoutput.n318 CSoutput.n317 103.111
R6925 CSoutput.n316 CSoutput.n315 103.111
R6926 CSoutput.n314 CSoutput.n313 103.111
R6927 CSoutput.n312 CSoutput.n311 103.111
R6928 CSoutput.n310 CSoutput.n309 103.111
R6929 CSoutput.n307 CSoutput.n306 103.111
R6930 CSoutput.n305 CSoutput.n304 103.111
R6931 CSoutput.n303 CSoutput.n302 103.111
R6932 CSoutput.n301 CSoutput.n300 103.111
R6933 CSoutput.n299 CSoutput.n298 103.111
R6934 CSoutput.n297 CSoutput.n296 103.111
R6935 CSoutput.n295 CSoutput.n294 103.111
R6936 CSoutput.n293 CSoutput.n292 103.111
R6937 CSoutput.n291 CSoutput.n290 103.111
R6938 CSoutput.n120 CSoutput.n119 103.111
R6939 CSoutput.n122 CSoutput.n121 103.111
R6940 CSoutput.n124 CSoutput.n123 103.111
R6941 CSoutput.n126 CSoutput.n125 103.111
R6942 CSoutput.n128 CSoutput.n127 103.111
R6943 CSoutput.n130 CSoutput.n129 103.111
R6944 CSoutput.n132 CSoutput.n131 103.111
R6945 CSoutput.n134 CSoutput.n133 103.111
R6946 CSoutput.n136 CSoutput.n135 103.111
R6947 CSoutput.n100 CSoutput.n99 103.111
R6948 CSoutput.n102 CSoutput.n101 103.111
R6949 CSoutput.n104 CSoutput.n103 103.111
R6950 CSoutput.n106 CSoutput.n105 103.111
R6951 CSoutput.n108 CSoutput.n107 103.111
R6952 CSoutput.n110 CSoutput.n109 103.111
R6953 CSoutput.n112 CSoutput.n111 103.111
R6954 CSoutput.n114 CSoutput.n113 103.111
R6955 CSoutput.n116 CSoutput.n115 103.111
R6956 CSoutput.n81 CSoutput.n80 103.111
R6957 CSoutput.n83 CSoutput.n82 103.111
R6958 CSoutput.n85 CSoutput.n84 103.111
R6959 CSoutput.n87 CSoutput.n86 103.111
R6960 CSoutput.n89 CSoutput.n88 103.111
R6961 CSoutput.n91 CSoutput.n90 103.111
R6962 CSoutput.n93 CSoutput.n92 103.111
R6963 CSoutput.n95 CSoutput.n94 103.111
R6964 CSoutput.n97 CSoutput.n96 103.111
R6965 CSoutput.n346 CSoutput.n345 103.111
R6966 CSoutput.n366 CSoutput.n364 81.5057
R6967 CSoutput.n351 CSoutput.n349 81.5057
R6968 CSoutput.n398 CSoutput.n396 81.5057
R6969 CSoutput.n383 CSoutput.n381 81.5057
R6970 CSoutput.n378 CSoutput.n377 80.9324
R6971 CSoutput.n376 CSoutput.n375 80.9324
R6972 CSoutput.n374 CSoutput.n373 80.9324
R6973 CSoutput.n372 CSoutput.n371 80.9324
R6974 CSoutput.n370 CSoutput.n369 80.9324
R6975 CSoutput.n368 CSoutput.n367 80.9324
R6976 CSoutput.n366 CSoutput.n365 80.9324
R6977 CSoutput.n363 CSoutput.n362 80.9324
R6978 CSoutput.n361 CSoutput.n360 80.9324
R6979 CSoutput.n359 CSoutput.n358 80.9324
R6980 CSoutput.n357 CSoutput.n356 80.9324
R6981 CSoutput.n355 CSoutput.n354 80.9324
R6982 CSoutput.n353 CSoutput.n352 80.9324
R6983 CSoutput.n351 CSoutput.n350 80.9324
R6984 CSoutput.n398 CSoutput.n397 80.9324
R6985 CSoutput.n400 CSoutput.n399 80.9324
R6986 CSoutput.n402 CSoutput.n401 80.9324
R6987 CSoutput.n404 CSoutput.n403 80.9324
R6988 CSoutput.n406 CSoutput.n405 80.9324
R6989 CSoutput.n408 CSoutput.n407 80.9324
R6990 CSoutput.n410 CSoutput.n409 80.9324
R6991 CSoutput.n383 CSoutput.n382 80.9324
R6992 CSoutput.n385 CSoutput.n384 80.9324
R6993 CSoutput.n387 CSoutput.n386 80.9324
R6994 CSoutput.n389 CSoutput.n388 80.9324
R6995 CSoutput.n391 CSoutput.n390 80.9324
R6996 CSoutput.n393 CSoutput.n392 80.9324
R6997 CSoutput.n395 CSoutput.n394 80.9324
R6998 CSoutput.n25 CSoutput.n24 48.1486
R6999 CSoutput.n69 CSoutput.n3 48.1486
R7000 CSoutput.n38 CSoutput.n37 48.1486
R7001 CSoutput.n42 CSoutput.n41 48.1486
R7002 CSoutput.n51 CSoutput.n50 48.1486
R7003 CSoutput.n55 CSoutput.n54 48.1486
R7004 CSoutput.n22 CSoutput.n17 46.462
R7005 CSoutput.n72 CSoutput.n71 46.462
R7006 CSoutput.n20 CSoutput.n19 44.9055
R7007 CSoutput.n29 CSoutput.n28 43.7635
R7008 CSoutput.n65 CSoutput.n63 43.7635
R7009 CSoutput.n35 CSoutput.n13 41.7396
R7010 CSoutput.n57 CSoutput.n5 41.7396
R7011 CSoutput.n44 CSoutput.n9 37.0171
R7012 CSoutput.n48 CSoutput.n9 37.0171
R7013 CSoutput.n76 CSoutput.n75 34.9932
R7014 CSoutput.n31 CSoutput.n13 32.2947
R7015 CSoutput.n61 CSoutput.n5 32.2947
R7016 CSoutput.n30 CSoutput.n29 29.6014
R7017 CSoutput.n63 CSoutput.n62 29.6014
R7018 CSoutput.n19 CSoutput.n18 28.4085
R7019 CSoutput.n18 CSoutput.n17 25.1176
R7020 CSoutput.n72 CSoutput.n1 25.1176
R7021 CSoutput.n43 CSoutput.n42 22.0922
R7022 CSoutput.n50 CSoutput.n49 22.0922
R7023 CSoutput.n77 CSoutput.n76 21.8586
R7024 CSoutput.n37 CSoutput.n36 18.9681
R7025 CSoutput.n56 CSoutput.n55 18.9681
R7026 CSoutput.n25 CSoutput.n15 17.6292
R7027 CSoutput.n64 CSoutput.n3 17.6292
R7028 CSoutput.n24 CSoutput.n23 15.844
R7029 CSoutput.n70 CSoutput.n69 15.844
R7030 CSoutput.n38 CSoutput.n11 14.5051
R7031 CSoutput.n54 CSoutput.n7 14.5051
R7032 CSoutput.n413 CSoutput.n78 11.6139
R7033 CSoutput.n41 CSoutput.n11 11.3811
R7034 CSoutput.n51 CSoutput.n7 11.3811
R7035 CSoutput.n23 CSoutput.n22 10.0422
R7036 CSoutput.n71 CSoutput.n70 10.0422
R7037 CSoutput.n327 CSoutput.n307 9.25285
R7038 CSoutput.n117 CSoutput.n97 9.25285
R7039 CSoutput.n379 CSoutput.n363 8.97993
R7040 CSoutput.n411 CSoutput.n395 8.97993
R7041 CSoutput.n380 CSoutput.n348 8.71993
R7042 CSoutput.n28 CSoutput.n15 8.25698
R7043 CSoutput.n65 CSoutput.n64 8.25698
R7044 CSoutput.n380 CSoutput.n379 7.89345
R7045 CSoutput.n412 CSoutput.n411 7.89345
R7046 CSoutput.n348 CSoutput.n347 7.12641
R7047 CSoutput.n138 CSoutput.n137 7.12641
R7048 CSoutput.n36 CSoutput.n35 6.91809
R7049 CSoutput.n57 CSoutput.n56 6.91809
R7050 CSoutput.n379 CSoutput.n378 5.25266
R7051 CSoutput.n411 CSoutput.n410 5.25266
R7052 CSoutput.n347 CSoutput.n346 5.1449
R7053 CSoutput.n327 CSoutput.n326 5.1449
R7054 CSoutput.n137 CSoutput.n136 5.1449
R7055 CSoutput.n117 CSoutput.n116 5.1449
R7056 CSoutput.n413 CSoutput.n138 5.12749
R7057 CSoutput.n229 CSoutput.n182 4.5005
R7058 CSoutput.n198 CSoutput.n182 4.5005
R7059 CSoutput.n193 CSoutput.n177 4.5005
R7060 CSoutput.n193 CSoutput.n179 4.5005
R7061 CSoutput.n193 CSoutput.n176 4.5005
R7062 CSoutput.n193 CSoutput.n180 4.5005
R7063 CSoutput.n193 CSoutput.n175 4.5005
R7064 CSoutput.n193 CSoutput.t199 4.5005
R7065 CSoutput.n193 CSoutput.n174 4.5005
R7066 CSoutput.n193 CSoutput.n181 4.5005
R7067 CSoutput.n193 CSoutput.n182 4.5005
R7068 CSoutput.n191 CSoutput.n177 4.5005
R7069 CSoutput.n191 CSoutput.n179 4.5005
R7070 CSoutput.n191 CSoutput.n176 4.5005
R7071 CSoutput.n191 CSoutput.n180 4.5005
R7072 CSoutput.n191 CSoutput.n175 4.5005
R7073 CSoutput.n191 CSoutput.t199 4.5005
R7074 CSoutput.n191 CSoutput.n174 4.5005
R7075 CSoutput.n191 CSoutput.n181 4.5005
R7076 CSoutput.n191 CSoutput.n182 4.5005
R7077 CSoutput.n190 CSoutput.n177 4.5005
R7078 CSoutput.n190 CSoutput.n179 4.5005
R7079 CSoutput.n190 CSoutput.n176 4.5005
R7080 CSoutput.n190 CSoutput.n180 4.5005
R7081 CSoutput.n190 CSoutput.n175 4.5005
R7082 CSoutput.n190 CSoutput.t199 4.5005
R7083 CSoutput.n190 CSoutput.n174 4.5005
R7084 CSoutput.n190 CSoutput.n181 4.5005
R7085 CSoutput.n190 CSoutput.n182 4.5005
R7086 CSoutput.n275 CSoutput.n177 4.5005
R7087 CSoutput.n275 CSoutput.n179 4.5005
R7088 CSoutput.n275 CSoutput.n176 4.5005
R7089 CSoutput.n275 CSoutput.n180 4.5005
R7090 CSoutput.n275 CSoutput.n175 4.5005
R7091 CSoutput.n275 CSoutput.t199 4.5005
R7092 CSoutput.n275 CSoutput.n174 4.5005
R7093 CSoutput.n275 CSoutput.n181 4.5005
R7094 CSoutput.n275 CSoutput.n182 4.5005
R7095 CSoutput.n273 CSoutput.n177 4.5005
R7096 CSoutput.n273 CSoutput.n179 4.5005
R7097 CSoutput.n273 CSoutput.n176 4.5005
R7098 CSoutput.n273 CSoutput.n180 4.5005
R7099 CSoutput.n273 CSoutput.n175 4.5005
R7100 CSoutput.n273 CSoutput.t199 4.5005
R7101 CSoutput.n273 CSoutput.n174 4.5005
R7102 CSoutput.n273 CSoutput.n181 4.5005
R7103 CSoutput.n271 CSoutput.n177 4.5005
R7104 CSoutput.n271 CSoutput.n179 4.5005
R7105 CSoutput.n271 CSoutput.n176 4.5005
R7106 CSoutput.n271 CSoutput.n180 4.5005
R7107 CSoutput.n271 CSoutput.n175 4.5005
R7108 CSoutput.n271 CSoutput.t199 4.5005
R7109 CSoutput.n271 CSoutput.n174 4.5005
R7110 CSoutput.n271 CSoutput.n181 4.5005
R7111 CSoutput.n201 CSoutput.n177 4.5005
R7112 CSoutput.n201 CSoutput.n179 4.5005
R7113 CSoutput.n201 CSoutput.n176 4.5005
R7114 CSoutput.n201 CSoutput.n180 4.5005
R7115 CSoutput.n201 CSoutput.n175 4.5005
R7116 CSoutput.n201 CSoutput.t199 4.5005
R7117 CSoutput.n201 CSoutput.n174 4.5005
R7118 CSoutput.n201 CSoutput.n181 4.5005
R7119 CSoutput.n201 CSoutput.n182 4.5005
R7120 CSoutput.n200 CSoutput.n177 4.5005
R7121 CSoutput.n200 CSoutput.n179 4.5005
R7122 CSoutput.n200 CSoutput.n176 4.5005
R7123 CSoutput.n200 CSoutput.n180 4.5005
R7124 CSoutput.n200 CSoutput.n175 4.5005
R7125 CSoutput.n200 CSoutput.t199 4.5005
R7126 CSoutput.n200 CSoutput.n174 4.5005
R7127 CSoutput.n200 CSoutput.n181 4.5005
R7128 CSoutput.n200 CSoutput.n182 4.5005
R7129 CSoutput.n204 CSoutput.n177 4.5005
R7130 CSoutput.n204 CSoutput.n179 4.5005
R7131 CSoutput.n204 CSoutput.n176 4.5005
R7132 CSoutput.n204 CSoutput.n180 4.5005
R7133 CSoutput.n204 CSoutput.n175 4.5005
R7134 CSoutput.n204 CSoutput.t199 4.5005
R7135 CSoutput.n204 CSoutput.n174 4.5005
R7136 CSoutput.n204 CSoutput.n181 4.5005
R7137 CSoutput.n204 CSoutput.n182 4.5005
R7138 CSoutput.n203 CSoutput.n177 4.5005
R7139 CSoutput.n203 CSoutput.n179 4.5005
R7140 CSoutput.n203 CSoutput.n176 4.5005
R7141 CSoutput.n203 CSoutput.n180 4.5005
R7142 CSoutput.n203 CSoutput.n175 4.5005
R7143 CSoutput.n203 CSoutput.t199 4.5005
R7144 CSoutput.n203 CSoutput.n174 4.5005
R7145 CSoutput.n203 CSoutput.n181 4.5005
R7146 CSoutput.n203 CSoutput.n182 4.5005
R7147 CSoutput.n186 CSoutput.n177 4.5005
R7148 CSoutput.n186 CSoutput.n179 4.5005
R7149 CSoutput.n186 CSoutput.n176 4.5005
R7150 CSoutput.n186 CSoutput.n180 4.5005
R7151 CSoutput.n186 CSoutput.n175 4.5005
R7152 CSoutput.n186 CSoutput.t199 4.5005
R7153 CSoutput.n186 CSoutput.n174 4.5005
R7154 CSoutput.n186 CSoutput.n181 4.5005
R7155 CSoutput.n186 CSoutput.n182 4.5005
R7156 CSoutput.n278 CSoutput.n177 4.5005
R7157 CSoutput.n278 CSoutput.n179 4.5005
R7158 CSoutput.n278 CSoutput.n176 4.5005
R7159 CSoutput.n278 CSoutput.n180 4.5005
R7160 CSoutput.n278 CSoutput.n175 4.5005
R7161 CSoutput.n278 CSoutput.t199 4.5005
R7162 CSoutput.n278 CSoutput.n174 4.5005
R7163 CSoutput.n278 CSoutput.n181 4.5005
R7164 CSoutput.n278 CSoutput.n182 4.5005
R7165 CSoutput.n265 CSoutput.n236 4.5005
R7166 CSoutput.n265 CSoutput.n242 4.5005
R7167 CSoutput.n223 CSoutput.n212 4.5005
R7168 CSoutput.n223 CSoutput.n214 4.5005
R7169 CSoutput.n223 CSoutput.n211 4.5005
R7170 CSoutput.n223 CSoutput.n215 4.5005
R7171 CSoutput.n223 CSoutput.n210 4.5005
R7172 CSoutput.n223 CSoutput.t195 4.5005
R7173 CSoutput.n223 CSoutput.n209 4.5005
R7174 CSoutput.n223 CSoutput.n216 4.5005
R7175 CSoutput.n265 CSoutput.n223 4.5005
R7176 CSoutput.n244 CSoutput.n212 4.5005
R7177 CSoutput.n244 CSoutput.n214 4.5005
R7178 CSoutput.n244 CSoutput.n211 4.5005
R7179 CSoutput.n244 CSoutput.n215 4.5005
R7180 CSoutput.n244 CSoutput.n210 4.5005
R7181 CSoutput.n244 CSoutput.t195 4.5005
R7182 CSoutput.n244 CSoutput.n209 4.5005
R7183 CSoutput.n244 CSoutput.n216 4.5005
R7184 CSoutput.n265 CSoutput.n244 4.5005
R7185 CSoutput.n222 CSoutput.n212 4.5005
R7186 CSoutput.n222 CSoutput.n214 4.5005
R7187 CSoutput.n222 CSoutput.n211 4.5005
R7188 CSoutput.n222 CSoutput.n215 4.5005
R7189 CSoutput.n222 CSoutput.n210 4.5005
R7190 CSoutput.n222 CSoutput.t195 4.5005
R7191 CSoutput.n222 CSoutput.n209 4.5005
R7192 CSoutput.n222 CSoutput.n216 4.5005
R7193 CSoutput.n265 CSoutput.n222 4.5005
R7194 CSoutput.n246 CSoutput.n212 4.5005
R7195 CSoutput.n246 CSoutput.n214 4.5005
R7196 CSoutput.n246 CSoutput.n211 4.5005
R7197 CSoutput.n246 CSoutput.n215 4.5005
R7198 CSoutput.n246 CSoutput.n210 4.5005
R7199 CSoutput.n246 CSoutput.t195 4.5005
R7200 CSoutput.n246 CSoutput.n209 4.5005
R7201 CSoutput.n246 CSoutput.n216 4.5005
R7202 CSoutput.n265 CSoutput.n246 4.5005
R7203 CSoutput.n212 CSoutput.n207 4.5005
R7204 CSoutput.n214 CSoutput.n207 4.5005
R7205 CSoutput.n211 CSoutput.n207 4.5005
R7206 CSoutput.n215 CSoutput.n207 4.5005
R7207 CSoutput.n210 CSoutput.n207 4.5005
R7208 CSoutput.t195 CSoutput.n207 4.5005
R7209 CSoutput.n209 CSoutput.n207 4.5005
R7210 CSoutput.n216 CSoutput.n207 4.5005
R7211 CSoutput.n268 CSoutput.n212 4.5005
R7212 CSoutput.n268 CSoutput.n214 4.5005
R7213 CSoutput.n268 CSoutput.n211 4.5005
R7214 CSoutput.n268 CSoutput.n215 4.5005
R7215 CSoutput.n268 CSoutput.n210 4.5005
R7216 CSoutput.n268 CSoutput.t195 4.5005
R7217 CSoutput.n268 CSoutput.n209 4.5005
R7218 CSoutput.n268 CSoutput.n216 4.5005
R7219 CSoutput.n266 CSoutput.n212 4.5005
R7220 CSoutput.n266 CSoutput.n214 4.5005
R7221 CSoutput.n266 CSoutput.n211 4.5005
R7222 CSoutput.n266 CSoutput.n215 4.5005
R7223 CSoutput.n266 CSoutput.n210 4.5005
R7224 CSoutput.n266 CSoutput.t195 4.5005
R7225 CSoutput.n266 CSoutput.n209 4.5005
R7226 CSoutput.n266 CSoutput.n216 4.5005
R7227 CSoutput.n266 CSoutput.n265 4.5005
R7228 CSoutput.n248 CSoutput.n212 4.5005
R7229 CSoutput.n248 CSoutput.n214 4.5005
R7230 CSoutput.n248 CSoutput.n211 4.5005
R7231 CSoutput.n248 CSoutput.n215 4.5005
R7232 CSoutput.n248 CSoutput.n210 4.5005
R7233 CSoutput.n248 CSoutput.t195 4.5005
R7234 CSoutput.n248 CSoutput.n209 4.5005
R7235 CSoutput.n248 CSoutput.n216 4.5005
R7236 CSoutput.n265 CSoutput.n248 4.5005
R7237 CSoutput.n220 CSoutput.n212 4.5005
R7238 CSoutput.n220 CSoutput.n214 4.5005
R7239 CSoutput.n220 CSoutput.n211 4.5005
R7240 CSoutput.n220 CSoutput.n215 4.5005
R7241 CSoutput.n220 CSoutput.n210 4.5005
R7242 CSoutput.n220 CSoutput.t195 4.5005
R7243 CSoutput.n220 CSoutput.n209 4.5005
R7244 CSoutput.n220 CSoutput.n216 4.5005
R7245 CSoutput.n265 CSoutput.n220 4.5005
R7246 CSoutput.n250 CSoutput.n212 4.5005
R7247 CSoutput.n250 CSoutput.n214 4.5005
R7248 CSoutput.n250 CSoutput.n211 4.5005
R7249 CSoutput.n250 CSoutput.n215 4.5005
R7250 CSoutput.n250 CSoutput.n210 4.5005
R7251 CSoutput.n250 CSoutput.t195 4.5005
R7252 CSoutput.n250 CSoutput.n209 4.5005
R7253 CSoutput.n250 CSoutput.n216 4.5005
R7254 CSoutput.n265 CSoutput.n250 4.5005
R7255 CSoutput.n219 CSoutput.n212 4.5005
R7256 CSoutput.n219 CSoutput.n214 4.5005
R7257 CSoutput.n219 CSoutput.n211 4.5005
R7258 CSoutput.n219 CSoutput.n215 4.5005
R7259 CSoutput.n219 CSoutput.n210 4.5005
R7260 CSoutput.n219 CSoutput.t195 4.5005
R7261 CSoutput.n219 CSoutput.n209 4.5005
R7262 CSoutput.n219 CSoutput.n216 4.5005
R7263 CSoutput.n265 CSoutput.n219 4.5005
R7264 CSoutput.n264 CSoutput.n212 4.5005
R7265 CSoutput.n264 CSoutput.n214 4.5005
R7266 CSoutput.n264 CSoutput.n211 4.5005
R7267 CSoutput.n264 CSoutput.n215 4.5005
R7268 CSoutput.n264 CSoutput.n210 4.5005
R7269 CSoutput.n264 CSoutput.t195 4.5005
R7270 CSoutput.n264 CSoutput.n209 4.5005
R7271 CSoutput.n264 CSoutput.n216 4.5005
R7272 CSoutput.n265 CSoutput.n264 4.5005
R7273 CSoutput.n263 CSoutput.n148 4.5005
R7274 CSoutput.n164 CSoutput.n148 4.5005
R7275 CSoutput.n159 CSoutput.n143 4.5005
R7276 CSoutput.n159 CSoutput.n145 4.5005
R7277 CSoutput.n159 CSoutput.n142 4.5005
R7278 CSoutput.n159 CSoutput.n146 4.5005
R7279 CSoutput.n159 CSoutput.n141 4.5005
R7280 CSoutput.n159 CSoutput.t185 4.5005
R7281 CSoutput.n159 CSoutput.n140 4.5005
R7282 CSoutput.n159 CSoutput.n147 4.5005
R7283 CSoutput.n159 CSoutput.n148 4.5005
R7284 CSoutput.n157 CSoutput.n143 4.5005
R7285 CSoutput.n157 CSoutput.n145 4.5005
R7286 CSoutput.n157 CSoutput.n142 4.5005
R7287 CSoutput.n157 CSoutput.n146 4.5005
R7288 CSoutput.n157 CSoutput.n141 4.5005
R7289 CSoutput.n157 CSoutput.t185 4.5005
R7290 CSoutput.n157 CSoutput.n140 4.5005
R7291 CSoutput.n157 CSoutput.n147 4.5005
R7292 CSoutput.n157 CSoutput.n148 4.5005
R7293 CSoutput.n156 CSoutput.n143 4.5005
R7294 CSoutput.n156 CSoutput.n145 4.5005
R7295 CSoutput.n156 CSoutput.n142 4.5005
R7296 CSoutput.n156 CSoutput.n146 4.5005
R7297 CSoutput.n156 CSoutput.n141 4.5005
R7298 CSoutput.n156 CSoutput.t185 4.5005
R7299 CSoutput.n156 CSoutput.n140 4.5005
R7300 CSoutput.n156 CSoutput.n147 4.5005
R7301 CSoutput.n156 CSoutput.n148 4.5005
R7302 CSoutput.n285 CSoutput.n143 4.5005
R7303 CSoutput.n285 CSoutput.n145 4.5005
R7304 CSoutput.n285 CSoutput.n142 4.5005
R7305 CSoutput.n285 CSoutput.n146 4.5005
R7306 CSoutput.n285 CSoutput.n141 4.5005
R7307 CSoutput.n285 CSoutput.t185 4.5005
R7308 CSoutput.n285 CSoutput.n140 4.5005
R7309 CSoutput.n285 CSoutput.n147 4.5005
R7310 CSoutput.n285 CSoutput.n148 4.5005
R7311 CSoutput.n283 CSoutput.n143 4.5005
R7312 CSoutput.n283 CSoutput.n145 4.5005
R7313 CSoutput.n283 CSoutput.n142 4.5005
R7314 CSoutput.n283 CSoutput.n146 4.5005
R7315 CSoutput.n283 CSoutput.n141 4.5005
R7316 CSoutput.n283 CSoutput.t185 4.5005
R7317 CSoutput.n283 CSoutput.n140 4.5005
R7318 CSoutput.n283 CSoutput.n147 4.5005
R7319 CSoutput.n281 CSoutput.n143 4.5005
R7320 CSoutput.n281 CSoutput.n145 4.5005
R7321 CSoutput.n281 CSoutput.n142 4.5005
R7322 CSoutput.n281 CSoutput.n146 4.5005
R7323 CSoutput.n281 CSoutput.n141 4.5005
R7324 CSoutput.n281 CSoutput.t185 4.5005
R7325 CSoutput.n281 CSoutput.n140 4.5005
R7326 CSoutput.n281 CSoutput.n147 4.5005
R7327 CSoutput.n167 CSoutput.n143 4.5005
R7328 CSoutput.n167 CSoutput.n145 4.5005
R7329 CSoutput.n167 CSoutput.n142 4.5005
R7330 CSoutput.n167 CSoutput.n146 4.5005
R7331 CSoutput.n167 CSoutput.n141 4.5005
R7332 CSoutput.n167 CSoutput.t185 4.5005
R7333 CSoutput.n167 CSoutput.n140 4.5005
R7334 CSoutput.n167 CSoutput.n147 4.5005
R7335 CSoutput.n167 CSoutput.n148 4.5005
R7336 CSoutput.n166 CSoutput.n143 4.5005
R7337 CSoutput.n166 CSoutput.n145 4.5005
R7338 CSoutput.n166 CSoutput.n142 4.5005
R7339 CSoutput.n166 CSoutput.n146 4.5005
R7340 CSoutput.n166 CSoutput.n141 4.5005
R7341 CSoutput.n166 CSoutput.t185 4.5005
R7342 CSoutput.n166 CSoutput.n140 4.5005
R7343 CSoutput.n166 CSoutput.n147 4.5005
R7344 CSoutput.n166 CSoutput.n148 4.5005
R7345 CSoutput.n170 CSoutput.n143 4.5005
R7346 CSoutput.n170 CSoutput.n145 4.5005
R7347 CSoutput.n170 CSoutput.n142 4.5005
R7348 CSoutput.n170 CSoutput.n146 4.5005
R7349 CSoutput.n170 CSoutput.n141 4.5005
R7350 CSoutput.n170 CSoutput.t185 4.5005
R7351 CSoutput.n170 CSoutput.n140 4.5005
R7352 CSoutput.n170 CSoutput.n147 4.5005
R7353 CSoutput.n170 CSoutput.n148 4.5005
R7354 CSoutput.n169 CSoutput.n143 4.5005
R7355 CSoutput.n169 CSoutput.n145 4.5005
R7356 CSoutput.n169 CSoutput.n142 4.5005
R7357 CSoutput.n169 CSoutput.n146 4.5005
R7358 CSoutput.n169 CSoutput.n141 4.5005
R7359 CSoutput.n169 CSoutput.t185 4.5005
R7360 CSoutput.n169 CSoutput.n140 4.5005
R7361 CSoutput.n169 CSoutput.n147 4.5005
R7362 CSoutput.n169 CSoutput.n148 4.5005
R7363 CSoutput.n152 CSoutput.n143 4.5005
R7364 CSoutput.n152 CSoutput.n145 4.5005
R7365 CSoutput.n152 CSoutput.n142 4.5005
R7366 CSoutput.n152 CSoutput.n146 4.5005
R7367 CSoutput.n152 CSoutput.n141 4.5005
R7368 CSoutput.n152 CSoutput.t185 4.5005
R7369 CSoutput.n152 CSoutput.n140 4.5005
R7370 CSoutput.n152 CSoutput.n147 4.5005
R7371 CSoutput.n152 CSoutput.n148 4.5005
R7372 CSoutput.n288 CSoutput.n143 4.5005
R7373 CSoutput.n288 CSoutput.n145 4.5005
R7374 CSoutput.n288 CSoutput.n142 4.5005
R7375 CSoutput.n288 CSoutput.n146 4.5005
R7376 CSoutput.n288 CSoutput.n141 4.5005
R7377 CSoutput.n288 CSoutput.t185 4.5005
R7378 CSoutput.n288 CSoutput.n140 4.5005
R7379 CSoutput.n288 CSoutput.n147 4.5005
R7380 CSoutput.n288 CSoutput.n148 4.5005
R7381 CSoutput.n347 CSoutput.n327 4.10845
R7382 CSoutput.n137 CSoutput.n117 4.10845
R7383 CSoutput.n345 CSoutput.t165 4.06363
R7384 CSoutput.n345 CSoutput.t77 4.06363
R7385 CSoutput.n343 CSoutput.t101 4.06363
R7386 CSoutput.n343 CSoutput.t128 4.06363
R7387 CSoutput.n341 CSoutput.t145 4.06363
R7388 CSoutput.n341 CSoutput.t62 4.06363
R7389 CSoutput.n339 CSoutput.t56 4.06363
R7390 CSoutput.n339 CSoutput.t104 4.06363
R7391 CSoutput.n337 CSoutput.t122 4.06363
R7392 CSoutput.n337 CSoutput.t147 4.06363
R7393 CSoutput.n335 CSoutput.t162 4.06363
R7394 CSoutput.n335 CSoutput.t74 4.06363
R7395 CSoutput.n333 CSoutput.t80 4.06363
R7396 CSoutput.n333 CSoutput.t148 4.06363
R7397 CSoutput.n331 CSoutput.t164 4.06363
R7398 CSoutput.n331 CSoutput.t166 4.06363
R7399 CSoutput.n329 CSoutput.t100 4.06363
R7400 CSoutput.n329 CSoutput.t102 4.06363
R7401 CSoutput.n328 CSoutput.t106 4.06363
R7402 CSoutput.n328 CSoutput.t170 4.06363
R7403 CSoutput.n325 CSoutput.t154 4.06363
R7404 CSoutput.n325 CSoutput.t63 4.06363
R7405 CSoutput.n323 CSoutput.t83 4.06363
R7406 CSoutput.n323 CSoutput.t120 4.06363
R7407 CSoutput.n321 CSoutput.t135 4.06363
R7408 CSoutput.n321 CSoutput.t171 4.06363
R7409 CSoutput.n319 CSoutput.t163 4.06363
R7410 CSoutput.n319 CSoutput.t89 4.06363
R7411 CSoutput.n317 CSoutput.t109 4.06363
R7412 CSoutput.n317 CSoutput.t136 4.06363
R7413 CSoutput.n315 CSoutput.t149 4.06363
R7414 CSoutput.n315 CSoutput.t61 4.06363
R7415 CSoutput.n313 CSoutput.t64 4.06363
R7416 CSoutput.n313 CSoutput.t139 4.06363
R7417 CSoutput.n311 CSoutput.t155 4.06363
R7418 CSoutput.n311 CSoutput.t156 4.06363
R7419 CSoutput.n309 CSoutput.t82 4.06363
R7420 CSoutput.n309 CSoutput.t84 4.06363
R7421 CSoutput.n308 CSoutput.t90 4.06363
R7422 CSoutput.n308 CSoutput.t158 4.06363
R7423 CSoutput.n306 CSoutput.t167 4.06363
R7424 CSoutput.n306 CSoutput.t121 4.06363
R7425 CSoutput.n304 CSoutput.t152 4.06363
R7426 CSoutput.n304 CSoutput.t105 4.06363
R7427 CSoutput.n302 CSoutput.t137 4.06363
R7428 CSoutput.n302 CSoutput.t87 4.06363
R7429 CSoutput.n300 CSoutput.t159 4.06363
R7430 CSoutput.n300 CSoutput.t113 4.06363
R7431 CSoutput.n298 CSoutput.t146 4.06363
R7432 CSoutput.n298 CSoutput.t97 4.06363
R7433 CSoutput.n296 CSoutput.t132 4.06363
R7434 CSoutput.n296 CSoutput.t73 4.06363
R7435 CSoutput.n294 CSoutput.t150 4.06363
R7436 CSoutput.n294 CSoutput.t68 4.06363
R7437 CSoutput.n292 CSoutput.t110 4.06363
R7438 CSoutput.n292 CSoutput.t85 4.06363
R7439 CSoutput.n290 CSoutput.t91 4.06363
R7440 CSoutput.n290 CSoutput.t65 4.06363
R7441 CSoutput.n289 CSoutput.t144 4.06363
R7442 CSoutput.n289 CSoutput.t58 4.06363
R7443 CSoutput.n118 CSoutput.t99 4.06363
R7444 CSoutput.n118 CSoutput.t173 4.06363
R7445 CSoutput.n119 CSoutput.t142 4.06363
R7446 CSoutput.n119 CSoutput.t140 4.06363
R7447 CSoutput.n121 CSoutput.t125 4.06363
R7448 CSoutput.n121 CSoutput.t95 4.06363
R7449 CSoutput.n123 CSoutput.t72 4.06363
R7450 CSoutput.n123 CSoutput.t127 4.06363
R7451 CSoutput.n125 CSoutput.t124 4.06363
R7452 CSoutput.n125 CSoutput.t92 4.06363
R7453 CSoutput.n127 CSoutput.t71 4.06363
R7454 CSoutput.n127 CSoutput.t70 4.06363
R7455 CSoutput.n129 CSoutput.t143 4.06363
R7456 CSoutput.n129 CSoutput.t108 4.06363
R7457 CSoutput.n131 CSoutput.t103 4.06363
R7458 CSoutput.n131 CSoutput.t66 4.06363
R7459 CSoutput.n133 CSoutput.t169 4.06363
R7460 CSoutput.n133 CSoutput.t141 4.06363
R7461 CSoutput.n135 CSoutput.t126 4.06363
R7462 CSoutput.n135 CSoutput.t96 4.06363
R7463 CSoutput.n98 CSoutput.t81 4.06363
R7464 CSoutput.n98 CSoutput.t161 4.06363
R7465 CSoutput.n99 CSoutput.t131 4.06363
R7466 CSoutput.n99 CSoutput.t129 4.06363
R7467 CSoutput.n101 CSoutput.t115 4.06363
R7468 CSoutput.n101 CSoutput.t78 4.06363
R7469 CSoutput.n103 CSoutput.t59 4.06363
R7470 CSoutput.n103 CSoutput.t117 4.06363
R7471 CSoutput.n105 CSoutput.t112 4.06363
R7472 CSoutput.n105 CSoutput.t75 4.06363
R7473 CSoutput.n107 CSoutput.t57 4.06363
R7474 CSoutput.n107 CSoutput.t55 4.06363
R7475 CSoutput.n109 CSoutput.t134 4.06363
R7476 CSoutput.n109 CSoutput.t94 4.06363
R7477 CSoutput.n111 CSoutput.t88 4.06363
R7478 CSoutput.n111 CSoutput.t54 4.06363
R7479 CSoutput.n113 CSoutput.t157 4.06363
R7480 CSoutput.n113 CSoutput.t130 4.06363
R7481 CSoutput.n115 CSoutput.t116 4.06363
R7482 CSoutput.n115 CSoutput.t79 4.06363
R7483 CSoutput.n79 CSoutput.t60 4.06363
R7484 CSoutput.n79 CSoutput.t118 4.06363
R7485 CSoutput.n80 CSoutput.t67 4.06363
R7486 CSoutput.n80 CSoutput.t93 4.06363
R7487 CSoutput.n82 CSoutput.t172 4.06363
R7488 CSoutput.n82 CSoutput.t111 4.06363
R7489 CSoutput.n84 CSoutput.t69 4.06363
R7490 CSoutput.n84 CSoutput.t151 4.06363
R7491 CSoutput.n86 CSoutput.t76 4.06363
R7492 CSoutput.n86 CSoutput.t133 4.06363
R7493 CSoutput.n88 CSoutput.t98 4.06363
R7494 CSoutput.n88 CSoutput.t119 4.06363
R7495 CSoutput.n90 CSoutput.t114 4.06363
R7496 CSoutput.n90 CSoutput.t160 4.06363
R7497 CSoutput.n92 CSoutput.t86 4.06363
R7498 CSoutput.n92 CSoutput.t138 4.06363
R7499 CSoutput.n94 CSoutput.t107 4.06363
R7500 CSoutput.n94 CSoutput.t153 4.06363
R7501 CSoutput.n96 CSoutput.t123 4.06363
R7502 CSoutput.n96 CSoutput.t168 4.06363
R7503 CSoutput.n44 CSoutput.n43 3.79402
R7504 CSoutput.n49 CSoutput.n48 3.79402
R7505 CSoutput.n413 CSoutput.n412 3.57343
R7506 CSoutput.n412 CSoutput.n380 3.3798
R7507 CSoutput.n348 CSoutput.n138 2.99158
R7508 CSoutput.n377 CSoutput.t43 2.82907
R7509 CSoutput.n377 CSoutput.t31 2.82907
R7510 CSoutput.n375 CSoutput.t42 2.82907
R7511 CSoutput.n375 CSoutput.t40 2.82907
R7512 CSoutput.n373 CSoutput.t7 2.82907
R7513 CSoutput.n373 CSoutput.t49 2.82907
R7514 CSoutput.n371 CSoutput.t36 2.82907
R7515 CSoutput.n371 CSoutput.t38 2.82907
R7516 CSoutput.n369 CSoutput.t21 2.82907
R7517 CSoutput.n369 CSoutput.t22 2.82907
R7518 CSoutput.n367 CSoutput.t181 2.82907
R7519 CSoutput.n367 CSoutput.t52 2.82907
R7520 CSoutput.n365 CSoutput.t29 2.82907
R7521 CSoutput.n365 CSoutput.t20 2.82907
R7522 CSoutput.n364 CSoutput.t17 2.82907
R7523 CSoutput.n364 CSoutput.t24 2.82907
R7524 CSoutput.n362 CSoutput.t1 2.82907
R7525 CSoutput.n362 CSoutput.t41 2.82907
R7526 CSoutput.n360 CSoutput.t53 2.82907
R7527 CSoutput.n360 CSoutput.t37 2.82907
R7528 CSoutput.n358 CSoutput.t45 2.82907
R7529 CSoutput.n358 CSoutput.t5 2.82907
R7530 CSoutput.n356 CSoutput.t35 2.82907
R7531 CSoutput.n356 CSoutput.t175 2.82907
R7532 CSoutput.n354 CSoutput.t51 2.82907
R7533 CSoutput.n354 CSoutput.t19 2.82907
R7534 CSoutput.n352 CSoutput.t0 2.82907
R7535 CSoutput.n352 CSoutput.t180 2.82907
R7536 CSoutput.n350 CSoutput.t176 2.82907
R7537 CSoutput.n350 CSoutput.t16 2.82907
R7538 CSoutput.n349 CSoutput.t4 2.82907
R7539 CSoutput.n349 CSoutput.t23 2.82907
R7540 CSoutput.n396 CSoutput.t26 2.82907
R7541 CSoutput.n396 CSoutput.t2 2.82907
R7542 CSoutput.n397 CSoutput.t6 2.82907
R7543 CSoutput.n397 CSoutput.t13 2.82907
R7544 CSoutput.n399 CSoutput.t177 2.82907
R7545 CSoutput.n399 CSoutput.t3 2.82907
R7546 CSoutput.n401 CSoutput.t18 2.82907
R7547 CSoutput.n401 CSoutput.t48 2.82907
R7548 CSoutput.n403 CSoutput.t8 2.82907
R7549 CSoutput.n403 CSoutput.t27 2.82907
R7550 CSoutput.n405 CSoutput.t182 2.82907
R7551 CSoutput.n405 CSoutput.t34 2.82907
R7552 CSoutput.n407 CSoutput.t179 2.82907
R7553 CSoutput.n407 CSoutput.t39 2.82907
R7554 CSoutput.n409 CSoutput.t10 2.82907
R7555 CSoutput.n409 CSoutput.t32 2.82907
R7556 CSoutput.n381 CSoutput.t9 2.82907
R7557 CSoutput.n381 CSoutput.t28 2.82907
R7558 CSoutput.n382 CSoutput.t30 2.82907
R7559 CSoutput.n382 CSoutput.t46 2.82907
R7560 CSoutput.n384 CSoutput.t47 2.82907
R7561 CSoutput.n384 CSoutput.t174 2.82907
R7562 CSoutput.n386 CSoutput.t15 2.82907
R7563 CSoutput.n386 CSoutput.t44 2.82907
R7564 CSoutput.n388 CSoutput.t11 2.82907
R7565 CSoutput.n388 CSoutput.t14 2.82907
R7566 CSoutput.n390 CSoutput.t178 2.82907
R7567 CSoutput.n390 CSoutput.t33 2.82907
R7568 CSoutput.n392 CSoutput.t12 2.82907
R7569 CSoutput.n392 CSoutput.t25 2.82907
R7570 CSoutput.n394 CSoutput.t183 2.82907
R7571 CSoutput.n394 CSoutput.t50 2.82907
R7572 CSoutput.n75 CSoutput.n1 2.45513
R7573 CSoutput.n229 CSoutput.n227 2.251
R7574 CSoutput.n229 CSoutput.n226 2.251
R7575 CSoutput.n229 CSoutput.n225 2.251
R7576 CSoutput.n229 CSoutput.n224 2.251
R7577 CSoutput.n198 CSoutput.n197 2.251
R7578 CSoutput.n198 CSoutput.n196 2.251
R7579 CSoutput.n198 CSoutput.n195 2.251
R7580 CSoutput.n198 CSoutput.n194 2.251
R7581 CSoutput.n271 CSoutput.n270 2.251
R7582 CSoutput.n236 CSoutput.n234 2.251
R7583 CSoutput.n236 CSoutput.n233 2.251
R7584 CSoutput.n236 CSoutput.n232 2.251
R7585 CSoutput.n254 CSoutput.n236 2.251
R7586 CSoutput.n242 CSoutput.n241 2.251
R7587 CSoutput.n242 CSoutput.n240 2.251
R7588 CSoutput.n242 CSoutput.n239 2.251
R7589 CSoutput.n242 CSoutput.n238 2.251
R7590 CSoutput.n268 CSoutput.n208 2.251
R7591 CSoutput.n263 CSoutput.n261 2.251
R7592 CSoutput.n263 CSoutput.n260 2.251
R7593 CSoutput.n263 CSoutput.n259 2.251
R7594 CSoutput.n263 CSoutput.n258 2.251
R7595 CSoutput.n164 CSoutput.n163 2.251
R7596 CSoutput.n164 CSoutput.n162 2.251
R7597 CSoutput.n164 CSoutput.n161 2.251
R7598 CSoutput.n164 CSoutput.n160 2.251
R7599 CSoutput.n281 CSoutput.n280 2.251
R7600 CSoutput.n198 CSoutput.n178 2.2505
R7601 CSoutput.n193 CSoutput.n178 2.2505
R7602 CSoutput.n191 CSoutput.n178 2.2505
R7603 CSoutput.n190 CSoutput.n178 2.2505
R7604 CSoutput.n275 CSoutput.n178 2.2505
R7605 CSoutput.n273 CSoutput.n178 2.2505
R7606 CSoutput.n271 CSoutput.n178 2.2505
R7607 CSoutput.n201 CSoutput.n178 2.2505
R7608 CSoutput.n200 CSoutput.n178 2.2505
R7609 CSoutput.n204 CSoutput.n178 2.2505
R7610 CSoutput.n203 CSoutput.n178 2.2505
R7611 CSoutput.n186 CSoutput.n178 2.2505
R7612 CSoutput.n278 CSoutput.n178 2.2505
R7613 CSoutput.n278 CSoutput.n277 2.2505
R7614 CSoutput.n242 CSoutput.n213 2.2505
R7615 CSoutput.n223 CSoutput.n213 2.2505
R7616 CSoutput.n244 CSoutput.n213 2.2505
R7617 CSoutput.n222 CSoutput.n213 2.2505
R7618 CSoutput.n246 CSoutput.n213 2.2505
R7619 CSoutput.n213 CSoutput.n207 2.2505
R7620 CSoutput.n268 CSoutput.n213 2.2505
R7621 CSoutput.n266 CSoutput.n213 2.2505
R7622 CSoutput.n248 CSoutput.n213 2.2505
R7623 CSoutput.n220 CSoutput.n213 2.2505
R7624 CSoutput.n250 CSoutput.n213 2.2505
R7625 CSoutput.n219 CSoutput.n213 2.2505
R7626 CSoutput.n264 CSoutput.n213 2.2505
R7627 CSoutput.n264 CSoutput.n217 2.2505
R7628 CSoutput.n164 CSoutput.n144 2.2505
R7629 CSoutput.n159 CSoutput.n144 2.2505
R7630 CSoutput.n157 CSoutput.n144 2.2505
R7631 CSoutput.n156 CSoutput.n144 2.2505
R7632 CSoutput.n285 CSoutput.n144 2.2505
R7633 CSoutput.n283 CSoutput.n144 2.2505
R7634 CSoutput.n281 CSoutput.n144 2.2505
R7635 CSoutput.n167 CSoutput.n144 2.2505
R7636 CSoutput.n166 CSoutput.n144 2.2505
R7637 CSoutput.n170 CSoutput.n144 2.2505
R7638 CSoutput.n169 CSoutput.n144 2.2505
R7639 CSoutput.n152 CSoutput.n144 2.2505
R7640 CSoutput.n288 CSoutput.n144 2.2505
R7641 CSoutput.n288 CSoutput.n287 2.2505
R7642 CSoutput.n206 CSoutput.n199 2.25024
R7643 CSoutput.n206 CSoutput.n192 2.25024
R7644 CSoutput.n274 CSoutput.n206 2.25024
R7645 CSoutput.n206 CSoutput.n202 2.25024
R7646 CSoutput.n206 CSoutput.n205 2.25024
R7647 CSoutput.n206 CSoutput.n173 2.25024
R7648 CSoutput.n256 CSoutput.n253 2.25024
R7649 CSoutput.n256 CSoutput.n252 2.25024
R7650 CSoutput.n256 CSoutput.n251 2.25024
R7651 CSoutput.n256 CSoutput.n218 2.25024
R7652 CSoutput.n256 CSoutput.n255 2.25024
R7653 CSoutput.n257 CSoutput.n256 2.25024
R7654 CSoutput.n172 CSoutput.n165 2.25024
R7655 CSoutput.n172 CSoutput.n158 2.25024
R7656 CSoutput.n284 CSoutput.n172 2.25024
R7657 CSoutput.n172 CSoutput.n168 2.25024
R7658 CSoutput.n172 CSoutput.n171 2.25024
R7659 CSoutput.n172 CSoutput.n139 2.25024
R7660 CSoutput.n273 CSoutput.n183 1.50111
R7661 CSoutput.n221 CSoutput.n207 1.50111
R7662 CSoutput.n283 CSoutput.n149 1.50111
R7663 CSoutput.n229 CSoutput.n228 1.501
R7664 CSoutput.n236 CSoutput.n235 1.501
R7665 CSoutput.n263 CSoutput.n262 1.501
R7666 CSoutput.n277 CSoutput.n188 1.12536
R7667 CSoutput.n277 CSoutput.n189 1.12536
R7668 CSoutput.n277 CSoutput.n276 1.12536
R7669 CSoutput.n237 CSoutput.n217 1.12536
R7670 CSoutput.n243 CSoutput.n217 1.12536
R7671 CSoutput.n245 CSoutput.n217 1.12536
R7672 CSoutput.n287 CSoutput.n154 1.12536
R7673 CSoutput.n287 CSoutput.n155 1.12536
R7674 CSoutput.n287 CSoutput.n286 1.12536
R7675 CSoutput.n277 CSoutput.n184 1.12536
R7676 CSoutput.n277 CSoutput.n185 1.12536
R7677 CSoutput.n277 CSoutput.n187 1.12536
R7678 CSoutput.n267 CSoutput.n217 1.12536
R7679 CSoutput.n247 CSoutput.n217 1.12536
R7680 CSoutput.n249 CSoutput.n217 1.12536
R7681 CSoutput.n287 CSoutput.n150 1.12536
R7682 CSoutput.n287 CSoutput.n151 1.12536
R7683 CSoutput.n287 CSoutput.n153 1.12536
R7684 CSoutput.n31 CSoutput.n30 0.669944
R7685 CSoutput.n62 CSoutput.n61 0.669944
R7686 CSoutput.n368 CSoutput.n366 0.573776
R7687 CSoutput.n370 CSoutput.n368 0.573776
R7688 CSoutput.n372 CSoutput.n370 0.573776
R7689 CSoutput.n374 CSoutput.n372 0.573776
R7690 CSoutput.n376 CSoutput.n374 0.573776
R7691 CSoutput.n378 CSoutput.n376 0.573776
R7692 CSoutput.n353 CSoutput.n351 0.573776
R7693 CSoutput.n355 CSoutput.n353 0.573776
R7694 CSoutput.n357 CSoutput.n355 0.573776
R7695 CSoutput.n359 CSoutput.n357 0.573776
R7696 CSoutput.n361 CSoutput.n359 0.573776
R7697 CSoutput.n363 CSoutput.n361 0.573776
R7698 CSoutput.n410 CSoutput.n408 0.573776
R7699 CSoutput.n408 CSoutput.n406 0.573776
R7700 CSoutput.n406 CSoutput.n404 0.573776
R7701 CSoutput.n404 CSoutput.n402 0.573776
R7702 CSoutput.n402 CSoutput.n400 0.573776
R7703 CSoutput.n400 CSoutput.n398 0.573776
R7704 CSoutput.n395 CSoutput.n393 0.573776
R7705 CSoutput.n393 CSoutput.n391 0.573776
R7706 CSoutput.n391 CSoutput.n389 0.573776
R7707 CSoutput.n389 CSoutput.n387 0.573776
R7708 CSoutput.n387 CSoutput.n385 0.573776
R7709 CSoutput.n385 CSoutput.n383 0.573776
R7710 CSoutput.n413 CSoutput.n288 0.53442
R7711 CSoutput.n332 CSoutput.n330 0.358259
R7712 CSoutput.n334 CSoutput.n332 0.358259
R7713 CSoutput.n336 CSoutput.n334 0.358259
R7714 CSoutput.n338 CSoutput.n336 0.358259
R7715 CSoutput.n340 CSoutput.n338 0.358259
R7716 CSoutput.n342 CSoutput.n340 0.358259
R7717 CSoutput.n344 CSoutput.n342 0.358259
R7718 CSoutput.n346 CSoutput.n344 0.358259
R7719 CSoutput.n312 CSoutput.n310 0.358259
R7720 CSoutput.n314 CSoutput.n312 0.358259
R7721 CSoutput.n316 CSoutput.n314 0.358259
R7722 CSoutput.n318 CSoutput.n316 0.358259
R7723 CSoutput.n320 CSoutput.n318 0.358259
R7724 CSoutput.n322 CSoutput.n320 0.358259
R7725 CSoutput.n324 CSoutput.n322 0.358259
R7726 CSoutput.n326 CSoutput.n324 0.358259
R7727 CSoutput.n293 CSoutput.n291 0.358259
R7728 CSoutput.n295 CSoutput.n293 0.358259
R7729 CSoutput.n297 CSoutput.n295 0.358259
R7730 CSoutput.n299 CSoutput.n297 0.358259
R7731 CSoutput.n301 CSoutput.n299 0.358259
R7732 CSoutput.n303 CSoutput.n301 0.358259
R7733 CSoutput.n305 CSoutput.n303 0.358259
R7734 CSoutput.n307 CSoutput.n305 0.358259
R7735 CSoutput.n136 CSoutput.n134 0.358259
R7736 CSoutput.n134 CSoutput.n132 0.358259
R7737 CSoutput.n132 CSoutput.n130 0.358259
R7738 CSoutput.n130 CSoutput.n128 0.358259
R7739 CSoutput.n128 CSoutput.n126 0.358259
R7740 CSoutput.n126 CSoutput.n124 0.358259
R7741 CSoutput.n124 CSoutput.n122 0.358259
R7742 CSoutput.n122 CSoutput.n120 0.358259
R7743 CSoutput.n116 CSoutput.n114 0.358259
R7744 CSoutput.n114 CSoutput.n112 0.358259
R7745 CSoutput.n112 CSoutput.n110 0.358259
R7746 CSoutput.n110 CSoutput.n108 0.358259
R7747 CSoutput.n108 CSoutput.n106 0.358259
R7748 CSoutput.n106 CSoutput.n104 0.358259
R7749 CSoutput.n104 CSoutput.n102 0.358259
R7750 CSoutput.n102 CSoutput.n100 0.358259
R7751 CSoutput.n97 CSoutput.n95 0.358259
R7752 CSoutput.n95 CSoutput.n93 0.358259
R7753 CSoutput.n93 CSoutput.n91 0.358259
R7754 CSoutput.n91 CSoutput.n89 0.358259
R7755 CSoutput.n89 CSoutput.n87 0.358259
R7756 CSoutput.n87 CSoutput.n85 0.358259
R7757 CSoutput.n85 CSoutput.n83 0.358259
R7758 CSoutput.n83 CSoutput.n81 0.358259
R7759 CSoutput.n21 CSoutput.n20 0.169105
R7760 CSoutput.n21 CSoutput.n16 0.169105
R7761 CSoutput.n26 CSoutput.n16 0.169105
R7762 CSoutput.n27 CSoutput.n26 0.169105
R7763 CSoutput.n27 CSoutput.n14 0.169105
R7764 CSoutput.n32 CSoutput.n14 0.169105
R7765 CSoutput.n33 CSoutput.n32 0.169105
R7766 CSoutput.n34 CSoutput.n33 0.169105
R7767 CSoutput.n34 CSoutput.n12 0.169105
R7768 CSoutput.n39 CSoutput.n12 0.169105
R7769 CSoutput.n40 CSoutput.n39 0.169105
R7770 CSoutput.n40 CSoutput.n10 0.169105
R7771 CSoutput.n45 CSoutput.n10 0.169105
R7772 CSoutput.n46 CSoutput.n45 0.169105
R7773 CSoutput.n47 CSoutput.n46 0.169105
R7774 CSoutput.n47 CSoutput.n8 0.169105
R7775 CSoutput.n52 CSoutput.n8 0.169105
R7776 CSoutput.n53 CSoutput.n52 0.169105
R7777 CSoutput.n53 CSoutput.n6 0.169105
R7778 CSoutput.n58 CSoutput.n6 0.169105
R7779 CSoutput.n59 CSoutput.n58 0.169105
R7780 CSoutput.n60 CSoutput.n59 0.169105
R7781 CSoutput.n60 CSoutput.n4 0.169105
R7782 CSoutput.n66 CSoutput.n4 0.169105
R7783 CSoutput.n67 CSoutput.n66 0.169105
R7784 CSoutput.n68 CSoutput.n67 0.169105
R7785 CSoutput.n68 CSoutput.n2 0.169105
R7786 CSoutput.n73 CSoutput.n2 0.169105
R7787 CSoutput.n74 CSoutput.n73 0.169105
R7788 CSoutput.n74 CSoutput.n0 0.169105
R7789 CSoutput.n78 CSoutput.n0 0.169105
R7790 CSoutput.n231 CSoutput.n230 0.0910737
R7791 CSoutput.n282 CSoutput.n279 0.0723685
R7792 CSoutput.n236 CSoutput.n231 0.0522944
R7793 CSoutput.n279 CSoutput.n278 0.0499135
R7794 CSoutput.n230 CSoutput.n229 0.0499135
R7795 CSoutput.n264 CSoutput.n263 0.0464294
R7796 CSoutput.n272 CSoutput.n269 0.0391444
R7797 CSoutput.n231 CSoutput.t202 0.023435
R7798 CSoutput.n279 CSoutput.t196 0.02262
R7799 CSoutput.n230 CSoutput.t187 0.02262
R7800 CSoutput CSoutput.n413 0.0052
R7801 CSoutput.n201 CSoutput.n184 0.00365111
R7802 CSoutput.n204 CSoutput.n185 0.00365111
R7803 CSoutput.n187 CSoutput.n186 0.00365111
R7804 CSoutput.n229 CSoutput.n188 0.00365111
R7805 CSoutput.n193 CSoutput.n189 0.00365111
R7806 CSoutput.n276 CSoutput.n190 0.00365111
R7807 CSoutput.n267 CSoutput.n266 0.00365111
R7808 CSoutput.n247 CSoutput.n220 0.00365111
R7809 CSoutput.n249 CSoutput.n219 0.00365111
R7810 CSoutput.n237 CSoutput.n236 0.00365111
R7811 CSoutput.n243 CSoutput.n223 0.00365111
R7812 CSoutput.n245 CSoutput.n222 0.00365111
R7813 CSoutput.n167 CSoutput.n150 0.00365111
R7814 CSoutput.n170 CSoutput.n151 0.00365111
R7815 CSoutput.n153 CSoutput.n152 0.00365111
R7816 CSoutput.n263 CSoutput.n154 0.00365111
R7817 CSoutput.n159 CSoutput.n155 0.00365111
R7818 CSoutput.n286 CSoutput.n156 0.00365111
R7819 CSoutput.n198 CSoutput.n188 0.00340054
R7820 CSoutput.n191 CSoutput.n189 0.00340054
R7821 CSoutput.n276 CSoutput.n275 0.00340054
R7822 CSoutput.n271 CSoutput.n184 0.00340054
R7823 CSoutput.n200 CSoutput.n185 0.00340054
R7824 CSoutput.n203 CSoutput.n187 0.00340054
R7825 CSoutput.n242 CSoutput.n237 0.00340054
R7826 CSoutput.n244 CSoutput.n243 0.00340054
R7827 CSoutput.n246 CSoutput.n245 0.00340054
R7828 CSoutput.n268 CSoutput.n267 0.00340054
R7829 CSoutput.n248 CSoutput.n247 0.00340054
R7830 CSoutput.n250 CSoutput.n249 0.00340054
R7831 CSoutput.n164 CSoutput.n154 0.00340054
R7832 CSoutput.n157 CSoutput.n155 0.00340054
R7833 CSoutput.n286 CSoutput.n285 0.00340054
R7834 CSoutput.n281 CSoutput.n150 0.00340054
R7835 CSoutput.n166 CSoutput.n151 0.00340054
R7836 CSoutput.n169 CSoutput.n153 0.00340054
R7837 CSoutput.n199 CSoutput.n193 0.00252698
R7838 CSoutput.n192 CSoutput.n190 0.00252698
R7839 CSoutput.n274 CSoutput.n273 0.00252698
R7840 CSoutput.n202 CSoutput.n200 0.00252698
R7841 CSoutput.n205 CSoutput.n203 0.00252698
R7842 CSoutput.n278 CSoutput.n173 0.00252698
R7843 CSoutput.n199 CSoutput.n198 0.00252698
R7844 CSoutput.n192 CSoutput.n191 0.00252698
R7845 CSoutput.n275 CSoutput.n274 0.00252698
R7846 CSoutput.n202 CSoutput.n201 0.00252698
R7847 CSoutput.n205 CSoutput.n204 0.00252698
R7848 CSoutput.n186 CSoutput.n173 0.00252698
R7849 CSoutput.n253 CSoutput.n223 0.00252698
R7850 CSoutput.n252 CSoutput.n222 0.00252698
R7851 CSoutput.n251 CSoutput.n207 0.00252698
R7852 CSoutput.n248 CSoutput.n218 0.00252698
R7853 CSoutput.n255 CSoutput.n250 0.00252698
R7854 CSoutput.n264 CSoutput.n257 0.00252698
R7855 CSoutput.n253 CSoutput.n242 0.00252698
R7856 CSoutput.n252 CSoutput.n244 0.00252698
R7857 CSoutput.n251 CSoutput.n246 0.00252698
R7858 CSoutput.n266 CSoutput.n218 0.00252698
R7859 CSoutput.n255 CSoutput.n220 0.00252698
R7860 CSoutput.n257 CSoutput.n219 0.00252698
R7861 CSoutput.n165 CSoutput.n159 0.00252698
R7862 CSoutput.n158 CSoutput.n156 0.00252698
R7863 CSoutput.n284 CSoutput.n283 0.00252698
R7864 CSoutput.n168 CSoutput.n166 0.00252698
R7865 CSoutput.n171 CSoutput.n169 0.00252698
R7866 CSoutput.n288 CSoutput.n139 0.00252698
R7867 CSoutput.n165 CSoutput.n164 0.00252698
R7868 CSoutput.n158 CSoutput.n157 0.00252698
R7869 CSoutput.n285 CSoutput.n284 0.00252698
R7870 CSoutput.n168 CSoutput.n167 0.00252698
R7871 CSoutput.n171 CSoutput.n170 0.00252698
R7872 CSoutput.n152 CSoutput.n139 0.00252698
R7873 CSoutput.n273 CSoutput.n272 0.0020275
R7874 CSoutput.n272 CSoutput.n271 0.0020275
R7875 CSoutput.n269 CSoutput.n207 0.0020275
R7876 CSoutput.n269 CSoutput.n268 0.0020275
R7877 CSoutput.n283 CSoutput.n282 0.0020275
R7878 CSoutput.n282 CSoutput.n281 0.0020275
R7879 CSoutput.n183 CSoutput.n182 0.00166668
R7880 CSoutput.n265 CSoutput.n221 0.00166668
R7881 CSoutput.n149 CSoutput.n148 0.00166668
R7882 CSoutput.n287 CSoutput.n149 0.00133328
R7883 CSoutput.n221 CSoutput.n217 0.00133328
R7884 CSoutput.n277 CSoutput.n183 0.00133328
R7885 CSoutput.n280 CSoutput.n172 0.001
R7886 CSoutput.n258 CSoutput.n172 0.001
R7887 CSoutput.n160 CSoutput.n140 0.001
R7888 CSoutput.n259 CSoutput.n140 0.001
R7889 CSoutput.n161 CSoutput.n141 0.001
R7890 CSoutput.n260 CSoutput.n141 0.001
R7891 CSoutput.n162 CSoutput.n142 0.001
R7892 CSoutput.n261 CSoutput.n142 0.001
R7893 CSoutput.n163 CSoutput.n143 0.001
R7894 CSoutput.n262 CSoutput.n143 0.001
R7895 CSoutput.n256 CSoutput.n208 0.001
R7896 CSoutput.n256 CSoutput.n254 0.001
R7897 CSoutput.n238 CSoutput.n209 0.001
R7898 CSoutput.n232 CSoutput.n209 0.001
R7899 CSoutput.n239 CSoutput.n210 0.001
R7900 CSoutput.n233 CSoutput.n210 0.001
R7901 CSoutput.n240 CSoutput.n211 0.001
R7902 CSoutput.n234 CSoutput.n211 0.001
R7903 CSoutput.n241 CSoutput.n212 0.001
R7904 CSoutput.n235 CSoutput.n212 0.001
R7905 CSoutput.n270 CSoutput.n206 0.001
R7906 CSoutput.n224 CSoutput.n206 0.001
R7907 CSoutput.n194 CSoutput.n174 0.001
R7908 CSoutput.n225 CSoutput.n174 0.001
R7909 CSoutput.n195 CSoutput.n175 0.001
R7910 CSoutput.n226 CSoutput.n175 0.001
R7911 CSoutput.n196 CSoutput.n176 0.001
R7912 CSoutput.n227 CSoutput.n176 0.001
R7913 CSoutput.n197 CSoutput.n177 0.001
R7914 CSoutput.n228 CSoutput.n177 0.001
R7915 CSoutput.n228 CSoutput.n178 0.001
R7916 CSoutput.n227 CSoutput.n179 0.001
R7917 CSoutput.n226 CSoutput.n180 0.001
R7918 CSoutput.n225 CSoutput.t199 0.001
R7919 CSoutput.n224 CSoutput.n181 0.001
R7920 CSoutput.n197 CSoutput.n179 0.001
R7921 CSoutput.n196 CSoutput.n180 0.001
R7922 CSoutput.n195 CSoutput.t199 0.001
R7923 CSoutput.n194 CSoutput.n181 0.001
R7924 CSoutput.n270 CSoutput.n182 0.001
R7925 CSoutput.n235 CSoutput.n213 0.001
R7926 CSoutput.n234 CSoutput.n214 0.001
R7927 CSoutput.n233 CSoutput.n215 0.001
R7928 CSoutput.n232 CSoutput.t195 0.001
R7929 CSoutput.n254 CSoutput.n216 0.001
R7930 CSoutput.n241 CSoutput.n214 0.001
R7931 CSoutput.n240 CSoutput.n215 0.001
R7932 CSoutput.n239 CSoutput.t195 0.001
R7933 CSoutput.n238 CSoutput.n216 0.001
R7934 CSoutput.n265 CSoutput.n208 0.001
R7935 CSoutput.n262 CSoutput.n144 0.001
R7936 CSoutput.n261 CSoutput.n145 0.001
R7937 CSoutput.n260 CSoutput.n146 0.001
R7938 CSoutput.n259 CSoutput.t185 0.001
R7939 CSoutput.n258 CSoutput.n147 0.001
R7940 CSoutput.n163 CSoutput.n145 0.001
R7941 CSoutput.n162 CSoutput.n146 0.001
R7942 CSoutput.n161 CSoutput.t185 0.001
R7943 CSoutput.n160 CSoutput.n147 0.001
R7944 CSoutput.n280 CSoutput.n148 0.001
R7945 a_n2650_13878.n114 a_n2650_13878.t80 512.366
R7946 a_n2650_13878.n113 a_n2650_13878.t70 512.366
R7947 a_n2650_13878.n112 a_n2650_13878.t60 512.366
R7948 a_n2650_13878.n116 a_n2650_13878.t88 512.366
R7949 a_n2650_13878.n115 a_n2650_13878.t77 512.366
R7950 a_n2650_13878.n111 a_n2650_13878.t76 512.366
R7951 a_n2650_13878.n118 a_n2650_13878.t84 512.366
R7952 a_n2650_13878.n117 a_n2650_13878.t68 512.366
R7953 a_n2650_13878.n110 a_n2650_13878.t69 512.366
R7954 a_n2650_13878.n120 a_n2650_13878.t71 512.366
R7955 a_n2650_13878.n119 a_n2650_13878.t81 512.366
R7956 a_n2650_13878.n109 a_n2650_13878.t95 512.366
R7957 a_n2650_13878.n96 a_n2650_13878.t94 512.366
R7958 a_n2650_13878.n95 a_n2650_13878.t73 512.366
R7959 a_n2650_13878.n88 a_n2650_13878.t78 512.366
R7960 a_n2650_13878.n94 a_n2650_13878.t67 512.366
R7961 a_n2650_13878.n93 a_n2650_13878.t83 512.366
R7962 a_n2650_13878.n89 a_n2650_13878.t91 512.366
R7963 a_n2650_13878.n92 a_n2650_13878.t92 512.366
R7964 a_n2650_13878.n91 a_n2650_13878.t62 512.366
R7965 a_n2650_13878.n90 a_n2650_13878.t75 512.366
R7966 a_n2650_13878.n102 a_n2650_13878.t11 512.366
R7967 a_n2650_13878.n101 a_n2650_13878.t17 512.366
R7968 a_n2650_13878.n75 a_n2650_13878.t45 512.366
R7969 a_n2650_13878.n100 a_n2650_13878.t31 512.366
R7970 a_n2650_13878.n99 a_n2650_13878.t39 512.366
R7971 a_n2650_13878.n76 a_n2650_13878.t33 512.366
R7972 a_n2650_13878.n98 a_n2650_13878.t13 512.366
R7973 a_n2650_13878.n97 a_n2650_13878.t37 512.366
R7974 a_n2650_13878.n77 a_n2650_13878.t23 512.366
R7975 a_n2650_13878.n129 a_n2650_13878.t29 512.366
R7976 a_n2650_13878.n130 a_n2650_13878.t43 512.366
R7977 a_n2650_13878.n72 a_n2650_13878.t47 512.366
R7978 a_n2650_13878.n131 a_n2650_13878.t35 512.366
R7979 a_n2650_13878.n132 a_n2650_13878.t9 512.366
R7980 a_n2650_13878.n133 a_n2650_13878.t27 512.366
R7981 a_n2650_13878.n134 a_n2650_13878.t15 512.366
R7982 a_n2650_13878.n71 a_n2650_13878.t21 512.366
R7983 a_n2650_13878.n135 a_n2650_13878.t41 512.366
R7984 a_n2650_13878.n122 a_n2650_13878.t66 512.366
R7985 a_n2650_13878.n123 a_n2650_13878.t89 512.366
R7986 a_n2650_13878.n74 a_n2650_13878.t90 512.366
R7987 a_n2650_13878.n124 a_n2650_13878.t64 512.366
R7988 a_n2650_13878.n125 a_n2650_13878.t86 512.366
R7989 a_n2650_13878.n126 a_n2650_13878.t87 512.366
R7990 a_n2650_13878.n127 a_n2650_13878.t61 512.366
R7991 a_n2650_13878.n73 a_n2650_13878.t72 512.366
R7992 a_n2650_13878.n128 a_n2650_13878.t82 512.366
R7993 a_n2650_13878.n4 a_n2650_13878.n68 70.1674
R7994 a_n2650_13878.n6 a_n2650_13878.n66 70.1674
R7995 a_n2650_13878.n8 a_n2650_13878.n64 70.1674
R7996 a_n2650_13878.n10 a_n2650_13878.n62 70.1674
R7997 a_n2650_13878.n24 a_n2650_13878.n41 70.1674
R7998 a_n2650_13878.n32 a_n2650_13878.n33 70.1674
R7999 a_n2650_13878.n33 a_n2650_13878.n77 20.9683
R8000 a_n2650_13878.n69 a_n2650_13878.n21 74.73
R8001 a_n2650_13878.n41 a_n2650_13878.n90 20.9683
R8002 a_n2650_13878.n39 a_n2650_13878.n24 74.73
R8003 a_n2650_13878.n91 a_n2650_13878.n39 11.843
R8004 a_n2650_13878.n38 a_n2650_13878.n23 80.4688
R8005 a_n2650_13878.n38 a_n2650_13878.n92 0.365327
R8006 a_n2650_13878.n23 a_n2650_13878.n37 75.0448
R8007 a_n2650_13878.n36 a_n2650_13878.n25 70.1674
R8008 a_n2650_13878.n94 a_n2650_13878.n36 20.9683
R8009 a_n2650_13878.n25 a_n2650_13878.n35 70.3058
R8010 a_n2650_13878.n35 a_n2650_13878.n88 20.6913
R8011 a_n2650_13878.n34 a_n2650_13878.n26 75.3623
R8012 a_n2650_13878.n95 a_n2650_13878.n34 10.5784
R8013 a_n2650_13878.n26 a_n2650_13878.n96 161.3
R8014 a_n2650_13878.n97 a_n2650_13878.n69 11.843
R8015 a_n2650_13878.n46 a_n2650_13878.n21 80.4688
R8016 a_n2650_13878.n46 a_n2650_13878.n98 0.365327
R8017 a_n2650_13878.n21 a_n2650_13878.n45 75.0448
R8018 a_n2650_13878.n44 a_n2650_13878.n20 70.1674
R8019 a_n2650_13878.n100 a_n2650_13878.n44 20.9683
R8020 a_n2650_13878.n20 a_n2650_13878.n43 70.3058
R8021 a_n2650_13878.n43 a_n2650_13878.n75 20.6913
R8022 a_n2650_13878.n42 a_n2650_13878.n22 75.3623
R8023 a_n2650_13878.n101 a_n2650_13878.n42 10.5784
R8024 a_n2650_13878.n22 a_n2650_13878.n102 161.3
R8025 a_n2650_13878.n13 a_n2650_13878.n60 70.1674
R8026 a_n2650_13878.n17 a_n2650_13878.n53 70.1674
R8027 a_n2650_13878.n128 a_n2650_13878.n53 20.9683
R8028 a_n2650_13878.n52 a_n2650_13878.n17 74.73
R8029 a_n2650_13878.n52 a_n2650_13878.n73 11.843
R8030 a_n2650_13878.n16 a_n2650_13878.n51 80.4688
R8031 a_n2650_13878.n127 a_n2650_13878.n51 0.365327
R8032 a_n2650_13878.n50 a_n2650_13878.n16 75.0448
R8033 a_n2650_13878.n18 a_n2650_13878.n49 70.1674
R8034 a_n2650_13878.n124 a_n2650_13878.n49 20.9683
R8035 a_n2650_13878.n48 a_n2650_13878.n18 70.3058
R8036 a_n2650_13878.n48 a_n2650_13878.n74 20.6913
R8037 a_n2650_13878.n19 a_n2650_13878.n47 75.3623
R8038 a_n2650_13878.n123 a_n2650_13878.n47 10.5784
R8039 a_n2650_13878.n122 a_n2650_13878.n19 161.3
R8040 a_n2650_13878.n135 a_n2650_13878.n60 20.9683
R8041 a_n2650_13878.n59 a_n2650_13878.n13 74.73
R8042 a_n2650_13878.n59 a_n2650_13878.n71 11.843
R8043 a_n2650_13878.n12 a_n2650_13878.n58 80.4688
R8044 a_n2650_13878.n134 a_n2650_13878.n58 0.365327
R8045 a_n2650_13878.n57 a_n2650_13878.n12 75.0448
R8046 a_n2650_13878.n14 a_n2650_13878.n56 70.1674
R8047 a_n2650_13878.n131 a_n2650_13878.n56 20.9683
R8048 a_n2650_13878.n55 a_n2650_13878.n14 70.3058
R8049 a_n2650_13878.n55 a_n2650_13878.n72 20.6913
R8050 a_n2650_13878.n15 a_n2650_13878.n54 75.3623
R8051 a_n2650_13878.n130 a_n2650_13878.n54 10.5784
R8052 a_n2650_13878.n129 a_n2650_13878.n15 161.3
R8053 a_n2650_13878.n62 a_n2650_13878.n109 20.9683
R8054 a_n2650_13878.n61 a_n2650_13878.n11 75.0448
R8055 a_n2650_13878.n119 a_n2650_13878.n61 11.2134
R8056 a_n2650_13878.n11 a_n2650_13878.n120 161.3
R8057 a_n2650_13878.n64 a_n2650_13878.n110 20.9683
R8058 a_n2650_13878.n63 a_n2650_13878.n9 75.0448
R8059 a_n2650_13878.n117 a_n2650_13878.n63 11.2134
R8060 a_n2650_13878.n9 a_n2650_13878.n118 161.3
R8061 a_n2650_13878.n66 a_n2650_13878.n111 20.9683
R8062 a_n2650_13878.n65 a_n2650_13878.n7 75.0448
R8063 a_n2650_13878.n115 a_n2650_13878.n65 11.2134
R8064 a_n2650_13878.n7 a_n2650_13878.n116 161.3
R8065 a_n2650_13878.n68 a_n2650_13878.n112 20.9683
R8066 a_n2650_13878.n67 a_n2650_13878.n5 75.0448
R8067 a_n2650_13878.n113 a_n2650_13878.n67 11.2134
R8068 a_n2650_13878.n5 a_n2650_13878.n114 161.3
R8069 a_n2650_13878.n3 a_n2650_13878.n86 81.4626
R8070 a_n2650_13878.n1 a_n2650_13878.n81 81.4626
R8071 a_n2650_13878.n0 a_n2650_13878.n78 81.4626
R8072 a_n2650_13878.n3 a_n2650_13878.n87 80.9324
R8073 a_n2650_13878.n3 a_n2650_13878.n85 80.9324
R8074 a_n2650_13878.n2 a_n2650_13878.n84 80.9324
R8075 a_n2650_13878.n2 a_n2650_13878.n83 80.9324
R8076 a_n2650_13878.n1 a_n2650_13878.n82 80.9324
R8077 a_n2650_13878.n1 a_n2650_13878.n80 80.9324
R8078 a_n2650_13878.n0 a_n2650_13878.n79 80.9324
R8079 a_n2650_13878.n30 a_n2650_13878.t30 74.6477
R8080 a_n2650_13878.n27 a_n2650_13878.t26 74.6477
R8081 a_n2650_13878.n107 a_n2650_13878.t12 74.2899
R8082 a_n2650_13878.n29 a_n2650_13878.t20 74.2897
R8083 a_n2650_13878.n29 a_n2650_13878.n137 70.6783
R8084 a_n2650_13878.n31 a_n2650_13878.n138 70.6783
R8085 a_n2650_13878.n30 a_n2650_13878.n70 70.6783
R8086 a_n2650_13878.n27 a_n2650_13878.n103 70.6783
R8087 a_n2650_13878.n27 a_n2650_13878.n104 70.6783
R8088 a_n2650_13878.n28 a_n2650_13878.n105 70.6783
R8089 a_n2650_13878.n28 a_n2650_13878.n106 70.6783
R8090 a_n2650_13878.n139 a_n2650_13878.n31 70.6782
R8091 a_n2650_13878.n114 a_n2650_13878.n113 48.2005
R8092 a_n2650_13878.t85 a_n2650_13878.n68 533.335
R8093 a_n2650_13878.n116 a_n2650_13878.n115 48.2005
R8094 a_n2650_13878.t93 a_n2650_13878.n66 533.335
R8095 a_n2650_13878.n118 a_n2650_13878.n117 48.2005
R8096 a_n2650_13878.t79 a_n2650_13878.n64 533.335
R8097 a_n2650_13878.n120 a_n2650_13878.n119 48.2005
R8098 a_n2650_13878.t74 a_n2650_13878.n62 533.335
R8099 a_n2650_13878.n96 a_n2650_13878.n95 48.2005
R8100 a_n2650_13878.n36 a_n2650_13878.n93 20.9683
R8101 a_n2650_13878.n92 a_n2650_13878.n89 48.2005
R8102 a_n2650_13878.t65 a_n2650_13878.n41 533.335
R8103 a_n2650_13878.n102 a_n2650_13878.n101 48.2005
R8104 a_n2650_13878.n44 a_n2650_13878.n99 20.9683
R8105 a_n2650_13878.n98 a_n2650_13878.n76 48.2005
R8106 a_n2650_13878.t25 a_n2650_13878.n33 533.335
R8107 a_n2650_13878.n130 a_n2650_13878.n129 48.2005
R8108 a_n2650_13878.n132 a_n2650_13878.n56 20.9683
R8109 a_n2650_13878.n134 a_n2650_13878.n133 48.2005
R8110 a_n2650_13878.t19 a_n2650_13878.n60 533.335
R8111 a_n2650_13878.n123 a_n2650_13878.n122 48.2005
R8112 a_n2650_13878.n125 a_n2650_13878.n49 20.9683
R8113 a_n2650_13878.n127 a_n2650_13878.n126 48.2005
R8114 a_n2650_13878.t63 a_n2650_13878.n53 533.335
R8115 a_n2650_13878.n94 a_n2650_13878.n35 21.4216
R8116 a_n2650_13878.n100 a_n2650_13878.n43 21.4216
R8117 a_n2650_13878.n131 a_n2650_13878.n55 21.4216
R8118 a_n2650_13878.n124 a_n2650_13878.n48 21.4216
R8119 a_n2650_13878.n2 a_n2650_13878.n1 32.7898
R8120 a_n2650_13878.n39 a_n2650_13878.n90 34.4824
R8121 a_n2650_13878.n69 a_n2650_13878.n77 34.4824
R8122 a_n2650_13878.n135 a_n2650_13878.n59 34.4824
R8123 a_n2650_13878.n128 a_n2650_13878.n52 34.4824
R8124 a_n2650_13878.n67 a_n2650_13878.n112 35.3134
R8125 a_n2650_13878.n65 a_n2650_13878.n111 35.3134
R8126 a_n2650_13878.n63 a_n2650_13878.n110 35.3134
R8127 a_n2650_13878.n61 a_n2650_13878.n109 35.3134
R8128 a_n2650_13878.n93 a_n2650_13878.n37 35.3134
R8129 a_n2650_13878.n37 a_n2650_13878.n89 11.2134
R8130 a_n2650_13878.n99 a_n2650_13878.n45 35.3134
R8131 a_n2650_13878.n45 a_n2650_13878.n76 11.2134
R8132 a_n2650_13878.n132 a_n2650_13878.n57 35.3134
R8133 a_n2650_13878.n133 a_n2650_13878.n57 11.2134
R8134 a_n2650_13878.n125 a_n2650_13878.n50 35.3134
R8135 a_n2650_13878.n126 a_n2650_13878.n50 11.2134
R8136 a_n2650_13878.n21 a_n2650_13878.n3 23.891
R8137 a_n2650_13878.n34 a_n2650_13878.n88 36.139
R8138 a_n2650_13878.n42 a_n2650_13878.n75 36.139
R8139 a_n2650_13878.n72 a_n2650_13878.n54 36.139
R8140 a_n2650_13878.n74 a_n2650_13878.n47 36.139
R8141 a_n2650_13878.n19 a_n2650_13878.n121 13.3641
R8142 a_n2650_13878.n24 a_n2650_13878.n40 13.1596
R8143 a_n2650_13878.n108 a_n2650_13878.n22 11.8547
R8144 a_n2650_13878.n29 a_n2650_13878.n136 10.2167
R8145 a_n2650_13878.n121 a_n2650_13878.n11 9.99103
R8146 a_n2650_13878.n4 a_n2650_13878.n40 9.99103
R8147 a_n2650_13878.n136 a_n2650_13878.n13 8.01944
R8148 a_n2650_13878.n108 a_n2650_13878.n107 6.37334
R8149 a_n2650_13878.n136 a_n2650_13878.n40 5.3452
R8150 a_n2650_13878.n32 a_n2650_13878.n26 4.07247
R8151 a_n2650_13878.n15 a_n2650_13878.n17 4.07247
R8152 a_n2650_13878.n137 a_n2650_13878.t22 3.61217
R8153 a_n2650_13878.n137 a_n2650_13878.t42 3.61217
R8154 a_n2650_13878.n138 a_n2650_13878.t28 3.61217
R8155 a_n2650_13878.n138 a_n2650_13878.t16 3.61217
R8156 a_n2650_13878.n70 a_n2650_13878.t44 3.61217
R8157 a_n2650_13878.n70 a_n2650_13878.t48 3.61217
R8158 a_n2650_13878.n103 a_n2650_13878.t38 3.61217
R8159 a_n2650_13878.n103 a_n2650_13878.t24 3.61217
R8160 a_n2650_13878.n104 a_n2650_13878.t34 3.61217
R8161 a_n2650_13878.n104 a_n2650_13878.t14 3.61217
R8162 a_n2650_13878.n105 a_n2650_13878.t32 3.61217
R8163 a_n2650_13878.n105 a_n2650_13878.t40 3.61217
R8164 a_n2650_13878.n106 a_n2650_13878.t18 3.61217
R8165 a_n2650_13878.n106 a_n2650_13878.t46 3.61217
R8166 a_n2650_13878.n139 a_n2650_13878.t36 3.61217
R8167 a_n2650_13878.t10 a_n2650_13878.n139 3.61217
R8168 a_n2650_13878.n86 a_n2650_13878.t5 2.82907
R8169 a_n2650_13878.n86 a_n2650_13878.t2 2.82907
R8170 a_n2650_13878.n87 a_n2650_13878.t51 2.82907
R8171 a_n2650_13878.n87 a_n2650_13878.t6 2.82907
R8172 a_n2650_13878.n85 a_n2650_13878.t4 2.82907
R8173 a_n2650_13878.n85 a_n2650_13878.t0 2.82907
R8174 a_n2650_13878.n84 a_n2650_13878.t58 2.82907
R8175 a_n2650_13878.n84 a_n2650_13878.t1 2.82907
R8176 a_n2650_13878.n83 a_n2650_13878.t55 2.82907
R8177 a_n2650_13878.n83 a_n2650_13878.t59 2.82907
R8178 a_n2650_13878.n81 a_n2650_13878.t50 2.82907
R8179 a_n2650_13878.n81 a_n2650_13878.t54 2.82907
R8180 a_n2650_13878.n82 a_n2650_13878.t56 2.82907
R8181 a_n2650_13878.n82 a_n2650_13878.t53 2.82907
R8182 a_n2650_13878.n80 a_n2650_13878.t52 2.82907
R8183 a_n2650_13878.n80 a_n2650_13878.t3 2.82907
R8184 a_n2650_13878.n79 a_n2650_13878.t7 2.82907
R8185 a_n2650_13878.n79 a_n2650_13878.t49 2.82907
R8186 a_n2650_13878.n78 a_n2650_13878.t8 2.82907
R8187 a_n2650_13878.n78 a_n2650_13878.t57 2.82907
R8188 a_n2650_13878.n121 a_n2650_13878.n108 1.30542
R8189 a_n2650_13878.n8 a_n2650_13878.n7 1.04595
R8190 a_n2650_13878.n38 a_n2650_13878.n91 47.835
R8191 a_n2650_13878.n46 a_n2650_13878.n97 47.835
R8192 a_n2650_13878.n71 a_n2650_13878.n58 47.835
R8193 a_n2650_13878.n73 a_n2650_13878.n51 47.835
R8194 a_n2650_13878.n3 a_n2650_13878.n2 1.59102
R8195 a_n2650_13878.n24 a_n2650_13878.n23 1.13686
R8196 a_n2650_13878.n17 a_n2650_13878.n16 1.13686
R8197 a_n2650_13878.n13 a_n2650_13878.n12 1.13686
R8198 a_n2650_13878.n21 a_n2650_13878.n32 1.09898
R8199 a_n2650_13878.n1 a_n2650_13878.n0 1.06084
R8200 a_n2650_13878.n26 a_n2650_13878.n25 0.758076
R8201 a_n2650_13878.n23 a_n2650_13878.n25 0.758076
R8202 a_n2650_13878.n22 a_n2650_13878.n20 0.758076
R8203 a_n2650_13878.n21 a_n2650_13878.n20 0.758076
R8204 a_n2650_13878.n18 a_n2650_13878.n19 0.758076
R8205 a_n2650_13878.n16 a_n2650_13878.n18 0.758076
R8206 a_n2650_13878.n14 a_n2650_13878.n15 0.758076
R8207 a_n2650_13878.n12 a_n2650_13878.n14 0.758076
R8208 a_n2650_13878.n11 a_n2650_13878.n10 0.758076
R8209 a_n2650_13878.n9 a_n2650_13878.n8 0.758076
R8210 a_n2650_13878.n7 a_n2650_13878.n6 0.758076
R8211 a_n2650_13878.n5 a_n2650_13878.n4 0.758076
R8212 a_n2650_13878.n31 a_n2650_13878.n29 0.716017
R8213 a_n2650_13878.n31 a_n2650_13878.n30 0.716017
R8214 a_n2650_13878.n28 a_n2650_13878.n27 0.716017
R8215 a_n2650_13878.n107 a_n2650_13878.n28 0.716017
R8216 a_n2650_13878.n10 a_n2650_13878.n9 0.67853
R8217 a_n2650_13878.n6 a_n2650_13878.n5 0.67853
R8218 a_n2472_13878.n2 a_n2472_13878.n0 98.9633
R8219 a_n2472_13878.n5 a_n2472_13878.n3 98.7517
R8220 a_n2472_13878.n23 a_n2472_13878.n22 98.6055
R8221 a_n2472_13878.n2 a_n2472_13878.n1 98.6055
R8222 a_n2472_13878.n11 a_n2472_13878.n10 98.6055
R8223 a_n2472_13878.n9 a_n2472_13878.n8 98.6055
R8224 a_n2472_13878.n7 a_n2472_13878.n6 98.6055
R8225 a_n2472_13878.n5 a_n2472_13878.n4 98.6055
R8226 a_n2472_13878.n25 a_n2472_13878.n24 98.6054
R8227 a_n2472_13878.n21 a_n2472_13878.n20 98.6054
R8228 a_n2472_13878.n13 a_n2472_13878.t1 74.6477
R8229 a_n2472_13878.n18 a_n2472_13878.t2 74.2899
R8230 a_n2472_13878.n15 a_n2472_13878.t3 74.2899
R8231 a_n2472_13878.n14 a_n2472_13878.t0 74.2899
R8232 a_n2472_13878.n17 a_n2472_13878.n16 70.6783
R8233 a_n2472_13878.n13 a_n2472_13878.n12 70.6783
R8234 a_n2472_13878.n19 a_n2472_13878.n11 15.0004
R8235 a_n2472_13878.n21 a_n2472_13878.n19 12.2917
R8236 a_n2472_13878.n19 a_n2472_13878.n18 7.67184
R8237 a_n2472_13878.n20 a_n2472_13878.t24 3.61217
R8238 a_n2472_13878.n20 a_n2472_13878.t13 3.61217
R8239 a_n2472_13878.n22 a_n2472_13878.t16 3.61217
R8240 a_n2472_13878.n22 a_n2472_13878.t17 3.61217
R8241 a_n2472_13878.n1 a_n2472_13878.t8 3.61217
R8242 a_n2472_13878.n1 a_n2472_13878.t18 3.61217
R8243 a_n2472_13878.n0 a_n2472_13878.t21 3.61217
R8244 a_n2472_13878.n0 a_n2472_13878.t27 3.61217
R8245 a_n2472_13878.n16 a_n2472_13878.t6 3.61217
R8246 a_n2472_13878.n16 a_n2472_13878.t7 3.61217
R8247 a_n2472_13878.n12 a_n2472_13878.t4 3.61217
R8248 a_n2472_13878.n12 a_n2472_13878.t5 3.61217
R8249 a_n2472_13878.n10 a_n2472_13878.t19 3.61217
R8250 a_n2472_13878.n10 a_n2472_13878.t9 3.61217
R8251 a_n2472_13878.n8 a_n2472_13878.t22 3.61217
R8252 a_n2472_13878.n8 a_n2472_13878.t11 3.61217
R8253 a_n2472_13878.n6 a_n2472_13878.t10 3.61217
R8254 a_n2472_13878.n6 a_n2472_13878.t12 3.61217
R8255 a_n2472_13878.n4 a_n2472_13878.t20 3.61217
R8256 a_n2472_13878.n4 a_n2472_13878.t14 3.61217
R8257 a_n2472_13878.n3 a_n2472_13878.t23 3.61217
R8258 a_n2472_13878.n3 a_n2472_13878.t15 3.61217
R8259 a_n2472_13878.n25 a_n2472_13878.t25 3.61217
R8260 a_n2472_13878.t26 a_n2472_13878.n25 3.61217
R8261 a_n2472_13878.n14 a_n2472_13878.n13 0.358259
R8262 a_n2472_13878.n17 a_n2472_13878.n15 0.358259
R8263 a_n2472_13878.n18 a_n2472_13878.n17 0.358259
R8264 a_n2472_13878.n24 a_n2472_13878.n2 0.358259
R8265 a_n2472_13878.n24 a_n2472_13878.n23 0.358259
R8266 a_n2472_13878.n23 a_n2472_13878.n21 0.358259
R8267 a_n2472_13878.n7 a_n2472_13878.n5 0.146627
R8268 a_n2472_13878.n9 a_n2472_13878.n7 0.146627
R8269 a_n2472_13878.n11 a_n2472_13878.n9 0.146627
R8270 a_n2472_13878.n15 a_n2472_13878.n14 0.101793
R8271 plus.n61 plus.t11 251.488
R8272 plus.n12 plus.t14 251.488
R8273 plus.n100 plus.t1 243.97
R8274 plus.n96 plus.t23 231.093
R8275 plus.n47 plus.t6 231.093
R8276 plus.n100 plus.n99 223.454
R8277 plus.n102 plus.n101 223.454
R8278 plus.n60 plus.t5 187.445
R8279 plus.n65 plus.t21 187.445
R8280 plus.n71 plus.t20 187.445
R8281 plus.n56 plus.t16 187.445
R8282 plus.n54 plus.t17 187.445
R8283 plus.n83 plus.t13 187.445
R8284 plus.n89 plus.t15 187.445
R8285 plus.n50 plus.t10 187.445
R8286 plus.n1 plus.t12 187.445
R8287 plus.n40 plus.t8 187.445
R8288 plus.n34 plus.t7 187.445
R8289 plus.n5 plus.t19 187.445
R8290 plus.n7 plus.t18 187.445
R8291 plus.n22 plus.t24 187.445
R8292 plus.n16 plus.t22 187.445
R8293 plus.n11 plus.t9 187.445
R8294 plus.n97 plus.n96 161.3
R8295 plus.n95 plus.n49 161.3
R8296 plus.n94 plus.n93 161.3
R8297 plus.n92 plus.n91 161.3
R8298 plus.n90 plus.n51 161.3
R8299 plus.n88 plus.n87 161.3
R8300 plus.n86 plus.n52 161.3
R8301 plus.n85 plus.n84 161.3
R8302 plus.n82 plus.n53 161.3
R8303 plus.n81 plus.n80 161.3
R8304 plus.n79 plus.n78 161.3
R8305 plus.n77 plus.n55 161.3
R8306 plus.n76 plus.n75 161.3
R8307 plus.n74 plus.n73 161.3
R8308 plus.n72 plus.n57 161.3
R8309 plus.n70 plus.n69 161.3
R8310 plus.n68 plus.n58 161.3
R8311 plus.n67 plus.n66 161.3
R8312 plus.n64 plus.n59 161.3
R8313 plus.n63 plus.n62 161.3
R8314 plus.n14 plus.n13 161.3
R8315 plus.n15 plus.n10 161.3
R8316 plus.n18 plus.n17 161.3
R8317 plus.n19 plus.n9 161.3
R8318 plus.n21 plus.n20 161.3
R8319 plus.n23 plus.n8 161.3
R8320 plus.n25 plus.n24 161.3
R8321 plus.n27 plus.n26 161.3
R8322 plus.n28 plus.n6 161.3
R8323 plus.n30 plus.n29 161.3
R8324 plus.n32 plus.n31 161.3
R8325 plus.n33 plus.n4 161.3
R8326 plus.n36 plus.n35 161.3
R8327 plus.n37 plus.n3 161.3
R8328 plus.n39 plus.n38 161.3
R8329 plus.n41 plus.n2 161.3
R8330 plus.n43 plus.n42 161.3
R8331 plus.n45 plus.n44 161.3
R8332 plus.n46 plus.n0 161.3
R8333 plus.n48 plus.n47 161.3
R8334 plus.n64 plus.n63 56.5617
R8335 plus.n91 plus.n90 56.5617
R8336 plus.n42 plus.n41 56.5617
R8337 plus.n15 plus.n14 56.5617
R8338 plus.n73 plus.n72 56.5617
R8339 plus.n82 plus.n81 56.5617
R8340 plus.n33 plus.n32 56.5617
R8341 plus.n24 plus.n23 56.5617
R8342 plus.n95 plus.n94 48.3272
R8343 plus.n46 plus.n45 48.3272
R8344 plus.n70 plus.n58 44.4521
R8345 plus.n84 plus.n52 44.4521
R8346 plus.n35 plus.n3 44.4521
R8347 plus.n21 plus.n9 44.4521
R8348 plus.n62 plus.n61 43.0014
R8349 plus.n13 plus.n12 43.0014
R8350 plus.n77 plus.n76 40.577
R8351 plus.n78 plus.n77 40.577
R8352 plus.n29 plus.n28 40.577
R8353 plus.n28 plus.n27 40.577
R8354 plus.n61 plus.n60 39.4345
R8355 plus.n12 plus.n11 39.4345
R8356 plus.n66 plus.n58 36.702
R8357 plus.n88 plus.n52 36.702
R8358 plus.n39 plus.n3 36.702
R8359 plus.n17 plus.n9 36.702
R8360 plus.n98 plus.n97 33.3471
R8361 plus.n65 plus.n64 20.9036
R8362 plus.n90 plus.n89 20.9036
R8363 plus.n41 plus.n40 20.9036
R8364 plus.n16 plus.n15 20.9036
R8365 plus.n99 plus.t3 19.8005
R8366 plus.n99 plus.t2 19.8005
R8367 plus.n101 plus.t4 19.8005
R8368 plus.n101 plus.t0 19.8005
R8369 plus.n73 plus.n56 18.9362
R8370 plus.n81 plus.n54 18.9362
R8371 plus.n32 plus.n5 18.9362
R8372 plus.n24 plus.n7 18.9362
R8373 plus.n72 plus.n71 16.9689
R8374 plus.n83 plus.n82 16.9689
R8375 plus.n34 plus.n33 16.9689
R8376 plus.n23 plus.n22 16.9689
R8377 plus.n63 plus.n60 15.0015
R8378 plus.n91 plus.n50 15.0015
R8379 plus.n42 plus.n1 15.0015
R8380 plus.n14 plus.n11 15.0015
R8381 plus plus.n103 14.8715
R8382 plus.n96 plus.n95 12.4157
R8383 plus.n47 plus.n46 12.4157
R8384 plus.n98 plus.n48 11.9418
R8385 plus.n94 plus.n50 9.59132
R8386 plus.n45 plus.n1 9.59132
R8387 plus.n71 plus.n70 7.62397
R8388 plus.n84 plus.n83 7.62397
R8389 plus.n35 plus.n34 7.62397
R8390 plus.n22 plus.n21 7.62397
R8391 plus.n76 plus.n56 5.65662
R8392 plus.n78 plus.n54 5.65662
R8393 plus.n29 plus.n5 5.65662
R8394 plus.n27 plus.n7 5.65662
R8395 plus.n103 plus.n102 5.40567
R8396 plus.n66 plus.n65 3.68928
R8397 plus.n89 plus.n88 3.68928
R8398 plus.n40 plus.n39 3.68928
R8399 plus.n17 plus.n16 3.68928
R8400 plus.n103 plus.n98 1.188
R8401 plus.n102 plus.n100 0.716017
R8402 plus.n62 plus.n59 0.189894
R8403 plus.n67 plus.n59 0.189894
R8404 plus.n68 plus.n67 0.189894
R8405 plus.n69 plus.n68 0.189894
R8406 plus.n69 plus.n57 0.189894
R8407 plus.n74 plus.n57 0.189894
R8408 plus.n75 plus.n74 0.189894
R8409 plus.n75 plus.n55 0.189894
R8410 plus.n79 plus.n55 0.189894
R8411 plus.n80 plus.n79 0.189894
R8412 plus.n80 plus.n53 0.189894
R8413 plus.n85 plus.n53 0.189894
R8414 plus.n86 plus.n85 0.189894
R8415 plus.n87 plus.n86 0.189894
R8416 plus.n87 plus.n51 0.189894
R8417 plus.n92 plus.n51 0.189894
R8418 plus.n93 plus.n92 0.189894
R8419 plus.n93 plus.n49 0.189894
R8420 plus.n97 plus.n49 0.189894
R8421 plus.n48 plus.n0 0.189894
R8422 plus.n44 plus.n0 0.189894
R8423 plus.n44 plus.n43 0.189894
R8424 plus.n43 plus.n2 0.189894
R8425 plus.n38 plus.n2 0.189894
R8426 plus.n38 plus.n37 0.189894
R8427 plus.n37 plus.n36 0.189894
R8428 plus.n36 plus.n4 0.189894
R8429 plus.n31 plus.n4 0.189894
R8430 plus.n31 plus.n30 0.189894
R8431 plus.n30 plus.n6 0.189894
R8432 plus.n26 plus.n6 0.189894
R8433 plus.n26 plus.n25 0.189894
R8434 plus.n25 plus.n8 0.189894
R8435 plus.n20 plus.n8 0.189894
R8436 plus.n20 plus.n19 0.189894
R8437 plus.n19 plus.n18 0.189894
R8438 plus.n18 plus.n10 0.189894
R8439 plus.n13 plus.n10 0.189894
R8440 a_n3827_n3924.n12 a_n3827_n3924.t17 214.994
R8441 a_n3827_n3924.n1 a_n3827_n3924.t15 214.766
R8442 a_n3827_n3924.n13 a_n3827_n3924.t12 214.321
R8443 a_n3827_n3924.n14 a_n3827_n3924.t10 214.321
R8444 a_n3827_n3924.n15 a_n3827_n3924.t42 214.321
R8445 a_n3827_n3924.n16 a_n3827_n3924.t14 214.321
R8446 a_n3827_n3924.n17 a_n3827_n3924.t48 214.321
R8447 a_n3827_n3924.n18 a_n3827_n3924.t9 214.321
R8448 a_n3827_n3924.n19 a_n3827_n3924.t8 214.321
R8449 a_n3827_n3924.n12 a_n3827_n3924.t7 214.321
R8450 a_n3827_n3924.n0 a_n3827_n3924.t33 55.8337
R8451 a_n3827_n3924.n2 a_n3827_n3924.t2 55.8337
R8452 a_n3827_n3924.n11 a_n3827_n3924.t44 55.8337
R8453 a_n3827_n3924.n43 a_n3827_n3924.t21 55.8335
R8454 a_n3827_n3924.n41 a_n3827_n3924.t43 55.8335
R8455 a_n3827_n3924.n32 a_n3827_n3924.t13 55.8335
R8456 a_n3827_n3924.n31 a_n3827_n3924.t30 55.8335
R8457 a_n3827_n3924.n22 a_n3827_n3924.t38 55.8335
R8458 a_n3827_n3924.n45 a_n3827_n3924.n44 53.0052
R8459 a_n3827_n3924.n47 a_n3827_n3924.n46 53.0052
R8460 a_n3827_n3924.n49 a_n3827_n3924.n48 53.0052
R8461 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R8462 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R8463 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R8464 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R8465 a_n3827_n3924.n40 a_n3827_n3924.n39 53.0051
R8466 a_n3827_n3924.n38 a_n3827_n3924.n37 53.0051
R8467 a_n3827_n3924.n36 a_n3827_n3924.n35 53.0051
R8468 a_n3827_n3924.n34 a_n3827_n3924.n33 53.0051
R8469 a_n3827_n3924.n30 a_n3827_n3924.n29 53.0051
R8470 a_n3827_n3924.n28 a_n3827_n3924.n27 53.0051
R8471 a_n3827_n3924.n26 a_n3827_n3924.n25 53.0051
R8472 a_n3827_n3924.n24 a_n3827_n3924.n23 53.0051
R8473 a_n3827_n3924.n51 a_n3827_n3924.n50 53.0051
R8474 a_n3827_n3924.n21 a_n3827_n3924.n11 12.2417
R8475 a_n3827_n3924.n43 a_n3827_n3924.n42 12.2417
R8476 a_n3827_n3924.n22 a_n3827_n3924.n21 5.16214
R8477 a_n3827_n3924.n42 a_n3827_n3924.n41 5.16214
R8478 a_n3827_n3924.n44 a_n3827_n3924.t29 2.82907
R8479 a_n3827_n3924.n44 a_n3827_n3924.t34 2.82907
R8480 a_n3827_n3924.n46 a_n3827_n3924.t27 2.82907
R8481 a_n3827_n3924.n46 a_n3827_n3924.t31 2.82907
R8482 a_n3827_n3924.n48 a_n3827_n3924.t24 2.82907
R8483 a_n3827_n3924.n48 a_n3827_n3924.t28 2.82907
R8484 a_n3827_n3924.n3 a_n3827_n3924.t6 2.82907
R8485 a_n3827_n3924.n3 a_n3827_n3924.t5 2.82907
R8486 a_n3827_n3924.n5 a_n3827_n3924.t0 2.82907
R8487 a_n3827_n3924.n5 a_n3827_n3924.t19 2.82907
R8488 a_n3827_n3924.n7 a_n3827_n3924.t1 2.82907
R8489 a_n3827_n3924.n7 a_n3827_n3924.t4 2.82907
R8490 a_n3827_n3924.n9 a_n3827_n3924.t49 2.82907
R8491 a_n3827_n3924.n9 a_n3827_n3924.t47 2.82907
R8492 a_n3827_n3924.n39 a_n3827_n3924.t41 2.82907
R8493 a_n3827_n3924.n39 a_n3827_n3924.t18 2.82907
R8494 a_n3827_n3924.n37 a_n3827_n3924.t3 2.82907
R8495 a_n3827_n3924.n37 a_n3827_n3924.t45 2.82907
R8496 a_n3827_n3924.n35 a_n3827_n3924.t16 2.82907
R8497 a_n3827_n3924.n35 a_n3827_n3924.t40 2.82907
R8498 a_n3827_n3924.n33 a_n3827_n3924.t46 2.82907
R8499 a_n3827_n3924.n33 a_n3827_n3924.t11 2.82907
R8500 a_n3827_n3924.n29 a_n3827_n3924.t22 2.82907
R8501 a_n3827_n3924.n29 a_n3827_n3924.t35 2.82907
R8502 a_n3827_n3924.n27 a_n3827_n3924.t26 2.82907
R8503 a_n3827_n3924.n27 a_n3827_n3924.t20 2.82907
R8504 a_n3827_n3924.n25 a_n3827_n3924.t37 2.82907
R8505 a_n3827_n3924.n25 a_n3827_n3924.t25 2.82907
R8506 a_n3827_n3924.n23 a_n3827_n3924.t32 2.82907
R8507 a_n3827_n3924.n23 a_n3827_n3924.t36 2.82907
R8508 a_n3827_n3924.t39 a_n3827_n3924.n51 2.82907
R8509 a_n3827_n3924.n51 a_n3827_n3924.t23 2.82907
R8510 a_n3827_n3924.n42 a_n3827_n3924.n1 1.95694
R8511 a_n3827_n3924.n21 a_n3827_n3924.n20 1.95694
R8512 a_n3827_n3924.n19 a_n3827_n3924.n18 0.672012
R8513 a_n3827_n3924.n18 a_n3827_n3924.n17 0.672012
R8514 a_n3827_n3924.n17 a_n3827_n3924.n16 0.672012
R8515 a_n3827_n3924.n16 a_n3827_n3924.n15 0.672012
R8516 a_n3827_n3924.n15 a_n3827_n3924.n14 0.672012
R8517 a_n3827_n3924.n14 a_n3827_n3924.n13 0.672012
R8518 a_n3827_n3924.n24 a_n3827_n3924.n22 0.530672
R8519 a_n3827_n3924.n26 a_n3827_n3924.n24 0.530672
R8520 a_n3827_n3924.n28 a_n3827_n3924.n26 0.530672
R8521 a_n3827_n3924.n30 a_n3827_n3924.n28 0.530672
R8522 a_n3827_n3924.n31 a_n3827_n3924.n30 0.530672
R8523 a_n3827_n3924.n34 a_n3827_n3924.n32 0.530672
R8524 a_n3827_n3924.n36 a_n3827_n3924.n34 0.530672
R8525 a_n3827_n3924.n38 a_n3827_n3924.n36 0.530672
R8526 a_n3827_n3924.n40 a_n3827_n3924.n38 0.530672
R8527 a_n3827_n3924.n41 a_n3827_n3924.n40 0.530672
R8528 a_n3827_n3924.n11 a_n3827_n3924.n10 0.530672
R8529 a_n3827_n3924.n10 a_n3827_n3924.n8 0.530672
R8530 a_n3827_n3924.n8 a_n3827_n3924.n6 0.530672
R8531 a_n3827_n3924.n6 a_n3827_n3924.n4 0.530672
R8532 a_n3827_n3924.n4 a_n3827_n3924.n2 0.530672
R8533 a_n3827_n3924.n50 a_n3827_n3924.n0 0.530672
R8534 a_n3827_n3924.n50 a_n3827_n3924.n49 0.530672
R8535 a_n3827_n3924.n49 a_n3827_n3924.n47 0.530672
R8536 a_n3827_n3924.n47 a_n3827_n3924.n45 0.530672
R8537 a_n3827_n3924.n45 a_n3827_n3924.n43 0.530672
R8538 a_n3827_n3924.n20 a_n3827_n3924.n19 0.370413
R8539 a_n3827_n3924.n20 a_n3827_n3924.n12 0.302099
R8540 a_n3827_n3924.n32 a_n3827_n3924.n31 0.235414
R8541 a_n3827_n3924.n2 a_n3827_n3924.n0 0.235414
R8542 a_n3827_n3924.n13 a_n3827_n3924.n1 0.227971
R8543 gnd.n7186 gnd.n447 1638.19
R8544 gnd.n6490 gnd.n5138 939.716
R8545 gnd.n7580 gnd.n107 795.207
R8546 gnd.n7744 gnd.n103 795.207
R8547 gnd.n4479 gnd.n4478 795.207
R8548 gnd.n1688 gnd.n1687 795.207
R8549 gnd.n4899 gnd.n1324 795.207
R8550 gnd.n2792 gnd.n1322 795.207
R8551 gnd.n3020 gnd.n1008 795.207
R8552 gnd.n3083 gnd.n3021 795.207
R8553 gnd.n7742 gnd.n109 775.989
R8554 gnd.n178 gnd.n105 775.989
R8555 gnd.n1986 gnd.n1984 775.989
R8556 gnd.n1909 gnd.n1482 775.989
R8557 gnd.n4901 gnd.n1319 775.989
R8558 gnd.n3457 gnd.n1321 775.989
R8559 gnd.n5060 gnd.n5059 775.989
R8560 gnd.n5136 gnd.n1012 775.989
R8561 gnd.n967 gnd.n953 766.379
R8562 gnd.n6406 gnd.n6405 766.379
R8563 gnd.n5621 gnd.n5520 766.379
R8564 gnd.n5619 gnd.n5522 766.379
R8565 gnd.n6491 gnd.n958 756.769
R8566 gnd.n6392 gnd.n6391 756.769
R8567 gnd.n5753 gnd.n5482 756.769
R8568 gnd.n5739 gnd.n5471 756.769
R8569 gnd.n2838 gnd.n1329 711.122
R8570 gnd.n4741 gnd.n1455 711.122
R8571 gnd.n2721 gnd.n2665 711.122
R8572 gnd.n1798 gnd.n1457 711.122
R8573 gnd.n6694 gnd.n739 703.915
R8574 gnd.n7185 gnd.n448 703.915
R8575 gnd.n7398 gnd.n7397 703.915
R8576 gnd.n2923 gnd.n2920 703.915
R8577 gnd.n6694 gnd.n6693 585
R8578 gnd.n6695 gnd.n6694 585
R8579 gnd.n6692 gnd.n741 585
R8580 gnd.n741 gnd.n740 585
R8581 gnd.n6691 gnd.n6690 585
R8582 gnd.n6690 gnd.n6689 585
R8583 gnd.n746 gnd.n745 585
R8584 gnd.n6688 gnd.n746 585
R8585 gnd.n6686 gnd.n6685 585
R8586 gnd.n6687 gnd.n6686 585
R8587 gnd.n6684 gnd.n748 585
R8588 gnd.n748 gnd.n747 585
R8589 gnd.n6683 gnd.n6682 585
R8590 gnd.n6682 gnd.n6681 585
R8591 gnd.n754 gnd.n753 585
R8592 gnd.n6680 gnd.n754 585
R8593 gnd.n6678 gnd.n6677 585
R8594 gnd.n6679 gnd.n6678 585
R8595 gnd.n6676 gnd.n756 585
R8596 gnd.n756 gnd.n755 585
R8597 gnd.n6675 gnd.n6674 585
R8598 gnd.n6674 gnd.n6673 585
R8599 gnd.n762 gnd.n761 585
R8600 gnd.n6672 gnd.n762 585
R8601 gnd.n6670 gnd.n6669 585
R8602 gnd.n6671 gnd.n6670 585
R8603 gnd.n6668 gnd.n764 585
R8604 gnd.n764 gnd.n763 585
R8605 gnd.n6667 gnd.n6666 585
R8606 gnd.n6666 gnd.n6665 585
R8607 gnd.n770 gnd.n769 585
R8608 gnd.n6664 gnd.n770 585
R8609 gnd.n6662 gnd.n6661 585
R8610 gnd.n6663 gnd.n6662 585
R8611 gnd.n6660 gnd.n772 585
R8612 gnd.n772 gnd.n771 585
R8613 gnd.n6659 gnd.n6658 585
R8614 gnd.n6658 gnd.n6657 585
R8615 gnd.n778 gnd.n777 585
R8616 gnd.n6656 gnd.n778 585
R8617 gnd.n6654 gnd.n6653 585
R8618 gnd.n6655 gnd.n6654 585
R8619 gnd.n6652 gnd.n780 585
R8620 gnd.n780 gnd.n779 585
R8621 gnd.n6651 gnd.n6650 585
R8622 gnd.n6650 gnd.n6649 585
R8623 gnd.n786 gnd.n785 585
R8624 gnd.n6648 gnd.n786 585
R8625 gnd.n6646 gnd.n6645 585
R8626 gnd.n6647 gnd.n6646 585
R8627 gnd.n6644 gnd.n788 585
R8628 gnd.n788 gnd.n787 585
R8629 gnd.n6643 gnd.n6642 585
R8630 gnd.n6642 gnd.n6641 585
R8631 gnd.n794 gnd.n793 585
R8632 gnd.n6640 gnd.n794 585
R8633 gnd.n6638 gnd.n6637 585
R8634 gnd.n6639 gnd.n6638 585
R8635 gnd.n6636 gnd.n796 585
R8636 gnd.n796 gnd.n795 585
R8637 gnd.n6635 gnd.n6634 585
R8638 gnd.n6634 gnd.n6633 585
R8639 gnd.n802 gnd.n801 585
R8640 gnd.n6632 gnd.n802 585
R8641 gnd.n6630 gnd.n6629 585
R8642 gnd.n6631 gnd.n6630 585
R8643 gnd.n6628 gnd.n804 585
R8644 gnd.n804 gnd.n803 585
R8645 gnd.n6627 gnd.n6626 585
R8646 gnd.n6626 gnd.n6625 585
R8647 gnd.n810 gnd.n809 585
R8648 gnd.n6624 gnd.n810 585
R8649 gnd.n6622 gnd.n6621 585
R8650 gnd.n6623 gnd.n6622 585
R8651 gnd.n6620 gnd.n812 585
R8652 gnd.n812 gnd.n811 585
R8653 gnd.n6619 gnd.n6618 585
R8654 gnd.n6618 gnd.n6617 585
R8655 gnd.n818 gnd.n817 585
R8656 gnd.n6616 gnd.n818 585
R8657 gnd.n6614 gnd.n6613 585
R8658 gnd.n6615 gnd.n6614 585
R8659 gnd.n6612 gnd.n820 585
R8660 gnd.n820 gnd.n819 585
R8661 gnd.n6611 gnd.n6610 585
R8662 gnd.n6610 gnd.n6609 585
R8663 gnd.n826 gnd.n825 585
R8664 gnd.n6608 gnd.n826 585
R8665 gnd.n6606 gnd.n6605 585
R8666 gnd.n6607 gnd.n6606 585
R8667 gnd.n6604 gnd.n828 585
R8668 gnd.n828 gnd.n827 585
R8669 gnd.n6603 gnd.n6602 585
R8670 gnd.n6602 gnd.n6601 585
R8671 gnd.n834 gnd.n833 585
R8672 gnd.n6600 gnd.n834 585
R8673 gnd.n6598 gnd.n6597 585
R8674 gnd.n6599 gnd.n6598 585
R8675 gnd.n6596 gnd.n836 585
R8676 gnd.n836 gnd.n835 585
R8677 gnd.n6595 gnd.n6594 585
R8678 gnd.n6594 gnd.n6593 585
R8679 gnd.n842 gnd.n841 585
R8680 gnd.n6592 gnd.n842 585
R8681 gnd.n6590 gnd.n6589 585
R8682 gnd.n6591 gnd.n6590 585
R8683 gnd.n6588 gnd.n844 585
R8684 gnd.n844 gnd.n843 585
R8685 gnd.n6587 gnd.n6586 585
R8686 gnd.n6586 gnd.n6585 585
R8687 gnd.n850 gnd.n849 585
R8688 gnd.n6584 gnd.n850 585
R8689 gnd.n6582 gnd.n6581 585
R8690 gnd.n6583 gnd.n6582 585
R8691 gnd.n6580 gnd.n852 585
R8692 gnd.n852 gnd.n851 585
R8693 gnd.n6579 gnd.n6578 585
R8694 gnd.n6578 gnd.n6577 585
R8695 gnd.n858 gnd.n857 585
R8696 gnd.n6576 gnd.n858 585
R8697 gnd.n6574 gnd.n6573 585
R8698 gnd.n6575 gnd.n6574 585
R8699 gnd.n6572 gnd.n860 585
R8700 gnd.n860 gnd.n859 585
R8701 gnd.n6571 gnd.n6570 585
R8702 gnd.n6570 gnd.n6569 585
R8703 gnd.n866 gnd.n865 585
R8704 gnd.n6568 gnd.n866 585
R8705 gnd.n6566 gnd.n6565 585
R8706 gnd.n6567 gnd.n6566 585
R8707 gnd.n6564 gnd.n868 585
R8708 gnd.n868 gnd.n867 585
R8709 gnd.n6563 gnd.n6562 585
R8710 gnd.n6562 gnd.n6561 585
R8711 gnd.n874 gnd.n873 585
R8712 gnd.n6560 gnd.n874 585
R8713 gnd.n6558 gnd.n6557 585
R8714 gnd.n6559 gnd.n6558 585
R8715 gnd.n6556 gnd.n876 585
R8716 gnd.n876 gnd.n875 585
R8717 gnd.n6555 gnd.n6554 585
R8718 gnd.n6554 gnd.n6553 585
R8719 gnd.n882 gnd.n881 585
R8720 gnd.n6552 gnd.n882 585
R8721 gnd.n6550 gnd.n6549 585
R8722 gnd.n6551 gnd.n6550 585
R8723 gnd.n6548 gnd.n884 585
R8724 gnd.n884 gnd.n883 585
R8725 gnd.n6547 gnd.n6546 585
R8726 gnd.n6546 gnd.n6545 585
R8727 gnd.n890 gnd.n889 585
R8728 gnd.n6544 gnd.n890 585
R8729 gnd.n6542 gnd.n6541 585
R8730 gnd.n6543 gnd.n6542 585
R8731 gnd.n6540 gnd.n892 585
R8732 gnd.n892 gnd.n891 585
R8733 gnd.n6539 gnd.n6538 585
R8734 gnd.n6538 gnd.n6537 585
R8735 gnd.n898 gnd.n897 585
R8736 gnd.n6536 gnd.n898 585
R8737 gnd.n6534 gnd.n6533 585
R8738 gnd.n6535 gnd.n6534 585
R8739 gnd.n6532 gnd.n900 585
R8740 gnd.n900 gnd.n899 585
R8741 gnd.n6531 gnd.n6530 585
R8742 gnd.n6530 gnd.n6529 585
R8743 gnd.n906 gnd.n905 585
R8744 gnd.n6528 gnd.n906 585
R8745 gnd.n739 gnd.n738 585
R8746 gnd.n6696 gnd.n739 585
R8747 gnd.n6699 gnd.n6698 585
R8748 gnd.n6698 gnd.n6697 585
R8749 gnd.n736 gnd.n735 585
R8750 gnd.n735 gnd.n734 585
R8751 gnd.n6704 gnd.n6703 585
R8752 gnd.n6705 gnd.n6704 585
R8753 gnd.n733 gnd.n732 585
R8754 gnd.n6706 gnd.n733 585
R8755 gnd.n6709 gnd.n6708 585
R8756 gnd.n6708 gnd.n6707 585
R8757 gnd.n730 gnd.n729 585
R8758 gnd.n729 gnd.n728 585
R8759 gnd.n6714 gnd.n6713 585
R8760 gnd.n6715 gnd.n6714 585
R8761 gnd.n727 gnd.n726 585
R8762 gnd.n6716 gnd.n727 585
R8763 gnd.n6719 gnd.n6718 585
R8764 gnd.n6718 gnd.n6717 585
R8765 gnd.n724 gnd.n723 585
R8766 gnd.n723 gnd.n722 585
R8767 gnd.n6724 gnd.n6723 585
R8768 gnd.n6725 gnd.n6724 585
R8769 gnd.n721 gnd.n720 585
R8770 gnd.n6726 gnd.n721 585
R8771 gnd.n6729 gnd.n6728 585
R8772 gnd.n6728 gnd.n6727 585
R8773 gnd.n718 gnd.n717 585
R8774 gnd.n717 gnd.n716 585
R8775 gnd.n6734 gnd.n6733 585
R8776 gnd.n6735 gnd.n6734 585
R8777 gnd.n715 gnd.n714 585
R8778 gnd.n6736 gnd.n715 585
R8779 gnd.n6739 gnd.n6738 585
R8780 gnd.n6738 gnd.n6737 585
R8781 gnd.n712 gnd.n711 585
R8782 gnd.n711 gnd.n710 585
R8783 gnd.n6744 gnd.n6743 585
R8784 gnd.n6745 gnd.n6744 585
R8785 gnd.n709 gnd.n708 585
R8786 gnd.n6746 gnd.n709 585
R8787 gnd.n6749 gnd.n6748 585
R8788 gnd.n6748 gnd.n6747 585
R8789 gnd.n706 gnd.n705 585
R8790 gnd.n705 gnd.n704 585
R8791 gnd.n6754 gnd.n6753 585
R8792 gnd.n6755 gnd.n6754 585
R8793 gnd.n703 gnd.n702 585
R8794 gnd.n6756 gnd.n703 585
R8795 gnd.n6759 gnd.n6758 585
R8796 gnd.n6758 gnd.n6757 585
R8797 gnd.n700 gnd.n699 585
R8798 gnd.n699 gnd.n698 585
R8799 gnd.n6764 gnd.n6763 585
R8800 gnd.n6765 gnd.n6764 585
R8801 gnd.n697 gnd.n696 585
R8802 gnd.n6766 gnd.n697 585
R8803 gnd.n6769 gnd.n6768 585
R8804 gnd.n6768 gnd.n6767 585
R8805 gnd.n694 gnd.n693 585
R8806 gnd.n693 gnd.n692 585
R8807 gnd.n6774 gnd.n6773 585
R8808 gnd.n6775 gnd.n6774 585
R8809 gnd.n691 gnd.n690 585
R8810 gnd.n6776 gnd.n691 585
R8811 gnd.n6779 gnd.n6778 585
R8812 gnd.n6778 gnd.n6777 585
R8813 gnd.n688 gnd.n687 585
R8814 gnd.n687 gnd.n686 585
R8815 gnd.n6784 gnd.n6783 585
R8816 gnd.n6785 gnd.n6784 585
R8817 gnd.n685 gnd.n684 585
R8818 gnd.n6786 gnd.n685 585
R8819 gnd.n6789 gnd.n6788 585
R8820 gnd.n6788 gnd.n6787 585
R8821 gnd.n682 gnd.n681 585
R8822 gnd.n681 gnd.n680 585
R8823 gnd.n6794 gnd.n6793 585
R8824 gnd.n6795 gnd.n6794 585
R8825 gnd.n679 gnd.n678 585
R8826 gnd.n6796 gnd.n679 585
R8827 gnd.n6799 gnd.n6798 585
R8828 gnd.n6798 gnd.n6797 585
R8829 gnd.n676 gnd.n675 585
R8830 gnd.n675 gnd.n674 585
R8831 gnd.n6804 gnd.n6803 585
R8832 gnd.n6805 gnd.n6804 585
R8833 gnd.n673 gnd.n672 585
R8834 gnd.n6806 gnd.n673 585
R8835 gnd.n6809 gnd.n6808 585
R8836 gnd.n6808 gnd.n6807 585
R8837 gnd.n670 gnd.n669 585
R8838 gnd.n669 gnd.n668 585
R8839 gnd.n6814 gnd.n6813 585
R8840 gnd.n6815 gnd.n6814 585
R8841 gnd.n667 gnd.n666 585
R8842 gnd.n6816 gnd.n667 585
R8843 gnd.n6819 gnd.n6818 585
R8844 gnd.n6818 gnd.n6817 585
R8845 gnd.n664 gnd.n663 585
R8846 gnd.n663 gnd.n662 585
R8847 gnd.n6824 gnd.n6823 585
R8848 gnd.n6825 gnd.n6824 585
R8849 gnd.n661 gnd.n660 585
R8850 gnd.n6826 gnd.n661 585
R8851 gnd.n6829 gnd.n6828 585
R8852 gnd.n6828 gnd.n6827 585
R8853 gnd.n658 gnd.n657 585
R8854 gnd.n657 gnd.n656 585
R8855 gnd.n6834 gnd.n6833 585
R8856 gnd.n6835 gnd.n6834 585
R8857 gnd.n655 gnd.n654 585
R8858 gnd.n6836 gnd.n655 585
R8859 gnd.n6839 gnd.n6838 585
R8860 gnd.n6838 gnd.n6837 585
R8861 gnd.n652 gnd.n651 585
R8862 gnd.n651 gnd.n650 585
R8863 gnd.n6844 gnd.n6843 585
R8864 gnd.n6845 gnd.n6844 585
R8865 gnd.n649 gnd.n648 585
R8866 gnd.n6846 gnd.n649 585
R8867 gnd.n6849 gnd.n6848 585
R8868 gnd.n6848 gnd.n6847 585
R8869 gnd.n646 gnd.n645 585
R8870 gnd.n645 gnd.n644 585
R8871 gnd.n6854 gnd.n6853 585
R8872 gnd.n6855 gnd.n6854 585
R8873 gnd.n643 gnd.n642 585
R8874 gnd.n6856 gnd.n643 585
R8875 gnd.n6859 gnd.n6858 585
R8876 gnd.n6858 gnd.n6857 585
R8877 gnd.n640 gnd.n639 585
R8878 gnd.n639 gnd.n638 585
R8879 gnd.n6864 gnd.n6863 585
R8880 gnd.n6865 gnd.n6864 585
R8881 gnd.n637 gnd.n636 585
R8882 gnd.n6866 gnd.n637 585
R8883 gnd.n6869 gnd.n6868 585
R8884 gnd.n6868 gnd.n6867 585
R8885 gnd.n634 gnd.n633 585
R8886 gnd.n633 gnd.n632 585
R8887 gnd.n6874 gnd.n6873 585
R8888 gnd.n6875 gnd.n6874 585
R8889 gnd.n631 gnd.n630 585
R8890 gnd.n6876 gnd.n631 585
R8891 gnd.n6879 gnd.n6878 585
R8892 gnd.n6878 gnd.n6877 585
R8893 gnd.n628 gnd.n627 585
R8894 gnd.n627 gnd.n626 585
R8895 gnd.n6884 gnd.n6883 585
R8896 gnd.n6885 gnd.n6884 585
R8897 gnd.n625 gnd.n624 585
R8898 gnd.n6886 gnd.n625 585
R8899 gnd.n6889 gnd.n6888 585
R8900 gnd.n6888 gnd.n6887 585
R8901 gnd.n622 gnd.n621 585
R8902 gnd.n621 gnd.n620 585
R8903 gnd.n6894 gnd.n6893 585
R8904 gnd.n6895 gnd.n6894 585
R8905 gnd.n619 gnd.n618 585
R8906 gnd.n6896 gnd.n619 585
R8907 gnd.n6899 gnd.n6898 585
R8908 gnd.n6898 gnd.n6897 585
R8909 gnd.n616 gnd.n615 585
R8910 gnd.n615 gnd.n614 585
R8911 gnd.n6904 gnd.n6903 585
R8912 gnd.n6905 gnd.n6904 585
R8913 gnd.n613 gnd.n612 585
R8914 gnd.n6906 gnd.n613 585
R8915 gnd.n6909 gnd.n6908 585
R8916 gnd.n6908 gnd.n6907 585
R8917 gnd.n610 gnd.n609 585
R8918 gnd.n609 gnd.n608 585
R8919 gnd.n6914 gnd.n6913 585
R8920 gnd.n6915 gnd.n6914 585
R8921 gnd.n607 gnd.n606 585
R8922 gnd.n6916 gnd.n607 585
R8923 gnd.n6919 gnd.n6918 585
R8924 gnd.n6918 gnd.n6917 585
R8925 gnd.n604 gnd.n603 585
R8926 gnd.n603 gnd.n602 585
R8927 gnd.n6924 gnd.n6923 585
R8928 gnd.n6925 gnd.n6924 585
R8929 gnd.n601 gnd.n600 585
R8930 gnd.n6926 gnd.n601 585
R8931 gnd.n6929 gnd.n6928 585
R8932 gnd.n6928 gnd.n6927 585
R8933 gnd.n598 gnd.n597 585
R8934 gnd.n597 gnd.n596 585
R8935 gnd.n6934 gnd.n6933 585
R8936 gnd.n6935 gnd.n6934 585
R8937 gnd.n595 gnd.n594 585
R8938 gnd.n6936 gnd.n595 585
R8939 gnd.n6939 gnd.n6938 585
R8940 gnd.n6938 gnd.n6937 585
R8941 gnd.n592 gnd.n591 585
R8942 gnd.n591 gnd.n590 585
R8943 gnd.n6944 gnd.n6943 585
R8944 gnd.n6945 gnd.n6944 585
R8945 gnd.n589 gnd.n588 585
R8946 gnd.n6946 gnd.n589 585
R8947 gnd.n6949 gnd.n6948 585
R8948 gnd.n6948 gnd.n6947 585
R8949 gnd.n586 gnd.n585 585
R8950 gnd.n585 gnd.n584 585
R8951 gnd.n6954 gnd.n6953 585
R8952 gnd.n6955 gnd.n6954 585
R8953 gnd.n583 gnd.n582 585
R8954 gnd.n6956 gnd.n583 585
R8955 gnd.n6959 gnd.n6958 585
R8956 gnd.n6958 gnd.n6957 585
R8957 gnd.n580 gnd.n579 585
R8958 gnd.n579 gnd.n578 585
R8959 gnd.n6964 gnd.n6963 585
R8960 gnd.n6965 gnd.n6964 585
R8961 gnd.n577 gnd.n576 585
R8962 gnd.n6966 gnd.n577 585
R8963 gnd.n6969 gnd.n6968 585
R8964 gnd.n6968 gnd.n6967 585
R8965 gnd.n574 gnd.n573 585
R8966 gnd.n573 gnd.n572 585
R8967 gnd.n6974 gnd.n6973 585
R8968 gnd.n6975 gnd.n6974 585
R8969 gnd.n571 gnd.n570 585
R8970 gnd.n6976 gnd.n571 585
R8971 gnd.n6979 gnd.n6978 585
R8972 gnd.n6978 gnd.n6977 585
R8973 gnd.n568 gnd.n567 585
R8974 gnd.n567 gnd.n566 585
R8975 gnd.n6984 gnd.n6983 585
R8976 gnd.n6985 gnd.n6984 585
R8977 gnd.n565 gnd.n564 585
R8978 gnd.n6986 gnd.n565 585
R8979 gnd.n6989 gnd.n6988 585
R8980 gnd.n6988 gnd.n6987 585
R8981 gnd.n562 gnd.n561 585
R8982 gnd.n561 gnd.n560 585
R8983 gnd.n6994 gnd.n6993 585
R8984 gnd.n6995 gnd.n6994 585
R8985 gnd.n559 gnd.n558 585
R8986 gnd.n6996 gnd.n559 585
R8987 gnd.n6999 gnd.n6998 585
R8988 gnd.n6998 gnd.n6997 585
R8989 gnd.n556 gnd.n555 585
R8990 gnd.n555 gnd.n554 585
R8991 gnd.n7004 gnd.n7003 585
R8992 gnd.n7005 gnd.n7004 585
R8993 gnd.n553 gnd.n552 585
R8994 gnd.n7006 gnd.n553 585
R8995 gnd.n7009 gnd.n7008 585
R8996 gnd.n7008 gnd.n7007 585
R8997 gnd.n550 gnd.n549 585
R8998 gnd.n549 gnd.n548 585
R8999 gnd.n7014 gnd.n7013 585
R9000 gnd.n7015 gnd.n7014 585
R9001 gnd.n547 gnd.n546 585
R9002 gnd.n7016 gnd.n547 585
R9003 gnd.n7019 gnd.n7018 585
R9004 gnd.n7018 gnd.n7017 585
R9005 gnd.n544 gnd.n543 585
R9006 gnd.n543 gnd.n542 585
R9007 gnd.n7024 gnd.n7023 585
R9008 gnd.n7025 gnd.n7024 585
R9009 gnd.n541 gnd.n540 585
R9010 gnd.n7026 gnd.n541 585
R9011 gnd.n7029 gnd.n7028 585
R9012 gnd.n7028 gnd.n7027 585
R9013 gnd.n538 gnd.n537 585
R9014 gnd.n537 gnd.n536 585
R9015 gnd.n7034 gnd.n7033 585
R9016 gnd.n7035 gnd.n7034 585
R9017 gnd.n535 gnd.n534 585
R9018 gnd.n7036 gnd.n535 585
R9019 gnd.n7039 gnd.n7038 585
R9020 gnd.n7038 gnd.n7037 585
R9021 gnd.n532 gnd.n531 585
R9022 gnd.n531 gnd.n530 585
R9023 gnd.n7044 gnd.n7043 585
R9024 gnd.n7045 gnd.n7044 585
R9025 gnd.n529 gnd.n528 585
R9026 gnd.n7046 gnd.n529 585
R9027 gnd.n7049 gnd.n7048 585
R9028 gnd.n7048 gnd.n7047 585
R9029 gnd.n526 gnd.n525 585
R9030 gnd.n525 gnd.n524 585
R9031 gnd.n7054 gnd.n7053 585
R9032 gnd.n7055 gnd.n7054 585
R9033 gnd.n523 gnd.n522 585
R9034 gnd.n7056 gnd.n523 585
R9035 gnd.n7059 gnd.n7058 585
R9036 gnd.n7058 gnd.n7057 585
R9037 gnd.n520 gnd.n519 585
R9038 gnd.n519 gnd.n518 585
R9039 gnd.n7064 gnd.n7063 585
R9040 gnd.n7065 gnd.n7064 585
R9041 gnd.n517 gnd.n516 585
R9042 gnd.n7066 gnd.n517 585
R9043 gnd.n7069 gnd.n7068 585
R9044 gnd.n7068 gnd.n7067 585
R9045 gnd.n514 gnd.n513 585
R9046 gnd.n513 gnd.n512 585
R9047 gnd.n7074 gnd.n7073 585
R9048 gnd.n7075 gnd.n7074 585
R9049 gnd.n511 gnd.n510 585
R9050 gnd.n7076 gnd.n511 585
R9051 gnd.n7079 gnd.n7078 585
R9052 gnd.n7078 gnd.n7077 585
R9053 gnd.n508 gnd.n507 585
R9054 gnd.n507 gnd.n506 585
R9055 gnd.n7084 gnd.n7083 585
R9056 gnd.n7085 gnd.n7084 585
R9057 gnd.n505 gnd.n504 585
R9058 gnd.n7086 gnd.n505 585
R9059 gnd.n7089 gnd.n7088 585
R9060 gnd.n7088 gnd.n7087 585
R9061 gnd.n502 gnd.n501 585
R9062 gnd.n501 gnd.n500 585
R9063 gnd.n7094 gnd.n7093 585
R9064 gnd.n7095 gnd.n7094 585
R9065 gnd.n499 gnd.n498 585
R9066 gnd.n7096 gnd.n499 585
R9067 gnd.n7099 gnd.n7098 585
R9068 gnd.n7098 gnd.n7097 585
R9069 gnd.n496 gnd.n495 585
R9070 gnd.n495 gnd.n494 585
R9071 gnd.n7104 gnd.n7103 585
R9072 gnd.n7105 gnd.n7104 585
R9073 gnd.n493 gnd.n492 585
R9074 gnd.n7106 gnd.n493 585
R9075 gnd.n7109 gnd.n7108 585
R9076 gnd.n7108 gnd.n7107 585
R9077 gnd.n490 gnd.n489 585
R9078 gnd.n489 gnd.n488 585
R9079 gnd.n7114 gnd.n7113 585
R9080 gnd.n7115 gnd.n7114 585
R9081 gnd.n487 gnd.n486 585
R9082 gnd.n7116 gnd.n487 585
R9083 gnd.n7119 gnd.n7118 585
R9084 gnd.n7118 gnd.n7117 585
R9085 gnd.n484 gnd.n483 585
R9086 gnd.n483 gnd.n482 585
R9087 gnd.n7124 gnd.n7123 585
R9088 gnd.n7125 gnd.n7124 585
R9089 gnd.n481 gnd.n480 585
R9090 gnd.n7126 gnd.n481 585
R9091 gnd.n7129 gnd.n7128 585
R9092 gnd.n7128 gnd.n7127 585
R9093 gnd.n478 gnd.n477 585
R9094 gnd.n477 gnd.n476 585
R9095 gnd.n7134 gnd.n7133 585
R9096 gnd.n7135 gnd.n7134 585
R9097 gnd.n475 gnd.n474 585
R9098 gnd.n7136 gnd.n475 585
R9099 gnd.n7139 gnd.n7138 585
R9100 gnd.n7138 gnd.n7137 585
R9101 gnd.n472 gnd.n471 585
R9102 gnd.n471 gnd.n470 585
R9103 gnd.n7144 gnd.n7143 585
R9104 gnd.n7145 gnd.n7144 585
R9105 gnd.n469 gnd.n468 585
R9106 gnd.n7146 gnd.n469 585
R9107 gnd.n7149 gnd.n7148 585
R9108 gnd.n7148 gnd.n7147 585
R9109 gnd.n466 gnd.n465 585
R9110 gnd.n465 gnd.n464 585
R9111 gnd.n7154 gnd.n7153 585
R9112 gnd.n7155 gnd.n7154 585
R9113 gnd.n463 gnd.n462 585
R9114 gnd.n7156 gnd.n463 585
R9115 gnd.n7159 gnd.n7158 585
R9116 gnd.n7158 gnd.n7157 585
R9117 gnd.n460 gnd.n459 585
R9118 gnd.n459 gnd.n458 585
R9119 gnd.n7164 gnd.n7163 585
R9120 gnd.n7165 gnd.n7164 585
R9121 gnd.n457 gnd.n456 585
R9122 gnd.n7166 gnd.n457 585
R9123 gnd.n7169 gnd.n7168 585
R9124 gnd.n7168 gnd.n7167 585
R9125 gnd.n454 gnd.n453 585
R9126 gnd.n453 gnd.n452 585
R9127 gnd.n7175 gnd.n7174 585
R9128 gnd.n7176 gnd.n7175 585
R9129 gnd.n451 gnd.n450 585
R9130 gnd.n7177 gnd.n451 585
R9131 gnd.n7180 gnd.n7179 585
R9132 gnd.n7179 gnd.n7178 585
R9133 gnd.n7181 gnd.n448 585
R9134 gnd.n448 gnd.n447 585
R9135 gnd.n323 gnd.n322 585
R9136 gnd.n7388 gnd.n322 585
R9137 gnd.n7391 gnd.n7390 585
R9138 gnd.n7390 gnd.n7389 585
R9139 gnd.n326 gnd.n325 585
R9140 gnd.n7387 gnd.n326 585
R9141 gnd.n7385 gnd.n7384 585
R9142 gnd.n7386 gnd.n7385 585
R9143 gnd.n329 gnd.n328 585
R9144 gnd.n328 gnd.n327 585
R9145 gnd.n7380 gnd.n7379 585
R9146 gnd.n7379 gnd.n7378 585
R9147 gnd.n332 gnd.n331 585
R9148 gnd.n7377 gnd.n332 585
R9149 gnd.n7375 gnd.n7374 585
R9150 gnd.n7376 gnd.n7375 585
R9151 gnd.n335 gnd.n334 585
R9152 gnd.n334 gnd.n333 585
R9153 gnd.n7370 gnd.n7369 585
R9154 gnd.n7369 gnd.n7368 585
R9155 gnd.n338 gnd.n337 585
R9156 gnd.n7367 gnd.n338 585
R9157 gnd.n7365 gnd.n7364 585
R9158 gnd.n7366 gnd.n7365 585
R9159 gnd.n341 gnd.n340 585
R9160 gnd.n340 gnd.n339 585
R9161 gnd.n7360 gnd.n7359 585
R9162 gnd.n7359 gnd.n7358 585
R9163 gnd.n344 gnd.n343 585
R9164 gnd.n7357 gnd.n344 585
R9165 gnd.n7355 gnd.n7354 585
R9166 gnd.n7356 gnd.n7355 585
R9167 gnd.n347 gnd.n346 585
R9168 gnd.n346 gnd.n345 585
R9169 gnd.n7350 gnd.n7349 585
R9170 gnd.n7349 gnd.n7348 585
R9171 gnd.n350 gnd.n349 585
R9172 gnd.n7347 gnd.n350 585
R9173 gnd.n7345 gnd.n7344 585
R9174 gnd.n7346 gnd.n7345 585
R9175 gnd.n353 gnd.n352 585
R9176 gnd.n352 gnd.n351 585
R9177 gnd.n7340 gnd.n7339 585
R9178 gnd.n7339 gnd.n7338 585
R9179 gnd.n356 gnd.n355 585
R9180 gnd.n7337 gnd.n356 585
R9181 gnd.n7335 gnd.n7334 585
R9182 gnd.n7336 gnd.n7335 585
R9183 gnd.n359 gnd.n358 585
R9184 gnd.n358 gnd.n357 585
R9185 gnd.n7330 gnd.n7329 585
R9186 gnd.n7329 gnd.n7328 585
R9187 gnd.n362 gnd.n361 585
R9188 gnd.n7327 gnd.n362 585
R9189 gnd.n7325 gnd.n7324 585
R9190 gnd.n7326 gnd.n7325 585
R9191 gnd.n365 gnd.n364 585
R9192 gnd.n364 gnd.n363 585
R9193 gnd.n7320 gnd.n7319 585
R9194 gnd.n7319 gnd.n7318 585
R9195 gnd.n368 gnd.n367 585
R9196 gnd.n7317 gnd.n368 585
R9197 gnd.n7315 gnd.n7314 585
R9198 gnd.n7316 gnd.n7315 585
R9199 gnd.n371 gnd.n370 585
R9200 gnd.n370 gnd.n369 585
R9201 gnd.n7310 gnd.n7309 585
R9202 gnd.n7309 gnd.n7308 585
R9203 gnd.n374 gnd.n373 585
R9204 gnd.n7307 gnd.n374 585
R9205 gnd.n7305 gnd.n7304 585
R9206 gnd.n7306 gnd.n7305 585
R9207 gnd.n377 gnd.n376 585
R9208 gnd.n376 gnd.n375 585
R9209 gnd.n7300 gnd.n7299 585
R9210 gnd.n7299 gnd.n7298 585
R9211 gnd.n380 gnd.n379 585
R9212 gnd.n7297 gnd.n380 585
R9213 gnd.n7295 gnd.n7294 585
R9214 gnd.n7296 gnd.n7295 585
R9215 gnd.n383 gnd.n382 585
R9216 gnd.n382 gnd.n381 585
R9217 gnd.n7290 gnd.n7289 585
R9218 gnd.n7289 gnd.n7288 585
R9219 gnd.n386 gnd.n385 585
R9220 gnd.n7287 gnd.n386 585
R9221 gnd.n7285 gnd.n7284 585
R9222 gnd.n7286 gnd.n7285 585
R9223 gnd.n389 gnd.n388 585
R9224 gnd.n388 gnd.n387 585
R9225 gnd.n7280 gnd.n7279 585
R9226 gnd.n7279 gnd.n7278 585
R9227 gnd.n392 gnd.n391 585
R9228 gnd.n7277 gnd.n392 585
R9229 gnd.n7275 gnd.n7274 585
R9230 gnd.n7276 gnd.n7275 585
R9231 gnd.n395 gnd.n394 585
R9232 gnd.n394 gnd.n393 585
R9233 gnd.n7270 gnd.n7269 585
R9234 gnd.n7269 gnd.n7268 585
R9235 gnd.n398 gnd.n397 585
R9236 gnd.n7267 gnd.n398 585
R9237 gnd.n7265 gnd.n7264 585
R9238 gnd.n7266 gnd.n7265 585
R9239 gnd.n401 gnd.n400 585
R9240 gnd.n400 gnd.n399 585
R9241 gnd.n7260 gnd.n7259 585
R9242 gnd.n7259 gnd.n7258 585
R9243 gnd.n404 gnd.n403 585
R9244 gnd.n7257 gnd.n404 585
R9245 gnd.n7255 gnd.n7254 585
R9246 gnd.n7256 gnd.n7255 585
R9247 gnd.n407 gnd.n406 585
R9248 gnd.n406 gnd.n405 585
R9249 gnd.n7250 gnd.n7249 585
R9250 gnd.n7249 gnd.n7248 585
R9251 gnd.n410 gnd.n409 585
R9252 gnd.n7247 gnd.n410 585
R9253 gnd.n7245 gnd.n7244 585
R9254 gnd.n7246 gnd.n7245 585
R9255 gnd.n413 gnd.n412 585
R9256 gnd.n412 gnd.n411 585
R9257 gnd.n7240 gnd.n7239 585
R9258 gnd.n7239 gnd.n7238 585
R9259 gnd.n416 gnd.n415 585
R9260 gnd.n7237 gnd.n416 585
R9261 gnd.n7235 gnd.n7234 585
R9262 gnd.n7236 gnd.n7235 585
R9263 gnd.n419 gnd.n418 585
R9264 gnd.n418 gnd.n417 585
R9265 gnd.n7230 gnd.n7229 585
R9266 gnd.n7229 gnd.n7228 585
R9267 gnd.n422 gnd.n421 585
R9268 gnd.n7227 gnd.n422 585
R9269 gnd.n7225 gnd.n7224 585
R9270 gnd.n7226 gnd.n7225 585
R9271 gnd.n425 gnd.n424 585
R9272 gnd.n424 gnd.n423 585
R9273 gnd.n7220 gnd.n7219 585
R9274 gnd.n7219 gnd.n7218 585
R9275 gnd.n428 gnd.n427 585
R9276 gnd.n7217 gnd.n428 585
R9277 gnd.n7215 gnd.n7214 585
R9278 gnd.n7216 gnd.n7215 585
R9279 gnd.n431 gnd.n430 585
R9280 gnd.n430 gnd.n429 585
R9281 gnd.n7210 gnd.n7209 585
R9282 gnd.n7209 gnd.n7208 585
R9283 gnd.n434 gnd.n433 585
R9284 gnd.n7207 gnd.n434 585
R9285 gnd.n7205 gnd.n7204 585
R9286 gnd.n7206 gnd.n7205 585
R9287 gnd.n437 gnd.n436 585
R9288 gnd.n436 gnd.n435 585
R9289 gnd.n7200 gnd.n7199 585
R9290 gnd.n7199 gnd.n7198 585
R9291 gnd.n440 gnd.n439 585
R9292 gnd.n7197 gnd.n440 585
R9293 gnd.n7195 gnd.n7194 585
R9294 gnd.n7196 gnd.n7195 585
R9295 gnd.n443 gnd.n442 585
R9296 gnd.n442 gnd.n441 585
R9297 gnd.n7190 gnd.n7189 585
R9298 gnd.n7189 gnd.n7188 585
R9299 gnd.n446 gnd.n445 585
R9300 gnd.n7187 gnd.n446 585
R9301 gnd.n7185 gnd.n7184 585
R9302 gnd.n7186 gnd.n7185 585
R9303 gnd.n4899 gnd.n4898 585
R9304 gnd.n4900 gnd.n4899 585
R9305 gnd.n1310 gnd.n1309 585
R9306 gnd.n3450 gnd.n1310 585
R9307 gnd.n4908 gnd.n4907 585
R9308 gnd.n4907 gnd.n4906 585
R9309 gnd.n4909 gnd.n1304 585
R9310 gnd.n3285 gnd.n1304 585
R9311 gnd.n4911 gnd.n4910 585
R9312 gnd.n4912 gnd.n4911 585
R9313 gnd.n1288 gnd.n1287 585
R9314 gnd.n3276 gnd.n1288 585
R9315 gnd.n4920 gnd.n4919 585
R9316 gnd.n4919 gnd.n4918 585
R9317 gnd.n4921 gnd.n1282 585
R9318 gnd.n3272 gnd.n1282 585
R9319 gnd.n4923 gnd.n4922 585
R9320 gnd.n4924 gnd.n4923 585
R9321 gnd.n1267 gnd.n1266 585
R9322 gnd.n3299 gnd.n1267 585
R9323 gnd.n4932 gnd.n4931 585
R9324 gnd.n4931 gnd.n4930 585
R9325 gnd.n4933 gnd.n1261 585
R9326 gnd.n3264 gnd.n1261 585
R9327 gnd.n4935 gnd.n4934 585
R9328 gnd.n4936 gnd.n4935 585
R9329 gnd.n1246 gnd.n1245 585
R9330 gnd.n3256 gnd.n1246 585
R9331 gnd.n4944 gnd.n4943 585
R9332 gnd.n4943 gnd.n4942 585
R9333 gnd.n4945 gnd.n1240 585
R9334 gnd.n3247 gnd.n1240 585
R9335 gnd.n4947 gnd.n4946 585
R9336 gnd.n4948 gnd.n4947 585
R9337 gnd.n1225 gnd.n1224 585
R9338 gnd.n3239 gnd.n1225 585
R9339 gnd.n4956 gnd.n4955 585
R9340 gnd.n4955 gnd.n4954 585
R9341 gnd.n4957 gnd.n1219 585
R9342 gnd.n3231 gnd.n1219 585
R9343 gnd.n4959 gnd.n4958 585
R9344 gnd.n4960 gnd.n4959 585
R9345 gnd.n1205 gnd.n1204 585
R9346 gnd.n3223 gnd.n1205 585
R9347 gnd.n4968 gnd.n4967 585
R9348 gnd.n4967 gnd.n4966 585
R9349 gnd.n4969 gnd.n1199 585
R9350 gnd.n3215 gnd.n1199 585
R9351 gnd.n4971 gnd.n4970 585
R9352 gnd.n4972 gnd.n4971 585
R9353 gnd.n1187 gnd.n1186 585
R9354 gnd.n3207 gnd.n1187 585
R9355 gnd.n4981 gnd.n4980 585
R9356 gnd.n4980 gnd.n4979 585
R9357 gnd.n4982 gnd.n1181 585
R9358 gnd.n3198 gnd.n1181 585
R9359 gnd.n4984 gnd.n4983 585
R9360 gnd.n4985 gnd.n4984 585
R9361 gnd.n1168 gnd.n1167 585
R9362 gnd.n3189 gnd.n1168 585
R9363 gnd.n4993 gnd.n4992 585
R9364 gnd.n4992 gnd.n4991 585
R9365 gnd.n4994 gnd.n1162 585
R9366 gnd.n3181 gnd.n1162 585
R9367 gnd.n4996 gnd.n4995 585
R9368 gnd.n4997 gnd.n4996 585
R9369 gnd.n1147 gnd.n1146 585
R9370 gnd.n3173 gnd.n1147 585
R9371 gnd.n5005 gnd.n5004 585
R9372 gnd.n5004 gnd.n5003 585
R9373 gnd.n5006 gnd.n1141 585
R9374 gnd.n3165 gnd.n1141 585
R9375 gnd.n5008 gnd.n5007 585
R9376 gnd.n5009 gnd.n5008 585
R9377 gnd.n1126 gnd.n1125 585
R9378 gnd.n3157 gnd.n1126 585
R9379 gnd.n5017 gnd.n5016 585
R9380 gnd.n5016 gnd.n5015 585
R9381 gnd.n5018 gnd.n1120 585
R9382 gnd.n3149 gnd.n1120 585
R9383 gnd.n5020 gnd.n5019 585
R9384 gnd.n5021 gnd.n5020 585
R9385 gnd.n1104 gnd.n1103 585
R9386 gnd.n3141 gnd.n1104 585
R9387 gnd.n5029 gnd.n5028 585
R9388 gnd.n5028 gnd.n5027 585
R9389 gnd.n5030 gnd.n1098 585
R9390 gnd.n1105 gnd.n1098 585
R9391 gnd.n5032 gnd.n5031 585
R9392 gnd.n5033 gnd.n5032 585
R9393 gnd.n1085 gnd.n1084 585
R9394 gnd.n1088 gnd.n1085 585
R9395 gnd.n5041 gnd.n5040 585
R9396 gnd.n5040 gnd.n5039 585
R9397 gnd.n5042 gnd.n1079 585
R9398 gnd.n1079 gnd.n1077 585
R9399 gnd.n5044 gnd.n5043 585
R9400 gnd.n5045 gnd.n5044 585
R9401 gnd.n1080 gnd.n1078 585
R9402 gnd.n1078 gnd.n1065 585
R9403 gnd.n3088 gnd.n1066 585
R9404 gnd.n5051 gnd.n1066 585
R9405 gnd.n3024 gnd.n3022 585
R9406 gnd.n3022 gnd.n1063 585
R9407 gnd.n3093 gnd.n3092 585
R9408 gnd.n3100 gnd.n3093 585
R9409 gnd.n3023 gnd.n3021 585
R9410 gnd.n3021 gnd.n1009 585
R9411 gnd.n3084 gnd.n3083 585
R9412 gnd.n3082 gnd.n3081 585
R9413 gnd.n3080 gnd.n3079 585
R9414 gnd.n3078 gnd.n3077 585
R9415 gnd.n3076 gnd.n3075 585
R9416 gnd.n3074 gnd.n3073 585
R9417 gnd.n3072 gnd.n3071 585
R9418 gnd.n3070 gnd.n3069 585
R9419 gnd.n3068 gnd.n3067 585
R9420 gnd.n3066 gnd.n3065 585
R9421 gnd.n3064 gnd.n3063 585
R9422 gnd.n3062 gnd.n3061 585
R9423 gnd.n3060 gnd.n3059 585
R9424 gnd.n3058 gnd.n3057 585
R9425 gnd.n3056 gnd.n3055 585
R9426 gnd.n3054 gnd.n3053 585
R9427 gnd.n3052 gnd.n3051 585
R9428 gnd.n3043 gnd.n3040 585
R9429 gnd.n3047 gnd.n1008 585
R9430 gnd.n5138 gnd.n1008 585
R9431 gnd.n2793 gnd.n2792 585
R9432 gnd.n2790 gnd.n2784 585
R9433 gnd.n2800 gnd.n2781 585
R9434 gnd.n2801 gnd.n2779 585
R9435 gnd.n2778 gnd.n2771 585
R9436 gnd.n2808 gnd.n2770 585
R9437 gnd.n2809 gnd.n2769 585
R9438 gnd.n2767 gnd.n2759 585
R9439 gnd.n2816 gnd.n2758 585
R9440 gnd.n2817 gnd.n2756 585
R9441 gnd.n2755 gnd.n2748 585
R9442 gnd.n2824 gnd.n2747 585
R9443 gnd.n2825 gnd.n2746 585
R9444 gnd.n2744 gnd.n2737 585
R9445 gnd.n2832 gnd.n2736 585
R9446 gnd.n2833 gnd.n2734 585
R9447 gnd.n2733 gnd.n2729 585
R9448 gnd.n2731 gnd.n2730 585
R9449 gnd.n1326 gnd.n1324 585
R9450 gnd.n2606 gnd.n1324 585
R9451 gnd.n2643 gnd.n1322 585
R9452 gnd.n4900 gnd.n1322 585
R9453 gnd.n3449 gnd.n3448 585
R9454 gnd.n3450 gnd.n3449 585
R9455 gnd.n2642 gnd.n1313 585
R9456 gnd.n4906 gnd.n1313 585
R9457 gnd.n3287 gnd.n3286 585
R9458 gnd.n3286 gnd.n3285 585
R9459 gnd.n2865 gnd.n1302 585
R9460 gnd.n4912 gnd.n1302 585
R9461 gnd.n3291 gnd.n2864 585
R9462 gnd.n3276 gnd.n2864 585
R9463 gnd.n3292 gnd.n1291 585
R9464 gnd.n4918 gnd.n1291 585
R9465 gnd.n3293 gnd.n2863 585
R9466 gnd.n3272 gnd.n2863 585
R9467 gnd.n2860 gnd.n1280 585
R9468 gnd.n4924 gnd.n1280 585
R9469 gnd.n3298 gnd.n3297 585
R9470 gnd.n3299 gnd.n3298 585
R9471 gnd.n2859 gnd.n1270 585
R9472 gnd.n4930 gnd.n1270 585
R9473 gnd.n3263 gnd.n3262 585
R9474 gnd.n3264 gnd.n3263 585
R9475 gnd.n2873 gnd.n1260 585
R9476 gnd.n4936 gnd.n1260 585
R9477 gnd.n3258 gnd.n3257 585
R9478 gnd.n3257 gnd.n3256 585
R9479 gnd.n2875 gnd.n1249 585
R9480 gnd.n4942 gnd.n1249 585
R9481 gnd.n3246 gnd.n3245 585
R9482 gnd.n3247 gnd.n3246 585
R9483 gnd.n2879 gnd.n1238 585
R9484 gnd.n4948 gnd.n1238 585
R9485 gnd.n3241 gnd.n3240 585
R9486 gnd.n3240 gnd.n3239 585
R9487 gnd.n2881 gnd.n1228 585
R9488 gnd.n4954 gnd.n1228 585
R9489 gnd.n3230 gnd.n3229 585
R9490 gnd.n3231 gnd.n3230 585
R9491 gnd.n2887 gnd.n1218 585
R9492 gnd.n4960 gnd.n1218 585
R9493 gnd.n3225 gnd.n3224 585
R9494 gnd.n3224 gnd.n3223 585
R9495 gnd.n2889 gnd.n1208 585
R9496 gnd.n4966 gnd.n1208 585
R9497 gnd.n3214 gnd.n3213 585
R9498 gnd.n3215 gnd.n3214 585
R9499 gnd.n2893 gnd.n1197 585
R9500 gnd.n4972 gnd.n1197 585
R9501 gnd.n3209 gnd.n3208 585
R9502 gnd.n3208 gnd.n3207 585
R9503 gnd.n2895 gnd.n1190 585
R9504 gnd.n4979 gnd.n1190 585
R9505 gnd.n3197 gnd.n3196 585
R9506 gnd.n3198 gnd.n3197 585
R9507 gnd.n2902 gnd.n1180 585
R9508 gnd.n4985 gnd.n1180 585
R9509 gnd.n3191 gnd.n3190 585
R9510 gnd.n3190 gnd.n3189 585
R9511 gnd.n2904 gnd.n1171 585
R9512 gnd.n4991 gnd.n1171 585
R9513 gnd.n3180 gnd.n3179 585
R9514 gnd.n3181 gnd.n3180 585
R9515 gnd.n2908 gnd.n1160 585
R9516 gnd.n4997 gnd.n1160 585
R9517 gnd.n3175 gnd.n3174 585
R9518 gnd.n3174 gnd.n3173 585
R9519 gnd.n2910 gnd.n1150 585
R9520 gnd.n5003 gnd.n1150 585
R9521 gnd.n3164 gnd.n3163 585
R9522 gnd.n3165 gnd.n3164 585
R9523 gnd.n3006 gnd.n1140 585
R9524 gnd.n5009 gnd.n1140 585
R9525 gnd.n3159 gnd.n3158 585
R9526 gnd.n3158 gnd.n3157 585
R9527 gnd.n3008 gnd.n1129 585
R9528 gnd.n5015 gnd.n1129 585
R9529 gnd.n3148 gnd.n3147 585
R9530 gnd.n3149 gnd.n3148 585
R9531 gnd.n3012 gnd.n1118 585
R9532 gnd.n5021 gnd.n1118 585
R9533 gnd.n3143 gnd.n3142 585
R9534 gnd.n3142 gnd.n3141 585
R9535 gnd.n3120 gnd.n1107 585
R9536 gnd.n5027 gnd.n1107 585
R9537 gnd.n3119 gnd.n3118 585
R9538 gnd.n3118 gnd.n1105 585
R9539 gnd.n3014 gnd.n1097 585
R9540 gnd.n5033 gnd.n1097 585
R9541 gnd.n3114 gnd.n3113 585
R9542 gnd.n3113 gnd.n1088 585
R9543 gnd.n3112 gnd.n1087 585
R9544 gnd.n5039 gnd.n1087 585
R9545 gnd.n3111 gnd.n3110 585
R9546 gnd.n3110 gnd.n1077 585
R9547 gnd.n3016 gnd.n1076 585
R9548 gnd.n5045 gnd.n1076 585
R9549 gnd.n3106 gnd.n3105 585
R9550 gnd.n3105 gnd.n1065 585
R9551 gnd.n3104 gnd.n1064 585
R9552 gnd.n5051 gnd.n1064 585
R9553 gnd.n3103 gnd.n3102 585
R9554 gnd.n3102 gnd.n1063 585
R9555 gnd.n3101 gnd.n3018 585
R9556 gnd.n3101 gnd.n3100 585
R9557 gnd.n3045 gnd.n3020 585
R9558 gnd.n3020 gnd.n1009 585
R9559 gnd.n7647 gnd.n107 585
R9560 gnd.n7743 gnd.n107 585
R9561 gnd.n7648 gnd.n7578 585
R9562 gnd.n7578 gnd.n104 585
R9563 gnd.n7649 gnd.n187 585
R9564 gnd.n7663 gnd.n187 585
R9565 gnd.n198 gnd.n196 585
R9566 gnd.n196 gnd.n186 585
R9567 gnd.n7654 gnd.n7653 585
R9568 gnd.n7655 gnd.n7654 585
R9569 gnd.n197 gnd.n195 585
R9570 gnd.n195 gnd.n193 585
R9571 gnd.n7574 gnd.n7573 585
R9572 gnd.n7573 gnd.n7572 585
R9573 gnd.n201 gnd.n200 585
R9574 gnd.n211 gnd.n201 585
R9575 gnd.n7563 gnd.n7562 585
R9576 gnd.n7564 gnd.n7563 585
R9577 gnd.n213 gnd.n212 585
R9578 gnd.n212 gnd.n208 585
R9579 gnd.n7558 gnd.n7557 585
R9580 gnd.n7557 gnd.n7556 585
R9581 gnd.n216 gnd.n215 585
R9582 gnd.n218 gnd.n216 585
R9583 gnd.n7547 gnd.n7546 585
R9584 gnd.n7548 gnd.n7547 585
R9585 gnd.n228 gnd.n227 585
R9586 gnd.n7450 gnd.n227 585
R9587 gnd.n7542 gnd.n7541 585
R9588 gnd.n7541 gnd.n7540 585
R9589 gnd.n231 gnd.n230 585
R9590 gnd.n7457 gnd.n231 585
R9591 gnd.n7531 gnd.n7530 585
R9592 gnd.n7532 gnd.n7531 585
R9593 gnd.n243 gnd.n242 585
R9594 gnd.n7417 gnd.n242 585
R9595 gnd.n7526 gnd.n7525 585
R9596 gnd.n7525 gnd.n7524 585
R9597 gnd.n246 gnd.n245 585
R9598 gnd.n7413 gnd.n246 585
R9599 gnd.n7515 gnd.n7514 585
R9600 gnd.n7516 gnd.n7515 585
R9601 gnd.n259 gnd.n258 585
R9602 gnd.n7406 gnd.n258 585
R9603 gnd.n7510 gnd.n7509 585
R9604 gnd.n7509 gnd.n7508 585
R9605 gnd.n262 gnd.n261 585
R9606 gnd.n7474 gnd.n262 585
R9607 gnd.n7487 gnd.n7486 585
R9608 gnd.n7486 gnd.n7485 585
R9609 gnd.n7488 gnd.n293 585
R9610 gnd.n7480 gnd.n293 585
R9611 gnd.n4647 gnd.n290 585
R9612 gnd.n4648 gnd.n4647 585
R9613 gnd.n7493 gnd.n289 585
R9614 gnd.n4660 gnd.n289 585
R9615 gnd.n7494 gnd.n288 585
R9616 gnd.n4664 gnd.n288 585
R9617 gnd.n7495 gnd.n287 585
R9618 gnd.n1541 gnd.n287 585
R9619 gnd.n284 gnd.n282 585
R9620 gnd.n4637 gnd.n282 585
R9621 gnd.n7500 gnd.n7499 585
R9622 gnd.n7501 gnd.n7500 585
R9623 gnd.n283 gnd.n281 585
R9624 gnd.n4625 gnd.n281 585
R9625 gnd.n4689 gnd.n4688 585
R9626 gnd.n4688 gnd.n4687 585
R9627 gnd.n4692 gnd.n1517 585
R9628 gnd.n1528 gnd.n1517 585
R9629 gnd.n4693 gnd.n1516 585
R9630 gnd.n4679 gnd.n1516 585
R9631 gnd.n4694 gnd.n1515 585
R9632 gnd.n4612 gnd.n1515 585
R9633 gnd.n1571 gnd.n1513 585
R9634 gnd.n1572 gnd.n1571 585
R9635 gnd.n4698 gnd.n1512 585
R9636 gnd.n4599 gnd.n1512 585
R9637 gnd.n4699 gnd.n1511 585
R9638 gnd.n1581 gnd.n1511 585
R9639 gnd.n4700 gnd.n1510 585
R9640 gnd.n4589 gnd.n1510 585
R9641 gnd.n4569 gnd.n1508 585
R9642 gnd.n4570 gnd.n4569 585
R9643 gnd.n4704 gnd.n1507 585
R9644 gnd.n1589 gnd.n1507 585
R9645 gnd.n4705 gnd.n1506 585
R9646 gnd.n4560 gnd.n1506 585
R9647 gnd.n4706 gnd.n1505 585
R9648 gnd.n1608 gnd.n1505 585
R9649 gnd.n4549 gnd.n1503 585
R9650 gnd.n4550 gnd.n4549 585
R9651 gnd.n4710 gnd.n1502 585
R9652 gnd.n4537 gnd.n1502 585
R9653 gnd.n4711 gnd.n1501 585
R9654 gnd.n1616 gnd.n1501 585
R9655 gnd.n4712 gnd.n1500 585
R9656 gnd.n4528 gnd.n1500 585
R9657 gnd.n1497 gnd.n1495 585
R9658 gnd.n1635 gnd.n1495 585
R9659 gnd.n4717 gnd.n4716 585
R9660 gnd.n4718 gnd.n4717 585
R9661 gnd.n1496 gnd.n1494 585
R9662 gnd.n4487 gnd.n1494 585
R9663 gnd.n1689 gnd.n1481 585
R9664 gnd.n4724 gnd.n1481 585
R9665 gnd.n1690 gnd.n1688 585
R9666 gnd.n1688 gnd.n1477 585
R9667 gnd.n1687 gnd.n1684 585
R9668 gnd.n1683 gnd.n1682 585
R9669 gnd.n1705 gnd.n1704 585
R9670 gnd.n1707 gnd.n1681 585
R9671 gnd.n1710 gnd.n1709 585
R9672 gnd.n1674 gnd.n1673 585
R9673 gnd.n1724 gnd.n1723 585
R9674 gnd.n1726 gnd.n1672 585
R9675 gnd.n1729 gnd.n1728 585
R9676 gnd.n1665 gnd.n1664 585
R9677 gnd.n1743 gnd.n1742 585
R9678 gnd.n1745 gnd.n1663 585
R9679 gnd.n1748 gnd.n1747 585
R9680 gnd.n1656 gnd.n1655 585
R9681 gnd.n1762 gnd.n1761 585
R9682 gnd.n1764 gnd.n1654 585
R9683 gnd.n1767 gnd.n1766 585
R9684 gnd.n1647 gnd.n1644 585
R9685 gnd.n4478 gnd.n4477 585
R9686 gnd.n4478 gnd.n1468 585
R9687 gnd.n7618 gnd.n103 585
R9688 gnd.n7619 gnd.n7616 585
R9689 gnd.n7620 gnd.n7612 585
R9690 gnd.n7610 gnd.n7608 585
R9691 gnd.n7624 gnd.n7607 585
R9692 gnd.n7625 gnd.n7605 585
R9693 gnd.n7626 gnd.n7604 585
R9694 gnd.n7602 gnd.n7600 585
R9695 gnd.n7630 gnd.n7599 585
R9696 gnd.n7631 gnd.n7597 585
R9697 gnd.n7632 gnd.n7596 585
R9698 gnd.n7594 gnd.n7592 585
R9699 gnd.n7636 gnd.n7591 585
R9700 gnd.n7637 gnd.n7589 585
R9701 gnd.n7638 gnd.n7588 585
R9702 gnd.n7586 gnd.n7584 585
R9703 gnd.n7642 gnd.n7583 585
R9704 gnd.n7643 gnd.n7581 585
R9705 gnd.n7644 gnd.n7580 585
R9706 gnd.n7580 gnd.n117 585
R9707 gnd.n7745 gnd.n7744 585
R9708 gnd.n7744 gnd.n7743 585
R9709 gnd.n7746 gnd.n101 585
R9710 gnd.n104 gnd.n101 585
R9711 gnd.n7747 gnd.n100 585
R9712 gnd.n7663 gnd.n100 585
R9713 gnd.n185 gnd.n98 585
R9714 gnd.n186 gnd.n185 585
R9715 gnd.n7751 gnd.n97 585
R9716 gnd.n7655 gnd.n97 585
R9717 gnd.n7752 gnd.n96 585
R9718 gnd.n193 gnd.n96 585
R9719 gnd.n7753 gnd.n95 585
R9720 gnd.n7572 gnd.n95 585
R9721 gnd.n210 gnd.n93 585
R9722 gnd.n211 gnd.n210 585
R9723 gnd.n7757 gnd.n92 585
R9724 gnd.n7564 gnd.n92 585
R9725 gnd.n7758 gnd.n91 585
R9726 gnd.n208 gnd.n91 585
R9727 gnd.n7759 gnd.n90 585
R9728 gnd.n7556 gnd.n90 585
R9729 gnd.n217 gnd.n88 585
R9730 gnd.n218 gnd.n217 585
R9731 gnd.n7763 gnd.n87 585
R9732 gnd.n7548 gnd.n87 585
R9733 gnd.n7764 gnd.n86 585
R9734 gnd.n7450 gnd.n86 585
R9735 gnd.n7765 gnd.n85 585
R9736 gnd.n7540 gnd.n85 585
R9737 gnd.n7456 gnd.n83 585
R9738 gnd.n7457 gnd.n7456 585
R9739 gnd.n7769 gnd.n82 585
R9740 gnd.n7532 gnd.n82 585
R9741 gnd.n7770 gnd.n81 585
R9742 gnd.n7417 gnd.n81 585
R9743 gnd.n7771 gnd.n80 585
R9744 gnd.n7524 gnd.n80 585
R9745 gnd.n7412 gnd.n78 585
R9746 gnd.n7413 gnd.n7412 585
R9747 gnd.n7775 gnd.n77 585
R9748 gnd.n7516 gnd.n77 585
R9749 gnd.n7776 gnd.n76 585
R9750 gnd.n7406 gnd.n76 585
R9751 gnd.n7777 gnd.n75 585
R9752 gnd.n7508 gnd.n75 585
R9753 gnd.n305 gnd.n73 585
R9754 gnd.n7474 gnd.n305 585
R9755 gnd.n7781 gnd.n72 585
R9756 gnd.n7485 gnd.n72 585
R9757 gnd.n7782 gnd.n71 585
R9758 gnd.n7480 gnd.n71 585
R9759 gnd.n7783 gnd.n70 585
R9760 gnd.n4648 gnd.n70 585
R9761 gnd.n4646 gnd.n69 585
R9762 gnd.n4660 gnd.n4646 585
R9763 gnd.n4630 gnd.n1543 585
R9764 gnd.n4664 gnd.n1543 585
R9765 gnd.n1553 gnd.n1551 585
R9766 gnd.n1551 gnd.n1541 585
R9767 gnd.n4635 gnd.n4634 585
R9768 gnd.n4637 gnd.n4635 585
R9769 gnd.n1552 gnd.n279 585
R9770 gnd.n7501 gnd.n279 585
R9771 gnd.n4627 gnd.n4626 585
R9772 gnd.n4626 gnd.n4625 585
R9773 gnd.n1555 gnd.n1519 585
R9774 gnd.n4687 gnd.n1519 585
R9775 gnd.n4605 gnd.n4604 585
R9776 gnd.n4604 gnd.n1528 585
R9777 gnd.n1564 gnd.n1527 585
R9778 gnd.n4679 gnd.n1527 585
R9779 gnd.n4610 gnd.n4609 585
R9780 gnd.n4612 gnd.n4610 585
R9781 gnd.n1563 gnd.n1562 585
R9782 gnd.n1572 gnd.n1562 585
R9783 gnd.n4601 gnd.n4600 585
R9784 gnd.n4600 gnd.n4599 585
R9785 gnd.n1567 gnd.n1566 585
R9786 gnd.n1581 gnd.n1567 585
R9787 gnd.n1593 gnd.n1580 585
R9788 gnd.n4589 gnd.n1580 585
R9789 gnd.n4568 gnd.n4567 585
R9790 gnd.n4570 gnd.n4568 585
R9791 gnd.n1592 gnd.n1591 585
R9792 gnd.n1591 gnd.n1589 585
R9793 gnd.n4562 gnd.n4561 585
R9794 gnd.n4561 gnd.n4560 585
R9795 gnd.n1596 gnd.n1595 585
R9796 gnd.n1608 gnd.n1596 585
R9797 gnd.n1620 gnd.n1607 585
R9798 gnd.n4550 gnd.n1607 585
R9799 gnd.n4536 gnd.n4535 585
R9800 gnd.n4537 gnd.n4536 585
R9801 gnd.n1619 gnd.n1618 585
R9802 gnd.n1618 gnd.n1616 585
R9803 gnd.n4530 gnd.n4529 585
R9804 gnd.n4529 gnd.n4528 585
R9805 gnd.n1623 gnd.n1622 585
R9806 gnd.n1635 gnd.n1623 585
R9807 gnd.n1642 gnd.n1492 585
R9808 gnd.n4718 gnd.n1492 585
R9809 gnd.n4486 gnd.n4485 585
R9810 gnd.n4487 gnd.n4486 585
R9811 gnd.n1641 gnd.n1479 585
R9812 gnd.n4724 gnd.n1479 585
R9813 gnd.n4480 gnd.n4479 585
R9814 gnd.n4479 gnd.n1477 585
R9815 gnd.n953 gnd.n952 585
R9816 gnd.n956 gnd.n953 585
R9817 gnd.n6501 gnd.n6500 585
R9818 gnd.n6500 gnd.n6499 585
R9819 gnd.n6502 gnd.n947 585
R9820 gnd.n6398 gnd.n947 585
R9821 gnd.n6504 gnd.n6503 585
R9822 gnd.n6505 gnd.n6504 585
R9823 gnd.n948 gnd.n946 585
R9824 gnd.n946 gnd.n942 585
R9825 gnd.n928 gnd.n927 585
R9826 gnd.n931 gnd.n928 585
R9827 gnd.n6515 gnd.n6514 585
R9828 gnd.n6514 gnd.n6513 585
R9829 gnd.n6516 gnd.n922 585
R9830 gnd.n6119 gnd.n922 585
R9831 gnd.n6518 gnd.n6517 585
R9832 gnd.n6519 gnd.n6518 585
R9833 gnd.n923 gnd.n921 585
R9834 gnd.n6103 gnd.n921 585
R9835 gnd.n6094 gnd.n6093 585
R9836 gnd.n6093 gnd.n909 585
R9837 gnd.n6092 gnd.n5211 585
R9838 gnd.n6092 gnd.n907 585
R9839 gnd.n6091 gnd.n5213 585
R9840 gnd.n6091 gnd.n6090 585
R9841 gnd.n6081 gnd.n5212 585
R9842 gnd.n5224 gnd.n5212 585
R9843 gnd.n6080 gnd.n6079 585
R9844 gnd.n6079 gnd.n6078 585
R9845 gnd.n5221 gnd.n5219 585
R9846 gnd.n6065 gnd.n5221 585
R9847 gnd.n6056 gnd.n6055 585
R9848 gnd.n6055 gnd.n6054 585
R9849 gnd.n5236 gnd.n5235 585
R9850 gnd.n5244 gnd.n5236 585
R9851 gnd.n6033 gnd.n6032 585
R9852 gnd.n6034 gnd.n6033 585
R9853 gnd.n5247 gnd.n5246 585
R9854 gnd.n5255 gnd.n5246 585
R9855 gnd.n6007 gnd.n5267 585
R9856 gnd.n5267 gnd.n5254 585
R9857 gnd.n6009 gnd.n6008 585
R9858 gnd.n6010 gnd.n6009 585
R9859 gnd.n5268 gnd.n5266 585
R9860 gnd.n5266 gnd.n5262 585
R9861 gnd.n5996 gnd.n5995 585
R9862 gnd.n5995 gnd.n5994 585
R9863 gnd.n5273 gnd.n5272 585
R9864 gnd.n5283 gnd.n5273 585
R9865 gnd.n5985 gnd.n5984 585
R9866 gnd.n5984 gnd.n5983 585
R9867 gnd.n5280 gnd.n5279 585
R9868 gnd.n5971 gnd.n5280 585
R9869 gnd.n5945 gnd.n5349 585
R9870 gnd.n5349 gnd.n5290 585
R9871 gnd.n5947 gnd.n5946 585
R9872 gnd.n5948 gnd.n5947 585
R9873 gnd.n5350 gnd.n5348 585
R9874 gnd.n5358 gnd.n5348 585
R9875 gnd.n5923 gnd.n5370 585
R9876 gnd.n5370 gnd.n5357 585
R9877 gnd.n5925 gnd.n5924 585
R9878 gnd.n5926 gnd.n5925 585
R9879 gnd.n5371 gnd.n5369 585
R9880 gnd.n5369 gnd.n5365 585
R9881 gnd.n5911 gnd.n5910 585
R9882 gnd.n5910 gnd.n5909 585
R9883 gnd.n5376 gnd.n5375 585
R9884 gnd.n5385 gnd.n5376 585
R9885 gnd.n5900 gnd.n5899 585
R9886 gnd.n5899 gnd.n5898 585
R9887 gnd.n5383 gnd.n5382 585
R9888 gnd.n5886 gnd.n5383 585
R9889 gnd.n5858 gnd.n5857 585
R9890 gnd.n5857 gnd.n5392 585
R9891 gnd.n5859 gnd.n5403 585
R9892 gnd.n5850 gnd.n5403 585
R9893 gnd.n5861 gnd.n5860 585
R9894 gnd.n5862 gnd.n5861 585
R9895 gnd.n5404 gnd.n5402 585
R9896 gnd.n5418 gnd.n5402 585
R9897 gnd.n5842 gnd.n5841 585
R9898 gnd.n5841 gnd.n5840 585
R9899 gnd.n5415 gnd.n5414 585
R9900 gnd.n5825 gnd.n5415 585
R9901 gnd.n5812 gnd.n5435 585
R9902 gnd.n5435 gnd.n5425 585
R9903 gnd.n5814 gnd.n5813 585
R9904 gnd.n5815 gnd.n5814 585
R9905 gnd.n5436 gnd.n5434 585
R9906 gnd.n5444 gnd.n5434 585
R9907 gnd.n5788 gnd.n5456 585
R9908 gnd.n5456 gnd.n5443 585
R9909 gnd.n5790 gnd.n5789 585
R9910 gnd.n5791 gnd.n5790 585
R9911 gnd.n5457 gnd.n5455 585
R9912 gnd.n5455 gnd.n5451 585
R9913 gnd.n5776 gnd.n5775 585
R9914 gnd.n5775 gnd.n5774 585
R9915 gnd.n5462 gnd.n5461 585
R9916 gnd.n5466 gnd.n5462 585
R9917 gnd.n5760 gnd.n5759 585
R9918 gnd.n5761 gnd.n5760 585
R9919 gnd.n5477 gnd.n5476 585
R9920 gnd.n5476 gnd.n5472 585
R9921 gnd.n5750 gnd.n5749 585
R9922 gnd.n5751 gnd.n5750 585
R9923 gnd.n5486 gnd.n5485 585
R9924 gnd.n5485 gnd.n5483 585
R9925 gnd.n5744 gnd.n5743 585
R9926 gnd.n5743 gnd.n5742 585
R9927 gnd.n5490 gnd.n5489 585
R9928 gnd.n5498 gnd.n5490 585
R9929 gnd.n5651 gnd.n5650 585
R9930 gnd.n5652 gnd.n5651 585
R9931 gnd.n5500 gnd.n5499 585
R9932 gnd.n5499 gnd.n5497 585
R9933 gnd.n5646 gnd.n5645 585
R9934 gnd.n5645 gnd.n5644 585
R9935 gnd.n5503 gnd.n5502 585
R9936 gnd.n5504 gnd.n5503 585
R9937 gnd.n5635 gnd.n5634 585
R9938 gnd.n5636 gnd.n5635 585
R9939 gnd.n5512 gnd.n5511 585
R9940 gnd.n5511 gnd.n5510 585
R9941 gnd.n5630 gnd.n5629 585
R9942 gnd.n5629 gnd.n5628 585
R9943 gnd.n5515 gnd.n5514 585
R9944 gnd.n5516 gnd.n5515 585
R9945 gnd.n5619 gnd.n5618 585
R9946 gnd.n5620 gnd.n5619 585
R9947 gnd.n5615 gnd.n5522 585
R9948 gnd.n5614 gnd.n5613 585
R9949 gnd.n5611 gnd.n5524 585
R9950 gnd.n5611 gnd.n5521 585
R9951 gnd.n5610 gnd.n5609 585
R9952 gnd.n5608 gnd.n5607 585
R9953 gnd.n5606 gnd.n5529 585
R9954 gnd.n5604 gnd.n5603 585
R9955 gnd.n5602 gnd.n5530 585
R9956 gnd.n5601 gnd.n5600 585
R9957 gnd.n5598 gnd.n5535 585
R9958 gnd.n5596 gnd.n5595 585
R9959 gnd.n5594 gnd.n5536 585
R9960 gnd.n5593 gnd.n5592 585
R9961 gnd.n5590 gnd.n5541 585
R9962 gnd.n5588 gnd.n5587 585
R9963 gnd.n5586 gnd.n5542 585
R9964 gnd.n5585 gnd.n5584 585
R9965 gnd.n5582 gnd.n5547 585
R9966 gnd.n5580 gnd.n5579 585
R9967 gnd.n5578 gnd.n5548 585
R9968 gnd.n5577 gnd.n5576 585
R9969 gnd.n5574 gnd.n5553 585
R9970 gnd.n5572 gnd.n5571 585
R9971 gnd.n5569 gnd.n5554 585
R9972 gnd.n5568 gnd.n5567 585
R9973 gnd.n5565 gnd.n5563 585
R9974 gnd.n5561 gnd.n5520 585
R9975 gnd.n6407 gnd.n6406 585
R9976 gnd.n6409 gnd.n6408 585
R9977 gnd.n6411 gnd.n6410 585
R9978 gnd.n6413 gnd.n6412 585
R9979 gnd.n6415 gnd.n6414 585
R9980 gnd.n6417 gnd.n6416 585
R9981 gnd.n6419 gnd.n6418 585
R9982 gnd.n6421 gnd.n6420 585
R9983 gnd.n6423 gnd.n6422 585
R9984 gnd.n6425 gnd.n6424 585
R9985 gnd.n6427 gnd.n6426 585
R9986 gnd.n6429 gnd.n6428 585
R9987 gnd.n6431 gnd.n6430 585
R9988 gnd.n6433 gnd.n6432 585
R9989 gnd.n6435 gnd.n6434 585
R9990 gnd.n6437 gnd.n6436 585
R9991 gnd.n6439 gnd.n6438 585
R9992 gnd.n6441 gnd.n6440 585
R9993 gnd.n6443 gnd.n6442 585
R9994 gnd.n6445 gnd.n6444 585
R9995 gnd.n6447 gnd.n6446 585
R9996 gnd.n6449 gnd.n6448 585
R9997 gnd.n6451 gnd.n6450 585
R9998 gnd.n6453 gnd.n6452 585
R9999 gnd.n6455 gnd.n6454 585
R10000 gnd.n6456 gnd.n5165 585
R10001 gnd.n6457 gnd.n967 585
R10002 gnd.n6490 gnd.n967 585
R10003 gnd.n6405 gnd.n6404 585
R10004 gnd.n6405 gnd.n956 585
R10005 gnd.n5194 gnd.n954 585
R10006 gnd.n6499 gnd.n954 585
R10007 gnd.n6400 gnd.n6399 585
R10008 gnd.n6399 gnd.n6398 585
R10009 gnd.n5196 gnd.n944 585
R10010 gnd.n6505 gnd.n944 585
R10011 gnd.n6113 gnd.n6112 585
R10012 gnd.n6113 gnd.n942 585
R10013 gnd.n6115 gnd.n6114 585
R10014 gnd.n6114 gnd.n931 585
R10015 gnd.n6116 gnd.n929 585
R10016 gnd.n6513 gnd.n929 585
R10017 gnd.n6118 gnd.n6117 585
R10018 gnd.n6119 gnd.n6118 585
R10019 gnd.n5205 gnd.n919 585
R10020 gnd.n6519 gnd.n919 585
R10021 gnd.n6105 gnd.n6104 585
R10022 gnd.n6104 gnd.n6103 585
R10023 gnd.n5208 gnd.n5207 585
R10024 gnd.n5208 gnd.n909 585
R10025 gnd.n6046 gnd.n6045 585
R10026 gnd.n6045 gnd.n907 585
R10027 gnd.n6047 gnd.n5215 585
R10028 gnd.n6090 gnd.n5215 585
R10029 gnd.n6049 gnd.n6048 585
R10030 gnd.n6048 gnd.n5224 585
R10031 gnd.n6050 gnd.n5222 585
R10032 gnd.n6078 gnd.n5222 585
R10033 gnd.n6051 gnd.n5232 585
R10034 gnd.n6065 gnd.n5232 585
R10035 gnd.n6053 gnd.n6052 585
R10036 gnd.n6054 gnd.n6053 585
R10037 gnd.n5239 gnd.n5238 585
R10038 gnd.n5244 gnd.n5238 585
R10039 gnd.n6036 gnd.n6035 585
R10040 gnd.n6035 gnd.n6034 585
R10041 gnd.n5242 gnd.n5241 585
R10042 gnd.n5255 gnd.n5242 585
R10043 gnd.n5961 gnd.n5960 585
R10044 gnd.n5960 gnd.n5254 585
R10045 gnd.n5962 gnd.n5264 585
R10046 gnd.n6010 gnd.n5264 585
R10047 gnd.n5964 gnd.n5963 585
R10048 gnd.n5963 gnd.n5262 585
R10049 gnd.n5965 gnd.n5275 585
R10050 gnd.n5994 gnd.n5275 585
R10051 gnd.n5967 gnd.n5966 585
R10052 gnd.n5966 gnd.n5283 585
R10053 gnd.n5968 gnd.n5282 585
R10054 gnd.n5983 gnd.n5282 585
R10055 gnd.n5970 gnd.n5969 585
R10056 gnd.n5971 gnd.n5970 585
R10057 gnd.n5294 gnd.n5293 585
R10058 gnd.n5293 gnd.n5290 585
R10059 gnd.n5950 gnd.n5949 585
R10060 gnd.n5949 gnd.n5948 585
R10061 gnd.n5345 gnd.n5344 585
R10062 gnd.n5358 gnd.n5345 585
R10063 gnd.n5871 gnd.n5870 585
R10064 gnd.n5870 gnd.n5357 585
R10065 gnd.n5872 gnd.n5367 585
R10066 gnd.n5926 gnd.n5367 585
R10067 gnd.n5875 gnd.n5874 585
R10068 gnd.n5874 gnd.n5365 585
R10069 gnd.n5876 gnd.n5378 585
R10070 gnd.n5909 gnd.n5378 585
R10071 gnd.n5879 gnd.n5878 585
R10072 gnd.n5878 gnd.n5385 585
R10073 gnd.n5880 gnd.n5384 585
R10074 gnd.n5898 gnd.n5384 585
R10075 gnd.n5883 gnd.n5882 585
R10076 gnd.n5886 gnd.n5883 585
R10077 gnd.n5868 gnd.n5394 585
R10078 gnd.n5394 gnd.n5392 585
R10079 gnd.n5399 gnd.n5395 585
R10080 gnd.n5850 gnd.n5399 585
R10081 gnd.n5864 gnd.n5863 585
R10082 gnd.n5863 gnd.n5862 585
R10083 gnd.n5398 gnd.n5397 585
R10084 gnd.n5418 gnd.n5398 585
R10085 gnd.n5822 gnd.n5417 585
R10086 gnd.n5840 gnd.n5417 585
R10087 gnd.n5824 gnd.n5823 585
R10088 gnd.n5825 gnd.n5824 585
R10089 gnd.n5428 gnd.n5427 585
R10090 gnd.n5427 gnd.n5425 585
R10091 gnd.n5817 gnd.n5816 585
R10092 gnd.n5816 gnd.n5815 585
R10093 gnd.n5431 gnd.n5430 585
R10094 gnd.n5444 gnd.n5431 585
R10095 gnd.n5668 gnd.n5667 585
R10096 gnd.n5667 gnd.n5443 585
R10097 gnd.n5669 gnd.n5453 585
R10098 gnd.n5791 gnd.n5453 585
R10099 gnd.n5671 gnd.n5670 585
R10100 gnd.n5670 gnd.n5451 585
R10101 gnd.n5672 gnd.n5463 585
R10102 gnd.n5774 gnd.n5463 585
R10103 gnd.n5674 gnd.n5673 585
R10104 gnd.n5673 gnd.n5466 585
R10105 gnd.n5675 gnd.n5474 585
R10106 gnd.n5761 gnd.n5474 585
R10107 gnd.n5677 gnd.n5676 585
R10108 gnd.n5676 gnd.n5472 585
R10109 gnd.n5678 gnd.n5484 585
R10110 gnd.n5751 gnd.n5484 585
R10111 gnd.n5679 gnd.n5492 585
R10112 gnd.n5492 gnd.n5483 585
R10113 gnd.n5681 gnd.n5680 585
R10114 gnd.n5742 gnd.n5681 585
R10115 gnd.n5493 gnd.n5491 585
R10116 gnd.n5498 gnd.n5491 585
R10117 gnd.n5654 gnd.n5653 585
R10118 gnd.n5653 gnd.n5652 585
R10119 gnd.n5496 gnd.n5495 585
R10120 gnd.n5497 gnd.n5496 585
R10121 gnd.n5643 gnd.n5642 585
R10122 gnd.n5644 gnd.n5643 585
R10123 gnd.n5506 gnd.n5505 585
R10124 gnd.n5505 gnd.n5504 585
R10125 gnd.n5638 gnd.n5637 585
R10126 gnd.n5637 gnd.n5636 585
R10127 gnd.n5509 gnd.n5508 585
R10128 gnd.n5510 gnd.n5509 585
R10129 gnd.n5627 gnd.n5626 585
R10130 gnd.n5628 gnd.n5627 585
R10131 gnd.n5518 gnd.n5517 585
R10132 gnd.n5517 gnd.n5516 585
R10133 gnd.n5622 gnd.n5621 585
R10134 gnd.n5621 gnd.n5620 585
R10135 gnd.n6495 gnd.n958 585
R10136 gnd.n966 gnd.n958 585
R10137 gnd.n6497 gnd.n6496 585
R10138 gnd.n6498 gnd.n6497 585
R10139 gnd.n959 gnd.n957 585
R10140 gnd.n6397 gnd.n957 585
R10141 gnd.n941 gnd.n940 585
R10142 gnd.n945 gnd.n941 585
R10143 gnd.n6508 gnd.n6507 585
R10144 gnd.n6507 gnd.n6506 585
R10145 gnd.n6509 gnd.n933 585
R10146 gnd.n5198 gnd.n933 585
R10147 gnd.n6511 gnd.n6510 585
R10148 gnd.n6512 gnd.n6511 585
R10149 gnd.n934 gnd.n932 585
R10150 gnd.n6120 gnd.n932 585
R10151 gnd.n917 gnd.n916 585
R10152 gnd.n920 gnd.n917 585
R10153 gnd.n6522 gnd.n6521 585
R10154 gnd.n6521 gnd.n6520 585
R10155 gnd.n6523 gnd.n911 585
R10156 gnd.n6102 gnd.n911 585
R10157 gnd.n6525 gnd.n6524 585
R10158 gnd.n6526 gnd.n6525 585
R10159 gnd.n912 gnd.n910 585
R10160 gnd.n6089 gnd.n910 585
R10161 gnd.n6074 gnd.n5226 585
R10162 gnd.n5226 gnd.n5214 585
R10163 gnd.n6076 gnd.n6075 585
R10164 gnd.n6077 gnd.n6076 585
R10165 gnd.n5227 gnd.n5225 585
R10166 gnd.n6064 gnd.n5225 585
R10167 gnd.n6068 gnd.n6067 585
R10168 gnd.n6067 gnd.n6066 585
R10169 gnd.n5230 gnd.n5229 585
R10170 gnd.n5237 gnd.n5230 585
R10171 gnd.n6020 gnd.n6019 585
R10172 gnd.n6019 gnd.n5245 585
R10173 gnd.n6021 gnd.n5257 585
R10174 gnd.n5257 gnd.n5243 585
R10175 gnd.n6023 gnd.n6022 585
R10176 gnd.n6024 gnd.n6023 585
R10177 gnd.n5258 gnd.n5256 585
R10178 gnd.n5265 gnd.n5256 585
R10179 gnd.n6013 gnd.n6012 585
R10180 gnd.n6012 gnd.n6011 585
R10181 gnd.n5261 gnd.n5260 585
R10182 gnd.n5993 gnd.n5261 585
R10183 gnd.n5979 gnd.n5285 585
R10184 gnd.n5285 gnd.n5274 585
R10185 gnd.n5981 gnd.n5980 585
R10186 gnd.n5982 gnd.n5981 585
R10187 gnd.n5286 gnd.n5284 585
R10188 gnd.n5284 gnd.n5281 585
R10189 gnd.n5974 gnd.n5973 585
R10190 gnd.n5973 gnd.n5972 585
R10191 gnd.n5289 gnd.n5288 585
R10192 gnd.n5347 gnd.n5289 585
R10193 gnd.n5934 gnd.n5360 585
R10194 gnd.n5360 gnd.n5346 585
R10195 gnd.n5936 gnd.n5935 585
R10196 gnd.n5937 gnd.n5936 585
R10197 gnd.n5361 gnd.n5359 585
R10198 gnd.n5368 gnd.n5359 585
R10199 gnd.n5929 gnd.n5928 585
R10200 gnd.n5928 gnd.n5927 585
R10201 gnd.n5364 gnd.n5363 585
R10202 gnd.n5908 gnd.n5364 585
R10203 gnd.n5894 gnd.n5387 585
R10204 gnd.n5387 gnd.n5377 585
R10205 gnd.n5896 gnd.n5895 585
R10206 gnd.n5897 gnd.n5896 585
R10207 gnd.n5388 gnd.n5386 585
R10208 gnd.n5885 gnd.n5386 585
R10209 gnd.n5889 gnd.n5888 585
R10210 gnd.n5888 gnd.n5887 585
R10211 gnd.n5391 gnd.n5390 585
R10212 gnd.n5851 gnd.n5391 585
R10213 gnd.n5835 gnd.n5834 585
R10214 gnd.n5834 gnd.n5401 585
R10215 gnd.n5836 gnd.n5420 585
R10216 gnd.n5420 gnd.n5400 585
R10217 gnd.n5838 gnd.n5837 585
R10218 gnd.n5839 gnd.n5838 585
R10219 gnd.n5421 gnd.n5419 585
R10220 gnd.n5419 gnd.n5416 585
R10221 gnd.n5828 gnd.n5827 585
R10222 gnd.n5827 gnd.n5826 585
R10223 gnd.n5424 gnd.n5423 585
R10224 gnd.n5433 gnd.n5424 585
R10225 gnd.n5799 gnd.n5446 585
R10226 gnd.n5446 gnd.n5432 585
R10227 gnd.n5801 gnd.n5800 585
R10228 gnd.n5802 gnd.n5801 585
R10229 gnd.n5447 gnd.n5445 585
R10230 gnd.n5454 gnd.n5445 585
R10231 gnd.n5794 gnd.n5793 585
R10232 gnd.n5793 gnd.n5792 585
R10233 gnd.n5450 gnd.n5449 585
R10234 gnd.n5773 gnd.n5450 585
R10235 gnd.n5769 gnd.n5768 585
R10236 gnd.n5770 gnd.n5769 585
R10237 gnd.n5468 gnd.n5467 585
R10238 gnd.n5475 gnd.n5467 585
R10239 gnd.n5764 gnd.n5763 585
R10240 gnd.n5763 gnd.n5762 585
R10241 gnd.n5471 gnd.n5470 585
R10242 gnd.n5752 gnd.n5471 585
R10243 gnd.n5739 gnd.n5738 585
R10244 gnd.n5737 gnd.n5690 585
R10245 gnd.n5736 gnd.n5689 585
R10246 gnd.n5741 gnd.n5689 585
R10247 gnd.n5735 gnd.n5734 585
R10248 gnd.n5733 gnd.n5732 585
R10249 gnd.n5731 gnd.n5730 585
R10250 gnd.n5729 gnd.n5728 585
R10251 gnd.n5727 gnd.n5726 585
R10252 gnd.n5725 gnd.n5724 585
R10253 gnd.n5723 gnd.n5722 585
R10254 gnd.n5721 gnd.n5720 585
R10255 gnd.n5719 gnd.n5718 585
R10256 gnd.n5717 gnd.n5716 585
R10257 gnd.n5715 gnd.n5714 585
R10258 gnd.n5713 gnd.n5712 585
R10259 gnd.n5711 gnd.n5710 585
R10260 gnd.n5706 gnd.n5482 585
R10261 gnd.n6391 gnd.n5160 585
R10262 gnd.n6463 gnd.n6462 585
R10263 gnd.n6465 gnd.n6464 585
R10264 gnd.n6467 gnd.n6466 585
R10265 gnd.n6469 gnd.n6468 585
R10266 gnd.n6471 gnd.n6470 585
R10267 gnd.n6473 gnd.n6472 585
R10268 gnd.n6475 gnd.n6474 585
R10269 gnd.n6477 gnd.n6476 585
R10270 gnd.n6479 gnd.n6478 585
R10271 gnd.n6481 gnd.n6480 585
R10272 gnd.n6483 gnd.n6482 585
R10273 gnd.n6485 gnd.n6484 585
R10274 gnd.n6486 gnd.n5146 585
R10275 gnd.n6488 gnd.n6487 585
R10276 gnd.n965 gnd.n964 585
R10277 gnd.n6492 gnd.n6491 585
R10278 gnd.n6491 gnd.n6490 585
R10279 gnd.n6393 gnd.n6392 585
R10280 gnd.n6392 gnd.n966 585
R10281 gnd.n6394 gnd.n955 585
R10282 gnd.n6498 gnd.n955 585
R10283 gnd.n6396 gnd.n6395 585
R10284 gnd.n6397 gnd.n6396 585
R10285 gnd.n6387 gnd.n5197 585
R10286 gnd.n5197 gnd.n945 585
R10287 gnd.n6385 gnd.n943 585
R10288 gnd.n6506 gnd.n943 585
R10289 gnd.n5200 gnd.n5199 585
R10290 gnd.n5199 gnd.n5198 585
R10291 gnd.n6123 gnd.n930 585
R10292 gnd.n6512 gnd.n930 585
R10293 gnd.n6122 gnd.n6121 585
R10294 gnd.n6121 gnd.n6120 585
R10295 gnd.n5204 gnd.n5202 585
R10296 gnd.n5204 gnd.n920 585
R10297 gnd.n6099 gnd.n918 585
R10298 gnd.n6520 gnd.n918 585
R10299 gnd.n6101 gnd.n6100 585
R10300 gnd.n6102 gnd.n6101 585
R10301 gnd.n5209 gnd.n908 585
R10302 gnd.n6526 gnd.n908 585
R10303 gnd.n6088 gnd.n6087 585
R10304 gnd.n6089 gnd.n6088 585
R10305 gnd.n5217 gnd.n5216 585
R10306 gnd.n5216 gnd.n5214 585
R10307 gnd.n6061 gnd.n5223 585
R10308 gnd.n6077 gnd.n5223 585
R10309 gnd.n6063 gnd.n6062 585
R10310 gnd.n6064 gnd.n6063 585
R10311 gnd.n5233 gnd.n5231 585
R10312 gnd.n6066 gnd.n5231 585
R10313 gnd.n6027 gnd.n5251 585
R10314 gnd.n6027 gnd.n5237 585
R10315 gnd.n6029 gnd.n6028 585
R10316 gnd.n6028 gnd.n5245 585
R10317 gnd.n6026 gnd.n5250 585
R10318 gnd.n6026 gnd.n5243 585
R10319 gnd.n6025 gnd.n5253 585
R10320 gnd.n6025 gnd.n6024 585
R10321 gnd.n6002 gnd.n5252 585
R10322 gnd.n5265 gnd.n5252 585
R10323 gnd.n6001 gnd.n5263 585
R10324 gnd.n6011 gnd.n5263 585
R10325 gnd.n5992 gnd.n5270 585
R10326 gnd.n5993 gnd.n5992 585
R10327 gnd.n5991 gnd.n5990 585
R10328 gnd.n5991 gnd.n5274 585
R10329 gnd.n5989 gnd.n5276 585
R10330 gnd.n5982 gnd.n5276 585
R10331 gnd.n5291 gnd.n5277 585
R10332 gnd.n5291 gnd.n5281 585
R10333 gnd.n5942 gnd.n5292 585
R10334 gnd.n5972 gnd.n5292 585
R10335 gnd.n5941 gnd.n5940 585
R10336 gnd.n5940 gnd.n5347 585
R10337 gnd.n5939 gnd.n5354 585
R10338 gnd.n5939 gnd.n5346 585
R10339 gnd.n5938 gnd.n5356 585
R10340 gnd.n5938 gnd.n5937 585
R10341 gnd.n5917 gnd.n5355 585
R10342 gnd.n5368 gnd.n5355 585
R10343 gnd.n5916 gnd.n5366 585
R10344 gnd.n5927 gnd.n5366 585
R10345 gnd.n5907 gnd.n5373 585
R10346 gnd.n5908 gnd.n5907 585
R10347 gnd.n5906 gnd.n5905 585
R10348 gnd.n5906 gnd.n5377 585
R10349 gnd.n5904 gnd.n5379 585
R10350 gnd.n5897 gnd.n5379 585
R10351 gnd.n5884 gnd.n5380 585
R10352 gnd.n5885 gnd.n5884 585
R10353 gnd.n5854 gnd.n5393 585
R10354 gnd.n5887 gnd.n5393 585
R10355 gnd.n5853 gnd.n5852 585
R10356 gnd.n5852 gnd.n5851 585
R10357 gnd.n5849 gnd.n5410 585
R10358 gnd.n5849 gnd.n5401 585
R10359 gnd.n5848 gnd.n5847 585
R10360 gnd.n5848 gnd.n5400 585
R10361 gnd.n5412 gnd.n5411 585
R10362 gnd.n5839 gnd.n5411 585
R10363 gnd.n5808 gnd.n5807 585
R10364 gnd.n5807 gnd.n5416 585
R10365 gnd.n5809 gnd.n5426 585
R10366 gnd.n5826 gnd.n5426 585
R10367 gnd.n5806 gnd.n5805 585
R10368 gnd.n5805 gnd.n5433 585
R10369 gnd.n5804 gnd.n5440 585
R10370 gnd.n5804 gnd.n5432 585
R10371 gnd.n5803 gnd.n5442 585
R10372 gnd.n5803 gnd.n5802 585
R10373 gnd.n5782 gnd.n5441 585
R10374 gnd.n5454 gnd.n5441 585
R10375 gnd.n5781 gnd.n5452 585
R10376 gnd.n5792 gnd.n5452 585
R10377 gnd.n5772 gnd.n5459 585
R10378 gnd.n5773 gnd.n5772 585
R10379 gnd.n5771 gnd.n5465 585
R10380 gnd.n5771 gnd.n5770 585
R10381 gnd.n5756 gnd.n5464 585
R10382 gnd.n5475 gnd.n5464 585
R10383 gnd.n5755 gnd.n5473 585
R10384 gnd.n5762 gnd.n5473 585
R10385 gnd.n5754 gnd.n5753 585
R10386 gnd.n5753 gnd.n5752 585
R10387 gnd.n4902 gnd.n4901 585
R10388 gnd.n4901 gnd.n4900 585
R10389 gnd.n4903 gnd.n1314 585
R10390 gnd.n3450 gnd.n1314 585
R10391 gnd.n4905 gnd.n4904 585
R10392 gnd.n4906 gnd.n4905 585
R10393 gnd.n1299 gnd.n1298 585
R10394 gnd.n3285 gnd.n1299 585
R10395 gnd.n4914 gnd.n4913 585
R10396 gnd.n4913 gnd.n4912 585
R10397 gnd.n4915 gnd.n1293 585
R10398 gnd.n3276 gnd.n1293 585
R10399 gnd.n4917 gnd.n4916 585
R10400 gnd.n4918 gnd.n4917 585
R10401 gnd.n1277 gnd.n1276 585
R10402 gnd.n3272 gnd.n1277 585
R10403 gnd.n4926 gnd.n4925 585
R10404 gnd.n4925 gnd.n4924 585
R10405 gnd.n4927 gnd.n1271 585
R10406 gnd.n3299 gnd.n1271 585
R10407 gnd.n4929 gnd.n4928 585
R10408 gnd.n4930 gnd.n4929 585
R10409 gnd.n1257 gnd.n1256 585
R10410 gnd.n3264 gnd.n1257 585
R10411 gnd.n4938 gnd.n4937 585
R10412 gnd.n4937 gnd.n4936 585
R10413 gnd.n4939 gnd.n1251 585
R10414 gnd.n3256 gnd.n1251 585
R10415 gnd.n4941 gnd.n4940 585
R10416 gnd.n4942 gnd.n4941 585
R10417 gnd.n1235 gnd.n1234 585
R10418 gnd.n3247 gnd.n1235 585
R10419 gnd.n4950 gnd.n4949 585
R10420 gnd.n4949 gnd.n4948 585
R10421 gnd.n4951 gnd.n1229 585
R10422 gnd.n3239 gnd.n1229 585
R10423 gnd.n4953 gnd.n4952 585
R10424 gnd.n4954 gnd.n4953 585
R10425 gnd.n1215 gnd.n1214 585
R10426 gnd.n3231 gnd.n1215 585
R10427 gnd.n4962 gnd.n4961 585
R10428 gnd.n4961 gnd.n4960 585
R10429 gnd.n4963 gnd.n1210 585
R10430 gnd.n3223 gnd.n1210 585
R10431 gnd.n4965 gnd.n4964 585
R10432 gnd.n4966 gnd.n4965 585
R10433 gnd.n1211 gnd.n1194 585
R10434 gnd.n3215 gnd.n1194 585
R10435 gnd.n4974 gnd.n4973 585
R10436 gnd.n4973 gnd.n4972 585
R10437 gnd.n4975 gnd.n1191 585
R10438 gnd.n3207 gnd.n1191 585
R10439 gnd.n4978 gnd.n4977 585
R10440 gnd.n4979 gnd.n4978 585
R10441 gnd.n1192 gnd.n1177 585
R10442 gnd.n3198 gnd.n1177 585
R10443 gnd.n4987 gnd.n4986 585
R10444 gnd.n4986 gnd.n4985 585
R10445 gnd.n4988 gnd.n1173 585
R10446 gnd.n3189 gnd.n1173 585
R10447 gnd.n4990 gnd.n4989 585
R10448 gnd.n4991 gnd.n4990 585
R10449 gnd.n1157 gnd.n1156 585
R10450 gnd.n3181 gnd.n1157 585
R10451 gnd.n4999 gnd.n4998 585
R10452 gnd.n4998 gnd.n4997 585
R10453 gnd.n5000 gnd.n1151 585
R10454 gnd.n3173 gnd.n1151 585
R10455 gnd.n5002 gnd.n5001 585
R10456 gnd.n5003 gnd.n5002 585
R10457 gnd.n1137 gnd.n1136 585
R10458 gnd.n3165 gnd.n1137 585
R10459 gnd.n5011 gnd.n5010 585
R10460 gnd.n5010 gnd.n5009 585
R10461 gnd.n5012 gnd.n1131 585
R10462 gnd.n3157 gnd.n1131 585
R10463 gnd.n5014 gnd.n5013 585
R10464 gnd.n5015 gnd.n5014 585
R10465 gnd.n1115 gnd.n1114 585
R10466 gnd.n3149 gnd.n1115 585
R10467 gnd.n5023 gnd.n5022 585
R10468 gnd.n5022 gnd.n5021 585
R10469 gnd.n5024 gnd.n1109 585
R10470 gnd.n3141 gnd.n1109 585
R10471 gnd.n5026 gnd.n5025 585
R10472 gnd.n5027 gnd.n5026 585
R10473 gnd.n1095 gnd.n1094 585
R10474 gnd.n1105 gnd.n1095 585
R10475 gnd.n5035 gnd.n5034 585
R10476 gnd.n5034 gnd.n5033 585
R10477 gnd.n5036 gnd.n1089 585
R10478 gnd.n1089 gnd.n1088 585
R10479 gnd.n5038 gnd.n5037 585
R10480 gnd.n5039 gnd.n5038 585
R10481 gnd.n1074 gnd.n1073 585
R10482 gnd.n1077 gnd.n1074 585
R10483 gnd.n5047 gnd.n5046 585
R10484 gnd.n5046 gnd.n5045 585
R10485 gnd.n5048 gnd.n1068 585
R10486 gnd.n1068 gnd.n1065 585
R10487 gnd.n5050 gnd.n5049 585
R10488 gnd.n5051 gnd.n5050 585
R10489 gnd.n1069 gnd.n1067 585
R10490 gnd.n1067 gnd.n1063 585
R10491 gnd.n3099 gnd.n3098 585
R10492 gnd.n3100 gnd.n3099 585
R10493 gnd.n3094 gnd.n1012 585
R10494 gnd.n1012 gnd.n1009 585
R10495 gnd.n5136 gnd.n5135 585
R10496 gnd.n5134 gnd.n1011 585
R10497 gnd.n5133 gnd.n1010 585
R10498 gnd.n5138 gnd.n1010 585
R10499 gnd.n5132 gnd.n5131 585
R10500 gnd.n5130 gnd.n5129 585
R10501 gnd.n5128 gnd.n5127 585
R10502 gnd.n5126 gnd.n5125 585
R10503 gnd.n5124 gnd.n5123 585
R10504 gnd.n5122 gnd.n5121 585
R10505 gnd.n5120 gnd.n5119 585
R10506 gnd.n5118 gnd.n5117 585
R10507 gnd.n5116 gnd.n5115 585
R10508 gnd.n5114 gnd.n5113 585
R10509 gnd.n5112 gnd.n5111 585
R10510 gnd.n5110 gnd.n5109 585
R10511 gnd.n5108 gnd.n5107 585
R10512 gnd.n5106 gnd.n5105 585
R10513 gnd.n5104 gnd.n5103 585
R10514 gnd.n5101 gnd.n5100 585
R10515 gnd.n5099 gnd.n5098 585
R10516 gnd.n5097 gnd.n5096 585
R10517 gnd.n5095 gnd.n5094 585
R10518 gnd.n5093 gnd.n5092 585
R10519 gnd.n5091 gnd.n5090 585
R10520 gnd.n5089 gnd.n5088 585
R10521 gnd.n5087 gnd.n5086 585
R10522 gnd.n5085 gnd.n5084 585
R10523 gnd.n5083 gnd.n5082 585
R10524 gnd.n5081 gnd.n5080 585
R10525 gnd.n5079 gnd.n5078 585
R10526 gnd.n5077 gnd.n5076 585
R10527 gnd.n5075 gnd.n5074 585
R10528 gnd.n5073 gnd.n5072 585
R10529 gnd.n5071 gnd.n5070 585
R10530 gnd.n5069 gnd.n5068 585
R10531 gnd.n5067 gnd.n5066 585
R10532 gnd.n5065 gnd.n1051 585
R10533 gnd.n1055 gnd.n1052 585
R10534 gnd.n5061 gnd.n5060 585
R10535 gnd.n3457 gnd.n3456 585
R10536 gnd.n3459 gnd.n2636 585
R10537 gnd.n3461 gnd.n3460 585
R10538 gnd.n3462 gnd.n2629 585
R10539 gnd.n3464 gnd.n3463 585
R10540 gnd.n3466 gnd.n2627 585
R10541 gnd.n3468 gnd.n3467 585
R10542 gnd.n3469 gnd.n2622 585
R10543 gnd.n3471 gnd.n3470 585
R10544 gnd.n3473 gnd.n2620 585
R10545 gnd.n3475 gnd.n3474 585
R10546 gnd.n3476 gnd.n2615 585
R10547 gnd.n3478 gnd.n3477 585
R10548 gnd.n3480 gnd.n2613 585
R10549 gnd.n3482 gnd.n3481 585
R10550 gnd.n3483 gnd.n2608 585
R10551 gnd.n3485 gnd.n3484 585
R10552 gnd.n3487 gnd.n2607 585
R10553 gnd.n3488 gnd.n2550 585
R10554 gnd.n3491 gnd.n3490 585
R10555 gnd.n2551 gnd.n2543 585
R10556 gnd.n2579 gnd.n2544 585
R10557 gnd.n2581 gnd.n2580 585
R10558 gnd.n2583 gnd.n2582 585
R10559 gnd.n2585 gnd.n2584 585
R10560 gnd.n2587 gnd.n2586 585
R10561 gnd.n2589 gnd.n2588 585
R10562 gnd.n2591 gnd.n2590 585
R10563 gnd.n2593 gnd.n2592 585
R10564 gnd.n2595 gnd.n2594 585
R10565 gnd.n2597 gnd.n2596 585
R10566 gnd.n2599 gnd.n2598 585
R10567 gnd.n2601 gnd.n2600 585
R10568 gnd.n2602 gnd.n2561 585
R10569 gnd.n2604 gnd.n2603 585
R10570 gnd.n2562 gnd.n2560 585
R10571 gnd.n2563 gnd.n1319 585
R10572 gnd.n2606 gnd.n1319 585
R10573 gnd.n3453 gnd.n1321 585
R10574 gnd.n4900 gnd.n1321 585
R10575 gnd.n3452 gnd.n3451 585
R10576 gnd.n3451 gnd.n3450 585
R10577 gnd.n2640 gnd.n1312 585
R10578 gnd.n4906 gnd.n1312 585
R10579 gnd.n3284 gnd.n3283 585
R10580 gnd.n3285 gnd.n3284 585
R10581 gnd.n2866 gnd.n1301 585
R10582 gnd.n4912 gnd.n1301 585
R10583 gnd.n3278 gnd.n3277 585
R10584 gnd.n3277 gnd.n3276 585
R10585 gnd.n3275 gnd.n1290 585
R10586 gnd.n4918 gnd.n1290 585
R10587 gnd.n3274 gnd.n3273 585
R10588 gnd.n3273 gnd.n3272 585
R10589 gnd.n2868 gnd.n1279 585
R10590 gnd.n4924 gnd.n1279 585
R10591 gnd.n3268 gnd.n2858 585
R10592 gnd.n3299 gnd.n2858 585
R10593 gnd.n3267 gnd.n1269 585
R10594 gnd.n4930 gnd.n1269 585
R10595 gnd.n3266 gnd.n3265 585
R10596 gnd.n3265 gnd.n3264 585
R10597 gnd.n2870 gnd.n1259 585
R10598 gnd.n4936 gnd.n1259 585
R10599 gnd.n3255 gnd.n3254 585
R10600 gnd.n3256 gnd.n3255 585
R10601 gnd.n2876 gnd.n1248 585
R10602 gnd.n4942 gnd.n1248 585
R10603 gnd.n3249 gnd.n3248 585
R10604 gnd.n3248 gnd.n3247 585
R10605 gnd.n2878 gnd.n1237 585
R10606 gnd.n4948 gnd.n1237 585
R10607 gnd.n3238 gnd.n3237 585
R10608 gnd.n3239 gnd.n3238 585
R10609 gnd.n2883 gnd.n1227 585
R10610 gnd.n4954 gnd.n1227 585
R10611 gnd.n3233 gnd.n3232 585
R10612 gnd.n3232 gnd.n3231 585
R10613 gnd.n2885 gnd.n1217 585
R10614 gnd.n4960 gnd.n1217 585
R10615 gnd.n3222 gnd.n3221 585
R10616 gnd.n3223 gnd.n3222 585
R10617 gnd.n2890 gnd.n1207 585
R10618 gnd.n4966 gnd.n1207 585
R10619 gnd.n3217 gnd.n3216 585
R10620 gnd.n3216 gnd.n3215 585
R10621 gnd.n2892 gnd.n1196 585
R10622 gnd.n4972 gnd.n1196 585
R10623 gnd.n3206 gnd.n3205 585
R10624 gnd.n3207 gnd.n3206 585
R10625 gnd.n2897 gnd.n1189 585
R10626 gnd.n4979 gnd.n1189 585
R10627 gnd.n3200 gnd.n3199 585
R10628 gnd.n3199 gnd.n3198 585
R10629 gnd.n2900 gnd.n1179 585
R10630 gnd.n4985 gnd.n1179 585
R10631 gnd.n3188 gnd.n3187 585
R10632 gnd.n3189 gnd.n3188 585
R10633 gnd.n2905 gnd.n1170 585
R10634 gnd.n4991 gnd.n1170 585
R10635 gnd.n3183 gnd.n3182 585
R10636 gnd.n3182 gnd.n3181 585
R10637 gnd.n2907 gnd.n1159 585
R10638 gnd.n4997 gnd.n1159 585
R10639 gnd.n3172 gnd.n3171 585
R10640 gnd.n3173 gnd.n3172 585
R10641 gnd.n2912 gnd.n1149 585
R10642 gnd.n5003 gnd.n1149 585
R10643 gnd.n3167 gnd.n3166 585
R10644 gnd.n3166 gnd.n3165 585
R10645 gnd.n2914 gnd.n1139 585
R10646 gnd.n5009 gnd.n1139 585
R10647 gnd.n3156 gnd.n3155 585
R10648 gnd.n3157 gnd.n3156 585
R10649 gnd.n3009 gnd.n1128 585
R10650 gnd.n5015 gnd.n1128 585
R10651 gnd.n3151 gnd.n3150 585
R10652 gnd.n3150 gnd.n3149 585
R10653 gnd.n3011 gnd.n1117 585
R10654 gnd.n5021 gnd.n1117 585
R10655 gnd.n3140 gnd.n3139 585
R10656 gnd.n3141 gnd.n3140 585
R10657 gnd.n3121 gnd.n1106 585
R10658 gnd.n5027 gnd.n1106 585
R10659 gnd.n3135 gnd.n3134 585
R10660 gnd.n3134 gnd.n1105 585
R10661 gnd.n3133 gnd.n1096 585
R10662 gnd.n5033 gnd.n1096 585
R10663 gnd.n3132 gnd.n3131 585
R10664 gnd.n3131 gnd.n1088 585
R10665 gnd.n3123 gnd.n1086 585
R10666 gnd.n5039 gnd.n1086 585
R10667 gnd.n3127 gnd.n3126 585
R10668 gnd.n3126 gnd.n1077 585
R10669 gnd.n3125 gnd.n1075 585
R10670 gnd.n5045 gnd.n1075 585
R10671 gnd.n1062 gnd.n1060 585
R10672 gnd.n1065 gnd.n1062 585
R10673 gnd.n5053 gnd.n5052 585
R10674 gnd.n5052 gnd.n5051 585
R10675 gnd.n1061 gnd.n1058 585
R10676 gnd.n1063 gnd.n1061 585
R10677 gnd.n5057 gnd.n1057 585
R10678 gnd.n3100 gnd.n1057 585
R10679 gnd.n5059 gnd.n5058 585
R10680 gnd.n5059 gnd.n1009 585
R10681 gnd.n7742 gnd.n7741 585
R10682 gnd.n7743 gnd.n7742 585
R10683 gnd.n110 gnd.n108 585
R10684 gnd.n108 gnd.n104 585
R10685 gnd.n7662 gnd.n7661 585
R10686 gnd.n7663 gnd.n7662 585
R10687 gnd.n189 gnd.n188 585
R10688 gnd.n188 gnd.n186 585
R10689 gnd.n7657 gnd.n7656 585
R10690 gnd.n7656 gnd.n7655 585
R10691 gnd.n192 gnd.n191 585
R10692 gnd.n193 gnd.n192 585
R10693 gnd.n7571 gnd.n7570 585
R10694 gnd.n7572 gnd.n7571 585
R10695 gnd.n204 gnd.n203 585
R10696 gnd.n211 gnd.n203 585
R10697 gnd.n7566 gnd.n7565 585
R10698 gnd.n7565 gnd.n7564 585
R10699 gnd.n207 gnd.n206 585
R10700 gnd.n208 gnd.n207 585
R10701 gnd.n7555 gnd.n7554 585
R10702 gnd.n7556 gnd.n7555 585
R10703 gnd.n221 gnd.n220 585
R10704 gnd.n220 gnd.n218 585
R10705 gnd.n7550 gnd.n7549 585
R10706 gnd.n7549 gnd.n7548 585
R10707 gnd.n224 gnd.n223 585
R10708 gnd.n7450 gnd.n224 585
R10709 gnd.n7539 gnd.n7538 585
R10710 gnd.n7540 gnd.n7539 585
R10711 gnd.n235 gnd.n234 585
R10712 gnd.n7457 gnd.n234 585
R10713 gnd.n7534 gnd.n7533 585
R10714 gnd.n7533 gnd.n7532 585
R10715 gnd.n238 gnd.n237 585
R10716 gnd.n7417 gnd.n238 585
R10717 gnd.n7523 gnd.n7522 585
R10718 gnd.n7524 gnd.n7523 585
R10719 gnd.n251 gnd.n250 585
R10720 gnd.n7413 gnd.n250 585
R10721 gnd.n7518 gnd.n7517 585
R10722 gnd.n7517 gnd.n7516 585
R10723 gnd.n254 gnd.n253 585
R10724 gnd.n7406 gnd.n254 585
R10725 gnd.n7507 gnd.n7506 585
R10726 gnd.n7508 gnd.n7507 585
R10727 gnd.n266 gnd.n265 585
R10728 gnd.n7474 gnd.n265 585
R10729 gnd.n7484 gnd.n7483 585
R10730 gnd.n7485 gnd.n7484 585
R10731 gnd.n7482 gnd.n7481 585
R10732 gnd.n7481 gnd.n7480 585
R10733 gnd.n1546 gnd.n297 585
R10734 gnd.n4648 gnd.n297 585
R10735 gnd.n4661 gnd.n1547 585
R10736 gnd.n4661 gnd.n4660 585
R10737 gnd.n4663 gnd.n4662 585
R10738 gnd.n4664 gnd.n4663 585
R10739 gnd.n1545 gnd.n272 585
R10740 gnd.n1545 gnd.n1541 585
R10741 gnd.n276 gnd.n273 585
R10742 gnd.n4637 gnd.n276 585
R10743 gnd.n7503 gnd.n7502 585
R10744 gnd.n7502 gnd.n7501 585
R10745 gnd.n275 gnd.n274 585
R10746 gnd.n4625 gnd.n275 585
R10747 gnd.n4686 gnd.n4685 585
R10748 gnd.n4687 gnd.n4686 585
R10749 gnd.n1522 gnd.n1521 585
R10750 gnd.n1528 gnd.n1521 585
R10751 gnd.n4681 gnd.n4680 585
R10752 gnd.n4680 gnd.n4679 585
R10753 gnd.n1525 gnd.n1524 585
R10754 gnd.n4612 gnd.n1525 585
R10755 gnd.n4596 gnd.n1573 585
R10756 gnd.n1573 gnd.n1572 585
R10757 gnd.n4598 gnd.n4597 585
R10758 gnd.n4599 gnd.n4598 585
R10759 gnd.n1574 gnd.n1570 585
R10760 gnd.n1581 gnd.n1570 585
R10761 gnd.n4591 gnd.n4590 585
R10762 gnd.n4590 gnd.n4589 585
R10763 gnd.n1577 gnd.n1576 585
R10764 gnd.n4570 gnd.n1577 585
R10765 gnd.n4557 gnd.n1600 585
R10766 gnd.n1600 gnd.n1589 585
R10767 gnd.n4559 gnd.n4558 585
R10768 gnd.n4560 gnd.n4559 585
R10769 gnd.n1601 gnd.n1599 585
R10770 gnd.n1608 gnd.n1599 585
R10771 gnd.n4552 gnd.n4551 585
R10772 gnd.n4551 gnd.n4550 585
R10773 gnd.n1604 gnd.n1603 585
R10774 gnd.n4537 gnd.n1604 585
R10775 gnd.n4525 gnd.n4521 585
R10776 gnd.n4521 gnd.n1616 585
R10777 gnd.n4527 gnd.n4526 585
R10778 gnd.n4528 gnd.n4527 585
R10779 gnd.n1489 gnd.n1488 585
R10780 gnd.n1635 gnd.n1489 585
R10781 gnd.n4720 gnd.n4719 585
R10782 gnd.n4719 gnd.n4718 585
R10783 gnd.n4721 gnd.n1483 585
R10784 gnd.n4487 gnd.n1483 585
R10785 gnd.n4723 gnd.n4722 585
R10786 gnd.n4724 gnd.n4723 585
R10787 gnd.n1484 gnd.n1482 585
R10788 gnd.n1482 gnd.n1477 585
R10789 gnd.n1909 gnd.n1908 585
R10790 gnd.n1912 gnd.n1911 585
R10791 gnd.n1905 gnd.n1904 585
R10792 gnd.n1904 gnd.n1468 585
R10793 gnd.n1917 gnd.n1916 585
R10794 gnd.n1919 gnd.n1903 585
R10795 gnd.n1922 gnd.n1921 585
R10796 gnd.n1901 gnd.n1900 585
R10797 gnd.n1927 gnd.n1926 585
R10798 gnd.n1929 gnd.n1899 585
R10799 gnd.n1932 gnd.n1931 585
R10800 gnd.n1897 gnd.n1896 585
R10801 gnd.n1938 gnd.n1937 585
R10802 gnd.n1940 gnd.n1895 585
R10803 gnd.n1941 gnd.n1892 585
R10804 gnd.n1944 gnd.n1943 585
R10805 gnd.n1894 gnd.n1889 585
R10806 gnd.n2029 gnd.n2028 585
R10807 gnd.n2026 gnd.n1951 585
R10808 gnd.n2024 gnd.n2023 585
R10809 gnd.n2022 gnd.n1952 585
R10810 gnd.n2021 gnd.n2020 585
R10811 gnd.n2018 gnd.n1957 585
R10812 gnd.n2016 gnd.n2015 585
R10813 gnd.n2014 gnd.n1958 585
R10814 gnd.n2013 gnd.n2012 585
R10815 gnd.n2010 gnd.n1963 585
R10816 gnd.n2008 gnd.n2007 585
R10817 gnd.n2006 gnd.n1964 585
R10818 gnd.n2005 gnd.n2004 585
R10819 gnd.n2002 gnd.n1969 585
R10820 gnd.n2000 gnd.n1999 585
R10821 gnd.n1998 gnd.n1970 585
R10822 gnd.n1997 gnd.n1996 585
R10823 gnd.n1994 gnd.n1975 585
R10824 gnd.n1992 gnd.n1991 585
R10825 gnd.n1979 gnd.n1976 585
R10826 gnd.n1987 gnd.n1986 585
R10827 gnd.n179 gnd.n178 585
R10828 gnd.n7671 gnd.n174 585
R10829 gnd.n7673 gnd.n7672 585
R10830 gnd.n7675 gnd.n172 585
R10831 gnd.n7677 gnd.n7676 585
R10832 gnd.n7678 gnd.n167 585
R10833 gnd.n7680 gnd.n7679 585
R10834 gnd.n7682 gnd.n165 585
R10835 gnd.n7684 gnd.n7683 585
R10836 gnd.n7685 gnd.n160 585
R10837 gnd.n7687 gnd.n7686 585
R10838 gnd.n7689 gnd.n158 585
R10839 gnd.n7691 gnd.n7690 585
R10840 gnd.n7692 gnd.n153 585
R10841 gnd.n7694 gnd.n7693 585
R10842 gnd.n7696 gnd.n151 585
R10843 gnd.n7698 gnd.n7697 585
R10844 gnd.n7699 gnd.n146 585
R10845 gnd.n7701 gnd.n7700 585
R10846 gnd.n7703 gnd.n144 585
R10847 gnd.n7705 gnd.n7704 585
R10848 gnd.n7709 gnd.n139 585
R10849 gnd.n7711 gnd.n7710 585
R10850 gnd.n7713 gnd.n137 585
R10851 gnd.n7715 gnd.n7714 585
R10852 gnd.n7716 gnd.n132 585
R10853 gnd.n7718 gnd.n7717 585
R10854 gnd.n7720 gnd.n130 585
R10855 gnd.n7722 gnd.n7721 585
R10856 gnd.n7723 gnd.n125 585
R10857 gnd.n7725 gnd.n7724 585
R10858 gnd.n7727 gnd.n123 585
R10859 gnd.n7729 gnd.n7728 585
R10860 gnd.n7730 gnd.n118 585
R10861 gnd.n7732 gnd.n7731 585
R10862 gnd.n7734 gnd.n115 585
R10863 gnd.n7736 gnd.n7735 585
R10864 gnd.n7737 gnd.n113 585
R10865 gnd.n7738 gnd.n109 585
R10866 gnd.n117 gnd.n109 585
R10867 gnd.n7667 gnd.n105 585
R10868 gnd.n7743 gnd.n105 585
R10869 gnd.n7666 gnd.n7665 585
R10870 gnd.n7665 gnd.n104 585
R10871 gnd.n7664 gnd.n183 585
R10872 gnd.n7664 gnd.n7663 585
R10873 gnd.n7436 gnd.n184 585
R10874 gnd.n186 gnd.n184 585
R10875 gnd.n7437 gnd.n194 585
R10876 gnd.n7655 gnd.n194 585
R10877 gnd.n7439 gnd.n7438 585
R10878 gnd.n7438 gnd.n193 585
R10879 gnd.n7440 gnd.n202 585
R10880 gnd.n7572 gnd.n202 585
R10881 gnd.n7442 gnd.n7441 585
R10882 gnd.n7441 gnd.n211 585
R10883 gnd.n7443 gnd.n209 585
R10884 gnd.n7564 gnd.n209 585
R10885 gnd.n7445 gnd.n7444 585
R10886 gnd.n7444 gnd.n208 585
R10887 gnd.n7446 gnd.n219 585
R10888 gnd.n7556 gnd.n219 585
R10889 gnd.n7448 gnd.n7447 585
R10890 gnd.n7447 gnd.n218 585
R10891 gnd.n7449 gnd.n226 585
R10892 gnd.n7548 gnd.n226 585
R10893 gnd.n7452 gnd.n7451 585
R10894 gnd.n7451 gnd.n7450 585
R10895 gnd.n7453 gnd.n232 585
R10896 gnd.n7540 gnd.n232 585
R10897 gnd.n7455 gnd.n7454 585
R10898 gnd.n7457 gnd.n7455 585
R10899 gnd.n7402 gnd.n240 585
R10900 gnd.n7532 gnd.n240 585
R10901 gnd.n7419 gnd.n7418 585
R10902 gnd.n7418 gnd.n7417 585
R10903 gnd.n7416 gnd.n248 585
R10904 gnd.n7524 gnd.n248 585
R10905 gnd.n7415 gnd.n7414 585
R10906 gnd.n7414 gnd.n7413 585
R10907 gnd.n7404 gnd.n256 585
R10908 gnd.n7516 gnd.n256 585
R10909 gnd.n7408 gnd.n7407 585
R10910 gnd.n7407 gnd.n7406 585
R10911 gnd.n304 gnd.n263 585
R10912 gnd.n7508 gnd.n263 585
R10913 gnd.n7476 gnd.n7475 585
R10914 gnd.n7475 gnd.n7474 585
R10915 gnd.n7477 gnd.n295 585
R10916 gnd.n7485 gnd.n295 585
R10917 gnd.n7479 gnd.n7478 585
R10918 gnd.n7480 gnd.n7479 585
R10919 gnd.n299 gnd.n298 585
R10920 gnd.n4648 gnd.n298 585
R10921 gnd.n4645 gnd.n4644 585
R10922 gnd.n4660 gnd.n4645 585
R10923 gnd.n1548 gnd.n1542 585
R10924 gnd.n4664 gnd.n1542 585
R10925 gnd.n4640 gnd.n4639 585
R10926 gnd.n4639 gnd.n1541 585
R10927 gnd.n4638 gnd.n1550 585
R10928 gnd.n4638 gnd.n4637 585
R10929 gnd.n4622 gnd.n278 585
R10930 gnd.n7501 gnd.n278 585
R10931 gnd.n4624 gnd.n4623 585
R10932 gnd.n4625 gnd.n4624 585
R10933 gnd.n1556 gnd.n1518 585
R10934 gnd.n4687 gnd.n1518 585
R10935 gnd.n4617 gnd.n4616 585
R10936 gnd.n4616 gnd.n1528 585
R10937 gnd.n4615 gnd.n1526 585
R10938 gnd.n4679 gnd.n1526 585
R10939 gnd.n4614 gnd.n4613 585
R10940 gnd.n4613 gnd.n4612 585
R10941 gnd.n1560 gnd.n1558 585
R10942 gnd.n1572 gnd.n1560 585
R10943 gnd.n4505 gnd.n1568 585
R10944 gnd.n4599 gnd.n1568 585
R10945 gnd.n4507 gnd.n4506 585
R10946 gnd.n4506 gnd.n1581 585
R10947 gnd.n4508 gnd.n1579 585
R10948 gnd.n4589 gnd.n1579 585
R10949 gnd.n4509 gnd.n1590 585
R10950 gnd.n4570 gnd.n1590 585
R10951 gnd.n4511 gnd.n4510 585
R10952 gnd.n4510 gnd.n1589 585
R10953 gnd.n4512 gnd.n1597 585
R10954 gnd.n4560 gnd.n1597 585
R10955 gnd.n4514 gnd.n4513 585
R10956 gnd.n4513 gnd.n1608 585
R10957 gnd.n4515 gnd.n1606 585
R10958 gnd.n4550 gnd.n1606 585
R10959 gnd.n4516 gnd.n1617 585
R10960 gnd.n4537 gnd.n1617 585
R10961 gnd.n4517 gnd.n1637 585
R10962 gnd.n1637 gnd.n1616 585
R10963 gnd.n4519 gnd.n4518 585
R10964 gnd.n4528 gnd.n4519 585
R10965 gnd.n1638 gnd.n1636 585
R10966 gnd.n1636 gnd.n1635 585
R10967 gnd.n4490 gnd.n1491 585
R10968 gnd.n4718 gnd.n1491 585
R10969 gnd.n4489 gnd.n4488 585
R10970 gnd.n4488 gnd.n4487 585
R10971 gnd.n1640 gnd.n1478 585
R10972 gnd.n4724 gnd.n1478 585
R10973 gnd.n1984 gnd.n1983 585
R10974 gnd.n1984 gnd.n1477 585
R10975 gnd.n4300 gnd.n4299 585
R10976 gnd.n4301 gnd.n4300 585
R10977 gnd.n4211 gnd.n2038 585
R10978 gnd.n4206 gnd.n2038 585
R10979 gnd.n4210 gnd.n4209 585
R10980 gnd.n4209 gnd.n4208 585
R10981 gnd.n2041 gnd.n2040 585
R10982 gnd.n4193 gnd.n2041 585
R10983 gnd.n4182 gnd.n2058 585
R10984 gnd.n2058 gnd.n2051 585
R10985 gnd.n4184 gnd.n4183 585
R10986 gnd.n4185 gnd.n4184 585
R10987 gnd.n4181 gnd.n2057 585
R10988 gnd.n2064 gnd.n2057 585
R10989 gnd.n4180 gnd.n4179 585
R10990 gnd.n4179 gnd.n4178 585
R10991 gnd.n2060 gnd.n2059 585
R10992 gnd.n4061 gnd.n2060 585
R10993 gnd.n4166 gnd.n4165 585
R10994 gnd.n4167 gnd.n4166 585
R10995 gnd.n4164 gnd.n2076 585
R10996 gnd.n2076 gnd.n2072 585
R10997 gnd.n4163 gnd.n4162 585
R10998 gnd.n4162 gnd.n4161 585
R10999 gnd.n2078 gnd.n2077 585
R11000 gnd.n4070 gnd.n2078 585
R11001 gnd.n4136 gnd.n4135 585
R11002 gnd.n4137 gnd.n4136 585
R11003 gnd.n4134 gnd.n2090 585
R11004 gnd.n2090 gnd.n2087 585
R11005 gnd.n4133 gnd.n4132 585
R11006 gnd.n4132 gnd.n4131 585
R11007 gnd.n2092 gnd.n2091 585
R11008 gnd.n4077 gnd.n2092 585
R11009 gnd.n4117 gnd.n4116 585
R11010 gnd.n4118 gnd.n4117 585
R11011 gnd.n4115 gnd.n2102 585
R11012 gnd.n4110 gnd.n2102 585
R11013 gnd.n4114 gnd.n4113 585
R11014 gnd.n4113 gnd.n4112 585
R11015 gnd.n2104 gnd.n2103 585
R11016 gnd.n2116 gnd.n2104 585
R11017 gnd.n4046 gnd.n4045 585
R11018 gnd.n4046 gnd.n2114 585
R11019 gnd.n4051 gnd.n4050 585
R11020 gnd.n4050 gnd.n4049 585
R11021 gnd.n4052 gnd.n2124 585
R11022 gnd.n4090 gnd.n2124 585
R11023 gnd.n4053 gnd.n2133 585
R11024 gnd.n2133 gnd.n2132 585
R11025 gnd.n4055 gnd.n4054 585
R11026 gnd.n4056 gnd.n4055 585
R11027 gnd.n4044 gnd.n2131 585
R11028 gnd.n4039 gnd.n2131 585
R11029 gnd.n4043 gnd.n4042 585
R11030 gnd.n4042 gnd.n4041 585
R11031 gnd.n2135 gnd.n2134 585
R11032 gnd.n4028 gnd.n2135 585
R11033 gnd.n4018 gnd.n2152 585
R11034 gnd.n2152 gnd.n2144 585
R11035 gnd.n4020 gnd.n4019 585
R11036 gnd.n4021 gnd.n4020 585
R11037 gnd.n4017 gnd.n2151 585
R11038 gnd.n2158 gnd.n2151 585
R11039 gnd.n4016 gnd.n4015 585
R11040 gnd.n4015 gnd.n4014 585
R11041 gnd.n2154 gnd.n2153 585
R11042 gnd.n3917 gnd.n2154 585
R11043 gnd.n4002 gnd.n4001 585
R11044 gnd.n4003 gnd.n4002 585
R11045 gnd.n4000 gnd.n2168 585
R11046 gnd.n2168 gnd.n2165 585
R11047 gnd.n3999 gnd.n3998 585
R11048 gnd.n3998 gnd.n3997 585
R11049 gnd.n2170 gnd.n2169 585
R11050 gnd.n3926 gnd.n2170 585
R11051 gnd.n3965 gnd.n3964 585
R11052 gnd.n3966 gnd.n3965 585
R11053 gnd.n3963 gnd.n2181 585
R11054 gnd.n2181 gnd.n2179 585
R11055 gnd.n3962 gnd.n3961 585
R11056 gnd.n3961 gnd.n3960 585
R11057 gnd.n2183 gnd.n2182 585
R11058 gnd.n3933 gnd.n2183 585
R11059 gnd.n3946 gnd.n3945 585
R11060 gnd.n3947 gnd.n3946 585
R11061 gnd.n3944 gnd.n2196 585
R11062 gnd.n3939 gnd.n2196 585
R11063 gnd.n3943 gnd.n3942 585
R11064 gnd.n3942 gnd.n3941 585
R11065 gnd.n2198 gnd.n2197 585
R11066 gnd.n3911 gnd.n2198 585
R11067 gnd.n3885 gnd.n3884 585
R11068 gnd.n3886 gnd.n3885 585
R11069 gnd.n3890 gnd.n3889 585
R11070 gnd.n3889 gnd.n3888 585
R11071 gnd.n3891 gnd.n2210 585
R11072 gnd.n3902 gnd.n2210 585
R11073 gnd.n3892 gnd.n2221 585
R11074 gnd.n2221 gnd.n2220 585
R11075 gnd.n3894 gnd.n3893 585
R11076 gnd.n3895 gnd.n3894 585
R11077 gnd.n3883 gnd.n2219 585
R11078 gnd.n3878 gnd.n2219 585
R11079 gnd.n3882 gnd.n3881 585
R11080 gnd.n3881 gnd.n3880 585
R11081 gnd.n2223 gnd.n2222 585
R11082 gnd.n3866 gnd.n2223 585
R11083 gnd.n3856 gnd.n2239 585
R11084 gnd.n2239 gnd.n2232 585
R11085 gnd.n3858 gnd.n3857 585
R11086 gnd.n3859 gnd.n3858 585
R11087 gnd.n3855 gnd.n2238 585
R11088 gnd.n2245 gnd.n2238 585
R11089 gnd.n3854 gnd.n3853 585
R11090 gnd.n3853 gnd.n3852 585
R11091 gnd.n2241 gnd.n2240 585
R11092 gnd.n3740 gnd.n2241 585
R11093 gnd.n3839 gnd.n3838 585
R11094 gnd.n3840 gnd.n3839 585
R11095 gnd.n3837 gnd.n2255 585
R11096 gnd.n2255 gnd.n2252 585
R11097 gnd.n3836 gnd.n3835 585
R11098 gnd.n3835 gnd.n3834 585
R11099 gnd.n2257 gnd.n2256 585
R11100 gnd.n3748 gnd.n2257 585
R11101 gnd.n3788 gnd.n3787 585
R11102 gnd.n3789 gnd.n3788 585
R11103 gnd.n3786 gnd.n2269 585
R11104 gnd.n2269 gnd.n2266 585
R11105 gnd.n3785 gnd.n3784 585
R11106 gnd.n3784 gnd.n3783 585
R11107 gnd.n2271 gnd.n2270 585
R11108 gnd.n3755 gnd.n2271 585
R11109 gnd.n3768 gnd.n3767 585
R11110 gnd.n3769 gnd.n3768 585
R11111 gnd.n3766 gnd.n2283 585
R11112 gnd.n3761 gnd.n2283 585
R11113 gnd.n3765 gnd.n3764 585
R11114 gnd.n3764 gnd.n3763 585
R11115 gnd.n2285 gnd.n2284 585
R11116 gnd.n3734 gnd.n2285 585
R11117 gnd.n3708 gnd.n3707 585
R11118 gnd.n3709 gnd.n3708 585
R11119 gnd.n3713 gnd.n3712 585
R11120 gnd.n3712 gnd.n3711 585
R11121 gnd.n3714 gnd.n2297 585
R11122 gnd.n3725 gnd.n2297 585
R11123 gnd.n3715 gnd.n2306 585
R11124 gnd.n3624 gnd.n2306 585
R11125 gnd.n3717 gnd.n3716 585
R11126 gnd.n3718 gnd.n3717 585
R11127 gnd.n3706 gnd.n2305 585
R11128 gnd.n3700 gnd.n2305 585
R11129 gnd.n3705 gnd.n3704 585
R11130 gnd.n3704 gnd.n3703 585
R11131 gnd.n2308 gnd.n2307 585
R11132 gnd.n3689 gnd.n2308 585
R11133 gnd.n3679 gnd.n2324 585
R11134 gnd.n2324 gnd.n2317 585
R11135 gnd.n3681 gnd.n3680 585
R11136 gnd.n3682 gnd.n3681 585
R11137 gnd.n3678 gnd.n2323 585
R11138 gnd.n2330 gnd.n2323 585
R11139 gnd.n3677 gnd.n3676 585
R11140 gnd.n3676 gnd.n3675 585
R11141 gnd.n2326 gnd.n2325 585
R11142 gnd.n2455 gnd.n2326 585
R11143 gnd.n3663 gnd.n3662 585
R11144 gnd.n3664 gnd.n3663 585
R11145 gnd.n3661 gnd.n2340 585
R11146 gnd.n2340 gnd.n2337 585
R11147 gnd.n3660 gnd.n3659 585
R11148 gnd.n3659 gnd.n3658 585
R11149 gnd.n2342 gnd.n2341 585
R11150 gnd.n2463 gnd.n2342 585
R11151 gnd.n3609 gnd.n3608 585
R11152 gnd.n3610 gnd.n3609 585
R11153 gnd.n3607 gnd.n2353 585
R11154 gnd.n2358 gnd.n2353 585
R11155 gnd.n3606 gnd.n3605 585
R11156 gnd.n3605 gnd.n3604 585
R11157 gnd.n2355 gnd.n2354 585
R11158 gnd.n2470 gnd.n2355 585
R11159 gnd.n3590 gnd.n3589 585
R11160 gnd.n3591 gnd.n3590 585
R11161 gnd.n3588 gnd.n2366 585
R11162 gnd.n3583 gnd.n2366 585
R11163 gnd.n3587 gnd.n3586 585
R11164 gnd.n3586 gnd.n3585 585
R11165 gnd.n2368 gnd.n2367 585
R11166 gnd.n2381 gnd.n2368 585
R11167 gnd.n2445 gnd.n2424 585
R11168 gnd.n2424 gnd.n2380 585
R11169 gnd.n3561 gnd.n3560 585
R11170 gnd.n3559 gnd.n2423 585
R11171 gnd.n3558 gnd.n2422 585
R11172 gnd.n3563 gnd.n2422 585
R11173 gnd.n3557 gnd.n3556 585
R11174 gnd.n3555 gnd.n3554 585
R11175 gnd.n3553 gnd.n3552 585
R11176 gnd.n3551 gnd.n3550 585
R11177 gnd.n3549 gnd.n3548 585
R11178 gnd.n3547 gnd.n3546 585
R11179 gnd.n3545 gnd.n3544 585
R11180 gnd.n3543 gnd.n3542 585
R11181 gnd.n3541 gnd.n3540 585
R11182 gnd.n3539 gnd.n3538 585
R11183 gnd.n3537 gnd.n3536 585
R11184 gnd.n3535 gnd.n3534 585
R11185 gnd.n3533 gnd.n3532 585
R11186 gnd.n3531 gnd.n3530 585
R11187 gnd.n3529 gnd.n3528 585
R11188 gnd.n3527 gnd.n3526 585
R11189 gnd.n3525 gnd.n3524 585
R11190 gnd.n3523 gnd.n3522 585
R11191 gnd.n3521 gnd.n3520 585
R11192 gnd.n3519 gnd.n3518 585
R11193 gnd.n3517 gnd.n3516 585
R11194 gnd.n3515 gnd.n3514 585
R11195 gnd.n3513 gnd.n3512 585
R11196 gnd.n3511 gnd.n3510 585
R11197 gnd.n3509 gnd.n3508 585
R11198 gnd.n3507 gnd.n3506 585
R11199 gnd.n3505 gnd.n3504 585
R11200 gnd.n3503 gnd.n3502 585
R11201 gnd.n3501 gnd.n3500 585
R11202 gnd.n3499 gnd.n3498 585
R11203 gnd.n3497 gnd.n2542 585
R11204 gnd.n2541 gnd.n2540 585
R11205 gnd.n2539 gnd.n2538 585
R11206 gnd.n2536 gnd.n2535 585
R11207 gnd.n2534 gnd.n2533 585
R11208 gnd.n2532 gnd.n2531 585
R11209 gnd.n2530 gnd.n2529 585
R11210 gnd.n2528 gnd.n2527 585
R11211 gnd.n2526 gnd.n2525 585
R11212 gnd.n2524 gnd.n2523 585
R11213 gnd.n2522 gnd.n2521 585
R11214 gnd.n2520 gnd.n2519 585
R11215 gnd.n2518 gnd.n2517 585
R11216 gnd.n2516 gnd.n2515 585
R11217 gnd.n2514 gnd.n2513 585
R11218 gnd.n2512 gnd.n2511 585
R11219 gnd.n2510 gnd.n2509 585
R11220 gnd.n2508 gnd.n2507 585
R11221 gnd.n2506 gnd.n2505 585
R11222 gnd.n2504 gnd.n2503 585
R11223 gnd.n2502 gnd.n2501 585
R11224 gnd.n2500 gnd.n2499 585
R11225 gnd.n2498 gnd.n2497 585
R11226 gnd.n2496 gnd.n2495 585
R11227 gnd.n2494 gnd.n2493 585
R11228 gnd.n2492 gnd.n2491 585
R11229 gnd.n2490 gnd.n2489 585
R11230 gnd.n2488 gnd.n2487 585
R11231 gnd.n2486 gnd.n2485 585
R11232 gnd.n2484 gnd.n2483 585
R11233 gnd.n2482 gnd.n2481 585
R11234 gnd.n2480 gnd.n2479 585
R11235 gnd.n4304 gnd.n4303 585
R11236 gnd.n4306 gnd.n4305 585
R11237 gnd.n4308 gnd.n4307 585
R11238 gnd.n4310 gnd.n4309 585
R11239 gnd.n4312 gnd.n4311 585
R11240 gnd.n4314 gnd.n4313 585
R11241 gnd.n4316 gnd.n4315 585
R11242 gnd.n4318 gnd.n4317 585
R11243 gnd.n4320 gnd.n4319 585
R11244 gnd.n4322 gnd.n4321 585
R11245 gnd.n4324 gnd.n4323 585
R11246 gnd.n4326 gnd.n4325 585
R11247 gnd.n4328 gnd.n4327 585
R11248 gnd.n4330 gnd.n4329 585
R11249 gnd.n4332 gnd.n4331 585
R11250 gnd.n4334 gnd.n4333 585
R11251 gnd.n4336 gnd.n4335 585
R11252 gnd.n4338 gnd.n4337 585
R11253 gnd.n4340 gnd.n4339 585
R11254 gnd.n4342 gnd.n4341 585
R11255 gnd.n4344 gnd.n4343 585
R11256 gnd.n4346 gnd.n4345 585
R11257 gnd.n4348 gnd.n4347 585
R11258 gnd.n4350 gnd.n4349 585
R11259 gnd.n4352 gnd.n4351 585
R11260 gnd.n4354 gnd.n4353 585
R11261 gnd.n4356 gnd.n4355 585
R11262 gnd.n4358 gnd.n4357 585
R11263 gnd.n4360 gnd.n4359 585
R11264 gnd.n4363 gnd.n4362 585
R11265 gnd.n4365 gnd.n4364 585
R11266 gnd.n4367 gnd.n4366 585
R11267 gnd.n4369 gnd.n4368 585
R11268 gnd.n4233 gnd.n2031 585
R11269 gnd.n4235 gnd.n4234 585
R11270 gnd.n4237 gnd.n4236 585
R11271 gnd.n4239 gnd.n4238 585
R11272 gnd.n4242 gnd.n4241 585
R11273 gnd.n4244 gnd.n4243 585
R11274 gnd.n4246 gnd.n4245 585
R11275 gnd.n4248 gnd.n4247 585
R11276 gnd.n4250 gnd.n4249 585
R11277 gnd.n4252 gnd.n4251 585
R11278 gnd.n4254 gnd.n4253 585
R11279 gnd.n4256 gnd.n4255 585
R11280 gnd.n4258 gnd.n4257 585
R11281 gnd.n4260 gnd.n4259 585
R11282 gnd.n4262 gnd.n4261 585
R11283 gnd.n4264 gnd.n4263 585
R11284 gnd.n4266 gnd.n4265 585
R11285 gnd.n4268 gnd.n4267 585
R11286 gnd.n4270 gnd.n4269 585
R11287 gnd.n4272 gnd.n4271 585
R11288 gnd.n4274 gnd.n4273 585
R11289 gnd.n4276 gnd.n4275 585
R11290 gnd.n4278 gnd.n4277 585
R11291 gnd.n4280 gnd.n4279 585
R11292 gnd.n4282 gnd.n4281 585
R11293 gnd.n4284 gnd.n4283 585
R11294 gnd.n4286 gnd.n4285 585
R11295 gnd.n4288 gnd.n4287 585
R11296 gnd.n4290 gnd.n4289 585
R11297 gnd.n4292 gnd.n4291 585
R11298 gnd.n4294 gnd.n4293 585
R11299 gnd.n4296 gnd.n4295 585
R11300 gnd.n4297 gnd.n2039 585
R11301 gnd.n4302 gnd.n2034 585
R11302 gnd.n4302 gnd.n4301 585
R11303 gnd.n4189 gnd.n2035 585
R11304 gnd.n4206 gnd.n2035 585
R11305 gnd.n4190 gnd.n2043 585
R11306 gnd.n4208 gnd.n2043 585
R11307 gnd.n4192 gnd.n4191 585
R11308 gnd.n4193 gnd.n4192 585
R11309 gnd.n4188 gnd.n2053 585
R11310 gnd.n2053 gnd.n2051 585
R11311 gnd.n4187 gnd.n4186 585
R11312 gnd.n4186 gnd.n4185 585
R11313 gnd.n2055 gnd.n2054 585
R11314 gnd.n2064 gnd.n2055 585
R11315 gnd.n4060 gnd.n2062 585
R11316 gnd.n4178 gnd.n2062 585
R11317 gnd.n4063 gnd.n4062 585
R11318 gnd.n4062 gnd.n4061 585
R11319 gnd.n4064 gnd.n2074 585
R11320 gnd.n4167 gnd.n2074 585
R11321 gnd.n4066 gnd.n4065 585
R11322 gnd.n4065 gnd.n2072 585
R11323 gnd.n4067 gnd.n2080 585
R11324 gnd.n4161 gnd.n2080 585
R11325 gnd.n4072 gnd.n4071 585
R11326 gnd.n4071 gnd.n4070 585
R11327 gnd.n4073 gnd.n2088 585
R11328 gnd.n4137 gnd.n2088 585
R11329 gnd.n4075 gnd.n4074 585
R11330 gnd.n4074 gnd.n2087 585
R11331 gnd.n4076 gnd.n2093 585
R11332 gnd.n4131 gnd.n2093 585
R11333 gnd.n4079 gnd.n4078 585
R11334 gnd.n4078 gnd.n4077 585
R11335 gnd.n4080 gnd.n2100 585
R11336 gnd.n4118 gnd.n2100 585
R11337 gnd.n4081 gnd.n2106 585
R11338 gnd.n4110 gnd.n2106 585
R11339 gnd.n4082 gnd.n2105 585
R11340 gnd.n4112 gnd.n2105 585
R11341 gnd.n4084 gnd.n4083 585
R11342 gnd.n4084 gnd.n2116 585
R11343 gnd.n4086 gnd.n4085 585
R11344 gnd.n4085 gnd.n2114 585
R11345 gnd.n4087 gnd.n2126 585
R11346 gnd.n4049 gnd.n2126 585
R11347 gnd.n4089 gnd.n4088 585
R11348 gnd.n4090 gnd.n4089 585
R11349 gnd.n4059 gnd.n2125 585
R11350 gnd.n2132 gnd.n2125 585
R11351 gnd.n4058 gnd.n4057 585
R11352 gnd.n4057 gnd.n4056 585
R11353 gnd.n2128 gnd.n2127 585
R11354 gnd.n4039 gnd.n2128 585
R11355 gnd.n4025 gnd.n2137 585
R11356 gnd.n4041 gnd.n2137 585
R11357 gnd.n4027 gnd.n4026 585
R11358 gnd.n4028 gnd.n4027 585
R11359 gnd.n4024 gnd.n2146 585
R11360 gnd.n2146 gnd.n2144 585
R11361 gnd.n4023 gnd.n4022 585
R11362 gnd.n4022 gnd.n4021 585
R11363 gnd.n2148 gnd.n2147 585
R11364 gnd.n2158 gnd.n2148 585
R11365 gnd.n3915 gnd.n2156 585
R11366 gnd.n4014 gnd.n2156 585
R11367 gnd.n3919 gnd.n3918 585
R11368 gnd.n3918 gnd.n3917 585
R11369 gnd.n3920 gnd.n2167 585
R11370 gnd.n4003 gnd.n2167 585
R11371 gnd.n3922 gnd.n3921 585
R11372 gnd.n3921 gnd.n2165 585
R11373 gnd.n3923 gnd.n2172 585
R11374 gnd.n3997 gnd.n2172 585
R11375 gnd.n3928 gnd.n3927 585
R11376 gnd.n3927 gnd.n3926 585
R11377 gnd.n3929 gnd.n2180 585
R11378 gnd.n3966 gnd.n2180 585
R11379 gnd.n3931 gnd.n3930 585
R11380 gnd.n3930 gnd.n2179 585
R11381 gnd.n3932 gnd.n2185 585
R11382 gnd.n3960 gnd.n2185 585
R11383 gnd.n3935 gnd.n3934 585
R11384 gnd.n3934 gnd.n3933 585
R11385 gnd.n3936 gnd.n2193 585
R11386 gnd.n3947 gnd.n2193 585
R11387 gnd.n3938 gnd.n3937 585
R11388 gnd.n3939 gnd.n3938 585
R11389 gnd.n3914 gnd.n2200 585
R11390 gnd.n3941 gnd.n2200 585
R11391 gnd.n3913 gnd.n3912 585
R11392 gnd.n3912 gnd.n3911 585
R11393 gnd.n2202 gnd.n2201 585
R11394 gnd.n3886 gnd.n2202 585
R11395 gnd.n3899 gnd.n2214 585
R11396 gnd.n3888 gnd.n2214 585
R11397 gnd.n3901 gnd.n3900 585
R11398 gnd.n3902 gnd.n3901 585
R11399 gnd.n3898 gnd.n2213 585
R11400 gnd.n2220 gnd.n2213 585
R11401 gnd.n3897 gnd.n3896 585
R11402 gnd.n3896 gnd.n3895 585
R11403 gnd.n2216 gnd.n2215 585
R11404 gnd.n3878 gnd.n2216 585
R11405 gnd.n3863 gnd.n2225 585
R11406 gnd.n3880 gnd.n2225 585
R11407 gnd.n3865 gnd.n3864 585
R11408 gnd.n3866 gnd.n3865 585
R11409 gnd.n3862 gnd.n2234 585
R11410 gnd.n2234 gnd.n2232 585
R11411 gnd.n3861 gnd.n3860 585
R11412 gnd.n3860 gnd.n3859 585
R11413 gnd.n2236 gnd.n2235 585
R11414 gnd.n2245 gnd.n2236 585
R11415 gnd.n3738 gnd.n2243 585
R11416 gnd.n3852 gnd.n2243 585
R11417 gnd.n3742 gnd.n3741 585
R11418 gnd.n3741 gnd.n3740 585
R11419 gnd.n3743 gnd.n2254 585
R11420 gnd.n3840 gnd.n2254 585
R11421 gnd.n3745 gnd.n3744 585
R11422 gnd.n3744 gnd.n2252 585
R11423 gnd.n3746 gnd.n2259 585
R11424 gnd.n3834 gnd.n2259 585
R11425 gnd.n3750 gnd.n3749 585
R11426 gnd.n3749 gnd.n3748 585
R11427 gnd.n3751 gnd.n2267 585
R11428 gnd.n3789 gnd.n2267 585
R11429 gnd.n3753 gnd.n3752 585
R11430 gnd.n3752 gnd.n2266 585
R11431 gnd.n3754 gnd.n2273 585
R11432 gnd.n3783 gnd.n2273 585
R11433 gnd.n3757 gnd.n3756 585
R11434 gnd.n3756 gnd.n3755 585
R11435 gnd.n3758 gnd.n2281 585
R11436 gnd.n3769 gnd.n2281 585
R11437 gnd.n3760 gnd.n3759 585
R11438 gnd.n3761 gnd.n3760 585
R11439 gnd.n3737 gnd.n2287 585
R11440 gnd.n3763 gnd.n2287 585
R11441 gnd.n3736 gnd.n3735 585
R11442 gnd.n3735 gnd.n3734 585
R11443 gnd.n2289 gnd.n2288 585
R11444 gnd.n3709 gnd.n2289 585
R11445 gnd.n3722 gnd.n2300 585
R11446 gnd.n3711 gnd.n2300 585
R11447 gnd.n3724 gnd.n3723 585
R11448 gnd.n3725 gnd.n3724 585
R11449 gnd.n3721 gnd.n2299 585
R11450 gnd.n3624 gnd.n2299 585
R11451 gnd.n3720 gnd.n3719 585
R11452 gnd.n3719 gnd.n3718 585
R11453 gnd.n2302 gnd.n2301 585
R11454 gnd.n3700 gnd.n2302 585
R11455 gnd.n3686 gnd.n2310 585
R11456 gnd.n3703 gnd.n2310 585
R11457 gnd.n3688 gnd.n3687 585
R11458 gnd.n3689 gnd.n3688 585
R11459 gnd.n3685 gnd.n2319 585
R11460 gnd.n2319 gnd.n2317 585
R11461 gnd.n3684 gnd.n3683 585
R11462 gnd.n3683 gnd.n3682 585
R11463 gnd.n2321 gnd.n2320 585
R11464 gnd.n2330 gnd.n2321 585
R11465 gnd.n2453 gnd.n2329 585
R11466 gnd.n3675 gnd.n2329 585
R11467 gnd.n2457 gnd.n2456 585
R11468 gnd.n2456 gnd.n2455 585
R11469 gnd.n2458 gnd.n2339 585
R11470 gnd.n3664 gnd.n2339 585
R11471 gnd.n2460 gnd.n2459 585
R11472 gnd.n2459 gnd.n2337 585
R11473 gnd.n2461 gnd.n2344 585
R11474 gnd.n3658 gnd.n2344 585
R11475 gnd.n2465 gnd.n2464 585
R11476 gnd.n2464 gnd.n2463 585
R11477 gnd.n2466 gnd.n2351 585
R11478 gnd.n3610 gnd.n2351 585
R11479 gnd.n2468 gnd.n2467 585
R11480 gnd.n2467 gnd.n2358 585
R11481 gnd.n2469 gnd.n2357 585
R11482 gnd.n3604 gnd.n2357 585
R11483 gnd.n2472 gnd.n2471 585
R11484 gnd.n2471 gnd.n2470 585
R11485 gnd.n2473 gnd.n2365 585
R11486 gnd.n3591 gnd.n2365 585
R11487 gnd.n2474 gnd.n2372 585
R11488 gnd.n3583 gnd.n2372 585
R11489 gnd.n2475 gnd.n2371 585
R11490 gnd.n3585 gnd.n2371 585
R11491 gnd.n2477 gnd.n2476 585
R11492 gnd.n2477 gnd.n2381 585
R11493 gnd.n2478 gnd.n2452 585
R11494 gnd.n2478 gnd.n2380 585
R11495 gnd.n2924 gnd.n2923 585
R11496 gnd.n2923 gnd.n1108 585
R11497 gnd.n7397 gnd.n7395 585
R11498 gnd.n7397 gnd.n7396 585
R11499 gnd.n7399 gnd.n7398 585
R11500 gnd.n7398 gnd.n225 585
R11501 gnd.n7400 gnd.n317 585
R11502 gnd.n317 gnd.n233 585
R11503 gnd.n7459 gnd.n7401 585
R11504 gnd.n7459 gnd.n7458 585
R11505 gnd.n7460 gnd.n316 585
R11506 gnd.n7460 gnd.n241 585
R11507 gnd.n7462 gnd.n7461 585
R11508 gnd.n7461 gnd.n239 585
R11509 gnd.n7463 gnd.n311 585
R11510 gnd.n311 gnd.n249 585
R11511 gnd.n7465 gnd.n7464 585
R11512 gnd.n7465 gnd.n247 585
R11513 gnd.n7466 gnd.n310 585
R11514 gnd.n7466 gnd.n257 585
R11515 gnd.n7468 gnd.n7467 585
R11516 gnd.n7467 gnd.n255 585
R11517 gnd.n7469 gnd.n307 585
R11518 gnd.n307 gnd.n264 585
R11519 gnd.n7472 gnd.n7471 585
R11520 gnd.n7473 gnd.n7472 585
R11521 gnd.n308 gnd.n306 585
R11522 gnd.n306 gnd.n296 585
R11523 gnd.n4654 gnd.n4653 585
R11524 gnd.n4653 gnd.n294 585
R11525 gnd.n4655 gnd.n4650 585
R11526 gnd.n4650 gnd.n4649 585
R11527 gnd.n4658 gnd.n4657 585
R11528 gnd.n4659 gnd.n4658 585
R11529 gnd.n4651 gnd.n1540 585
R11530 gnd.n1544 gnd.n1540 585
R11531 gnd.n4667 gnd.n4666 585
R11532 gnd.n4666 gnd.n4665 585
R11533 gnd.n4668 gnd.n1538 585
R11534 gnd.n4636 gnd.n1538 585
R11535 gnd.n4671 gnd.n4670 585
R11536 gnd.n4671 gnd.n280 585
R11537 gnd.n4672 gnd.n1537 585
R11538 gnd.n4672 gnd.n277 585
R11539 gnd.n4674 gnd.n4673 585
R11540 gnd.n4673 gnd.n1520 585
R11541 gnd.n4675 gnd.n1531 585
R11542 gnd.n1531 gnd.n1530 585
R11543 gnd.n4677 gnd.n4676 585
R11544 gnd.n4678 gnd.n4677 585
R11545 gnd.n1532 gnd.n1529 585
R11546 gnd.n4611 gnd.n1529 585
R11547 gnd.n4582 gnd.n4581 585
R11548 gnd.n4582 gnd.n1561 585
R11549 gnd.n4584 gnd.n4583 585
R11550 gnd.n4583 gnd.n1569 585
R11551 gnd.n4585 gnd.n1584 585
R11552 gnd.n1584 gnd.n1583 585
R11553 gnd.n4587 gnd.n4586 585
R11554 gnd.n4588 gnd.n4587 585
R11555 gnd.n1585 gnd.n1582 585
R11556 gnd.n1582 gnd.n1578 585
R11557 gnd.n4573 gnd.n4572 585
R11558 gnd.n4572 gnd.n4571 585
R11559 gnd.n1588 gnd.n1587 585
R11560 gnd.n1598 gnd.n1588 585
R11561 gnd.n4545 gnd.n1611 585
R11562 gnd.n1611 gnd.n1610 585
R11563 gnd.n4547 gnd.n4546 585
R11564 gnd.n4548 gnd.n4547 585
R11565 gnd.n1612 gnd.n1609 585
R11566 gnd.n1609 gnd.n1605 585
R11567 gnd.n4540 gnd.n4539 585
R11568 gnd.n4539 gnd.n4538 585
R11569 gnd.n1615 gnd.n1614 585
R11570 gnd.n4520 gnd.n1615 585
R11571 gnd.n1633 gnd.n1632 585
R11572 gnd.n1634 gnd.n1633 585
R11573 gnd.n1625 gnd.n1624 585
R11574 gnd.n1624 gnd.n1493 585
R11575 gnd.n1628 gnd.n1627 585
R11576 gnd.n1627 gnd.n1490 585
R11577 gnd.n1475 gnd.n1474 585
R11578 gnd.n1480 gnd.n1475 585
R11579 gnd.n4727 gnd.n4726 585
R11580 gnd.n4726 gnd.n4725 585
R11581 gnd.n4728 gnd.n1469 585
R11582 gnd.n1476 gnd.n1469 585
R11583 gnd.n4730 gnd.n4729 585
R11584 gnd.n4731 gnd.n4730 585
R11585 gnd.n1466 gnd.n1465 585
R11586 gnd.n4732 gnd.n1466 585
R11587 gnd.n4735 gnd.n4734 585
R11588 gnd.n4734 gnd.n4733 585
R11589 gnd.n4736 gnd.n1460 585
R11590 gnd.n1460 gnd.n1458 585
R11591 gnd.n4738 gnd.n4737 585
R11592 gnd.n4739 gnd.n4738 585
R11593 gnd.n1461 gnd.n1459 585
R11594 gnd.n1459 gnd.n1456 585
R11595 gnd.n4451 gnd.n4450 585
R11596 gnd.n4452 gnd.n4451 585
R11597 gnd.n1804 gnd.n1803 585
R11598 gnd.n4441 gnd.n1803 585
R11599 gnd.n4445 gnd.n4444 585
R11600 gnd.n4444 gnd.n4443 585
R11601 gnd.n1807 gnd.n1806 585
R11602 gnd.n4429 gnd.n1807 585
R11603 gnd.n4427 gnd.n4426 585
R11604 gnd.n4428 gnd.n4427 585
R11605 gnd.n1817 gnd.n1816 585
R11606 gnd.n4418 gnd.n1816 585
R11607 gnd.n4422 gnd.n4421 585
R11608 gnd.n4421 gnd.n4420 585
R11609 gnd.n1820 gnd.n1819 585
R11610 gnd.n4409 gnd.n1820 585
R11611 gnd.n4407 gnd.n4406 585
R11612 gnd.n4408 gnd.n4407 585
R11613 gnd.n1830 gnd.n1829 585
R11614 gnd.n4398 gnd.n1829 585
R11615 gnd.n4402 gnd.n4401 585
R11616 gnd.n4401 gnd.n4400 585
R11617 gnd.n1833 gnd.n1832 585
R11618 gnd.n4389 gnd.n1833 585
R11619 gnd.n4387 gnd.n4386 585
R11620 gnd.n4388 gnd.n4387 585
R11621 gnd.n1843 gnd.n1842 585
R11622 gnd.n4378 gnd.n1842 585
R11623 gnd.n4382 gnd.n4381 585
R11624 gnd.n4381 gnd.n4380 585
R11625 gnd.n1846 gnd.n1845 585
R11626 gnd.n1871 gnd.n1846 585
R11627 gnd.n4202 gnd.n2046 585
R11628 gnd.n2046 gnd.n1852 585
R11629 gnd.n4204 gnd.n4203 585
R11630 gnd.n4205 gnd.n4204 585
R11631 gnd.n2047 gnd.n2045 585
R11632 gnd.n2045 gnd.n2042 585
R11633 gnd.n4197 gnd.n4196 585
R11634 gnd.n4196 gnd.n4195 585
R11635 gnd.n2050 gnd.n2049 585
R11636 gnd.n2063 gnd.n2050 585
R11637 gnd.n4176 gnd.n4175 585
R11638 gnd.n4177 gnd.n4176 585
R11639 gnd.n2068 gnd.n2067 585
R11640 gnd.n2075 gnd.n2067 585
R11641 gnd.n4171 gnd.n4170 585
R11642 gnd.n4170 gnd.n4169 585
R11643 gnd.n2071 gnd.n2070 585
R11644 gnd.n2079 gnd.n2071 585
R11645 gnd.n4126 gnd.n2095 585
R11646 gnd.n2095 gnd.n2089 585
R11647 gnd.n4128 gnd.n4127 585
R11648 gnd.n4129 gnd.n4128 585
R11649 gnd.n2096 gnd.n2094 585
R11650 gnd.n2094 gnd.t180 585
R11651 gnd.n4121 gnd.n4120 585
R11652 gnd.n4120 gnd.n4119 585
R11653 gnd.n2099 gnd.n2098 585
R11654 gnd.n4111 gnd.n2099 585
R11655 gnd.n4097 gnd.n4096 585
R11656 gnd.n4098 gnd.n4097 585
R11657 gnd.n2118 gnd.n2117 585
R11658 gnd.n4048 gnd.n2117 585
R11659 gnd.n4092 gnd.n4091 585
R11660 gnd.n4091 gnd.n4090 585
R11661 gnd.n2121 gnd.n2120 585
R11662 gnd.n2130 gnd.n2121 585
R11663 gnd.n4037 gnd.n4036 585
R11664 gnd.n4038 gnd.n4037 585
R11665 gnd.n2140 gnd.n2139 585
R11666 gnd.n2139 gnd.n2136 585
R11667 gnd.n4032 gnd.n4031 585
R11668 gnd.n4031 gnd.n4030 585
R11669 gnd.n2143 gnd.n2142 585
R11670 gnd.n2157 gnd.n2143 585
R11671 gnd.n4012 gnd.n4011 585
R11672 gnd.n4013 gnd.n4012 585
R11673 gnd.n2161 gnd.n2160 585
R11674 gnd.n3916 gnd.n2160 585
R11675 gnd.n4007 gnd.n4006 585
R11676 gnd.n4006 gnd.n4005 585
R11677 gnd.n2164 gnd.n2163 585
R11678 gnd.n2171 gnd.n2164 585
R11679 gnd.n3955 gnd.n2187 585
R11680 gnd.n3924 gnd.n2187 585
R11681 gnd.n3957 gnd.n3956 585
R11682 gnd.n3958 gnd.n3957 585
R11683 gnd.n2188 gnd.n2186 585
R11684 gnd.n2186 gnd.n2184 585
R11685 gnd.n3950 gnd.n3949 585
R11686 gnd.n3949 gnd.n3948 585
R11687 gnd.n2191 gnd.n2190 585
R11688 gnd.n3940 gnd.n2191 585
R11689 gnd.n3909 gnd.n3908 585
R11690 gnd.n3910 gnd.n3909 585
R11691 gnd.n2205 gnd.n2204 585
R11692 gnd.n3887 gnd.n2204 585
R11693 gnd.n3904 gnd.n3903 585
R11694 gnd.n3903 gnd.n3902 585
R11695 gnd.n2208 gnd.n2207 585
R11696 gnd.n2218 gnd.n2208 585
R11697 gnd.n3876 gnd.n3875 585
R11698 gnd.n3877 gnd.n3876 585
R11699 gnd.n2228 gnd.n2227 585
R11700 gnd.n2227 gnd.n2224 585
R11701 gnd.n3871 gnd.n3870 585
R11702 gnd.n3870 gnd.n3869 585
R11703 gnd.n2231 gnd.n2230 585
R11704 gnd.n2244 gnd.n2231 585
R11705 gnd.n3850 gnd.n3849 585
R11706 gnd.n3851 gnd.n3850 585
R11707 gnd.n2248 gnd.n2247 585
R11708 gnd.n3739 gnd.n2247 585
R11709 gnd.n3845 gnd.n3844 585
R11710 gnd.n3844 gnd.n3843 585
R11711 gnd.n2251 gnd.n2250 585
R11712 gnd.n2258 gnd.n2251 585
R11713 gnd.n3777 gnd.n2275 585
R11714 gnd.n2275 gnd.n2268 585
R11715 gnd.n3779 gnd.n3778 585
R11716 gnd.n3780 gnd.n3779 585
R11717 gnd.n2276 gnd.n2274 585
R11718 gnd.n2274 gnd.n2272 585
R11719 gnd.n3772 gnd.n3771 585
R11720 gnd.n3771 gnd.n3770 585
R11721 gnd.n2279 gnd.n2278 585
R11722 gnd.n3762 gnd.n2279 585
R11723 gnd.n3732 gnd.n3731 585
R11724 gnd.n3733 gnd.n3732 585
R11725 gnd.n2293 gnd.n2292 585
R11726 gnd.n3710 gnd.n2292 585
R11727 gnd.n3727 gnd.n3726 585
R11728 gnd.n3726 gnd.n3725 585
R11729 gnd.n2296 gnd.n2295 585
R11730 gnd.n2304 gnd.n2296 585
R11731 gnd.n3698 gnd.n3697 585
R11732 gnd.n3699 gnd.n3698 585
R11733 gnd.n2313 gnd.n2312 585
R11734 gnd.n2312 gnd.n2309 585
R11735 gnd.n3693 gnd.n3692 585
R11736 gnd.n3692 gnd.n3691 585
R11737 gnd.n2316 gnd.n2315 585
R11738 gnd.t298 gnd.n2316 585
R11739 gnd.n3673 gnd.n3672 585
R11740 gnd.n3674 gnd.n3673 585
R11741 gnd.n2333 gnd.n2332 585
R11742 gnd.n2454 gnd.n2332 585
R11743 gnd.n3668 gnd.n3667 585
R11744 gnd.n3667 gnd.n3666 585
R11745 gnd.n2336 gnd.n2335 585
R11746 gnd.n2343 gnd.n2336 585
R11747 gnd.n3599 gnd.n2360 585
R11748 gnd.n2360 gnd.n2352 585
R11749 gnd.n3601 gnd.n3600 585
R11750 gnd.n3602 gnd.n3601 585
R11751 gnd.n2361 gnd.n2359 585
R11752 gnd.n2359 gnd.n2356 585
R11753 gnd.n3594 gnd.n3593 585
R11754 gnd.n3593 gnd.n3592 585
R11755 gnd.n2364 gnd.n2363 585
R11756 gnd.n3584 gnd.n2364 585
R11757 gnd.n3571 gnd.n3570 585
R11758 gnd.n3572 gnd.n3571 585
R11759 gnd.n2383 gnd.n2382 585
R11760 gnd.n2420 gnd.n2382 585
R11761 gnd.n3566 gnd.n3565 585
R11762 gnd.n3565 gnd.n3564 585
R11763 gnd.n2386 gnd.n2385 585
R11764 gnd.n3397 gnd.n2386 585
R11765 gnd.n3395 gnd.n3394 585
R11766 gnd.n3396 gnd.n3395 585
R11767 gnd.n2686 gnd.n2685 585
R11768 gnd.n3386 gnd.n2685 585
R11769 gnd.n3390 gnd.n3389 585
R11770 gnd.n3389 gnd.n3388 585
R11771 gnd.n2689 gnd.n2688 585
R11772 gnd.n3384 gnd.n2689 585
R11773 gnd.n3379 gnd.n3378 585
R11774 gnd.n3380 gnd.n3379 585
R11775 gnd.n2692 gnd.n2691 585
R11776 gnd.n3370 gnd.n2691 585
R11777 gnd.n3374 gnd.n3373 585
R11778 gnd.n3373 gnd.n3372 585
R11779 gnd.n2695 gnd.n2694 585
R11780 gnd.n3368 gnd.n2695 585
R11781 gnd.n3363 gnd.n3362 585
R11782 gnd.n3364 gnd.n3363 585
R11783 gnd.n2698 gnd.n2697 585
R11784 gnd.n3354 gnd.n2697 585
R11785 gnd.n3358 gnd.n3357 585
R11786 gnd.n3357 gnd.n3356 585
R11787 gnd.n2701 gnd.n2700 585
R11788 gnd.n3352 gnd.n2701 585
R11789 gnd.n3347 gnd.n3346 585
R11790 gnd.n3348 gnd.n3347 585
R11791 gnd.n2704 gnd.n2703 585
R11792 gnd.n3338 gnd.n2703 585
R11793 gnd.n3342 gnd.n3341 585
R11794 gnd.n3341 gnd.n3340 585
R11795 gnd.n2707 gnd.n2706 585
R11796 gnd.n3336 gnd.n2707 585
R11797 gnd.n3334 gnd.n3333 585
R11798 gnd.n3335 gnd.n3334 585
R11799 gnd.n2842 gnd.n2841 585
R11800 gnd.n3326 gnd.n2841 585
R11801 gnd.n3329 gnd.n3328 585
R11802 gnd.n3328 gnd.n3327 585
R11803 gnd.n3324 gnd.n2844 585
R11804 gnd.n3325 gnd.n3324 585
R11805 gnd.n3323 gnd.n3322 585
R11806 gnd.n3323 gnd.n1323 585
R11807 gnd.n2846 gnd.n2845 585
R11808 gnd.n2845 gnd.n1320 585
R11809 gnd.n3318 gnd.n3317 585
R11810 gnd.n3317 gnd.n2641 585
R11811 gnd.n3316 gnd.n2848 585
R11812 gnd.n3316 gnd.n1311 585
R11813 gnd.n3315 gnd.n3314 585
R11814 gnd.n3315 gnd.n1303 585
R11815 gnd.n2850 gnd.n2849 585
R11816 gnd.n2849 gnd.n1300 585
R11817 gnd.n3310 gnd.n3309 585
R11818 gnd.n3309 gnd.n1292 585
R11819 gnd.n3308 gnd.n2852 585
R11820 gnd.n3308 gnd.n1289 585
R11821 gnd.n3307 gnd.n3306 585
R11822 gnd.n3307 gnd.n1281 585
R11823 gnd.n2854 gnd.n2853 585
R11824 gnd.n2853 gnd.n1278 585
R11825 gnd.n3302 gnd.n3301 585
R11826 gnd.n3301 gnd.n3300 585
R11827 gnd.n2857 gnd.n2856 585
R11828 gnd.n2857 gnd.n1268 585
R11829 gnd.n2962 gnd.n2961 585
R11830 gnd.n2962 gnd.n2872 585
R11831 gnd.n2964 gnd.n2963 585
R11832 gnd.n2963 gnd.n1258 585
R11833 gnd.n2965 gnd.n2955 585
R11834 gnd.n2955 gnd.n1250 585
R11835 gnd.n2967 gnd.n2966 585
R11836 gnd.n2967 gnd.n1247 585
R11837 gnd.n2968 gnd.n2954 585
R11838 gnd.n2968 gnd.n1239 585
R11839 gnd.n2970 gnd.n2969 585
R11840 gnd.n2969 gnd.n1236 585
R11841 gnd.n2971 gnd.n2949 585
R11842 gnd.n2949 gnd.n2882 585
R11843 gnd.n2973 gnd.n2972 585
R11844 gnd.n2973 gnd.n1226 585
R11845 gnd.n2974 gnd.n2948 585
R11846 gnd.n2974 gnd.n2886 585
R11847 gnd.n2976 gnd.n2975 585
R11848 gnd.n2975 gnd.n1216 585
R11849 gnd.n2977 gnd.n2946 585
R11850 gnd.n2946 gnd.n1209 585
R11851 gnd.n2979 gnd.n2978 585
R11852 gnd.n2979 gnd.n1206 585
R11853 gnd.n2981 gnd.n2980 585
R11854 gnd.n2980 gnd.n1198 585
R11855 gnd.n2983 gnd.n2982 585
R11856 gnd.n2983 gnd.n1195 585
R11857 gnd.n2985 gnd.n2984 585
R11858 gnd.n2984 gnd.n2896 585
R11859 gnd.n2987 gnd.n2986 585
R11860 gnd.n2987 gnd.n1188 585
R11861 gnd.n2989 gnd.n2988 585
R11862 gnd.n2989 gnd.n2901 585
R11863 gnd.n2990 gnd.n2945 585
R11864 gnd.n2990 gnd.n1178 585
R11865 gnd.n2992 gnd.n2991 585
R11866 gnd.n2991 gnd.n1172 585
R11867 gnd.n2940 gnd.n2939 585
R11868 gnd.n2939 gnd.n1169 585
R11869 gnd.n2998 gnd.n2997 585
R11870 gnd.n2998 gnd.n1161 585
R11871 gnd.n2999 gnd.n2938 585
R11872 gnd.n2999 gnd.n1158 585
R11873 gnd.n3001 gnd.n3000 585
R11874 gnd.n3000 gnd.n2911 585
R11875 gnd.n3002 gnd.n2916 585
R11876 gnd.n2916 gnd.n1148 585
R11877 gnd.n3004 gnd.n3003 585
R11878 gnd.n3005 gnd.n3004 585
R11879 gnd.n2917 gnd.n2915 585
R11880 gnd.n2915 gnd.n1138 585
R11881 gnd.n2932 gnd.n2931 585
R11882 gnd.n2931 gnd.n1130 585
R11883 gnd.n2930 gnd.n2919 585
R11884 gnd.n2930 gnd.n1127 585
R11885 gnd.n2929 gnd.n2928 585
R11886 gnd.n2929 gnd.n1119 585
R11887 gnd.n2921 gnd.n2920 585
R11888 gnd.n2920 gnd.n1116 585
R11889 gnd.n4742 gnd.n4741 585
R11890 gnd.n4741 gnd.n4740 585
R11891 gnd.n4743 gnd.n1454 585
R11892 gnd.n4453 gnd.n1454 585
R11893 gnd.n4439 gnd.n1452 585
R11894 gnd.n4440 gnd.n4439 585
R11895 gnd.n4747 gnd.n1451 585
R11896 gnd.n4442 gnd.n1451 585
R11897 gnd.n4748 gnd.n1450 585
R11898 gnd.n1808 gnd.n1450 585
R11899 gnd.n4749 gnd.n1449 585
R11900 gnd.n4430 gnd.n1449 585
R11901 gnd.n1814 gnd.n1447 585
R11902 gnd.n1815 gnd.n1814 585
R11903 gnd.n4753 gnd.n1446 585
R11904 gnd.n4419 gnd.n1446 585
R11905 gnd.n4754 gnd.n1445 585
R11906 gnd.n1821 gnd.n1445 585
R11907 gnd.n4755 gnd.n1444 585
R11908 gnd.n4410 gnd.n1444 585
R11909 gnd.n1827 gnd.n1442 585
R11910 gnd.n1828 gnd.n1827 585
R11911 gnd.n4759 gnd.n1441 585
R11912 gnd.n4399 gnd.n1441 585
R11913 gnd.n4760 gnd.n1440 585
R11914 gnd.n1834 gnd.n1440 585
R11915 gnd.n4761 gnd.n1439 585
R11916 gnd.n4390 gnd.n1439 585
R11917 gnd.n1840 gnd.n1437 585
R11918 gnd.n1841 gnd.n1840 585
R11919 gnd.n4765 gnd.n1436 585
R11920 gnd.n4379 gnd.n1436 585
R11921 gnd.n4766 gnd.n1435 585
R11922 gnd.n1870 gnd.n1435 585
R11923 gnd.n4767 gnd.n1434 585
R11924 gnd.n4370 gnd.n1434 585
R11925 gnd.n2036 gnd.n1432 585
R11926 gnd.n2037 gnd.n2036 585
R11927 gnd.n4771 gnd.n1431 585
R11928 gnd.n4207 gnd.n1431 585
R11929 gnd.n4772 gnd.n1430 585
R11930 gnd.n4194 gnd.n1430 585
R11931 gnd.n4773 gnd.n1429 585
R11932 gnd.n2056 gnd.n1429 585
R11933 gnd.n2065 gnd.n1427 585
R11934 gnd.n2066 gnd.n2065 585
R11935 gnd.n4777 gnd.n1426 585
R11936 gnd.n2061 gnd.n1426 585
R11937 gnd.n4778 gnd.n1425 585
R11938 gnd.n4168 gnd.n1425 585
R11939 gnd.n4779 gnd.n1424 585
R11940 gnd.n4160 gnd.n1424 585
R11941 gnd.n4068 gnd.n1422 585
R11942 gnd.n4069 gnd.n4068 585
R11943 gnd.n4783 gnd.n1421 585
R11944 gnd.n4138 gnd.n1421 585
R11945 gnd.n4784 gnd.n1420 585
R11946 gnd.n4130 gnd.n1420 585
R11947 gnd.n4785 gnd.n1419 585
R11948 gnd.n2101 gnd.n1419 585
R11949 gnd.n4108 gnd.n1417 585
R11950 gnd.n4109 gnd.n4108 585
R11951 gnd.n4789 gnd.n1416 585
R11952 gnd.n2115 gnd.n1416 585
R11953 gnd.n4790 gnd.n1415 585
R11954 gnd.n4099 gnd.n1415 585
R11955 gnd.n4791 gnd.n1414 585
R11956 gnd.n4047 gnd.n1414 585
R11957 gnd.n2122 gnd.n1412 585
R11958 gnd.n2123 gnd.n2122 585
R11959 gnd.n4795 gnd.n1411 585
R11960 gnd.n2129 gnd.n1411 585
R11961 gnd.n4796 gnd.n1410 585
R11962 gnd.n4040 gnd.n1410 585
R11963 gnd.n4797 gnd.n1409 585
R11964 gnd.n4029 gnd.n1409 585
R11965 gnd.n2149 gnd.n1407 585
R11966 gnd.n2150 gnd.n2149 585
R11967 gnd.n4801 gnd.n1406 585
R11968 gnd.n2159 gnd.n1406 585
R11969 gnd.n4802 gnd.n1405 585
R11970 gnd.n2155 gnd.n1405 585
R11971 gnd.n4803 gnd.n1404 585
R11972 gnd.n4004 gnd.n1404 585
R11973 gnd.n3995 gnd.n1402 585
R11974 gnd.n3996 gnd.n3995 585
R11975 gnd.n4807 gnd.n1401 585
R11976 gnd.n3925 gnd.n1401 585
R11977 gnd.n4808 gnd.n1400 585
R11978 gnd.n3967 gnd.n1400 585
R11979 gnd.n4809 gnd.n1399 585
R11980 gnd.n3959 gnd.n1399 585
R11981 gnd.n2194 gnd.n1397 585
R11982 gnd.n2195 gnd.n2194 585
R11983 gnd.n4813 gnd.n1396 585
R11984 gnd.n2192 gnd.n1396 585
R11985 gnd.n4814 gnd.n1395 585
R11986 gnd.n2199 gnd.n1395 585
R11987 gnd.n4815 gnd.n1394 585
R11988 gnd.n2203 gnd.n1394 585
R11989 gnd.n2211 gnd.n1392 585
R11990 gnd.n2212 gnd.n2211 585
R11991 gnd.n4819 gnd.n1391 585
R11992 gnd.n2209 gnd.n1391 585
R11993 gnd.n4820 gnd.n1390 585
R11994 gnd.n2217 gnd.n1390 585
R11995 gnd.n4821 gnd.n1389 585
R11996 gnd.n3879 gnd.n1389 585
R11997 gnd.n3867 gnd.n1387 585
R11998 gnd.n3868 gnd.n3867 585
R11999 gnd.n4825 gnd.n1386 585
R12000 gnd.n2237 gnd.n1386 585
R12001 gnd.n4826 gnd.n1385 585
R12002 gnd.n2246 gnd.n1385 585
R12003 gnd.n4827 gnd.n1384 585
R12004 gnd.n2242 gnd.n1384 585
R12005 gnd.n3841 gnd.n1382 585
R12006 gnd.n3842 gnd.n3841 585
R12007 gnd.n4831 gnd.n1381 585
R12008 gnd.n3833 gnd.n1381 585
R12009 gnd.n4832 gnd.n1380 585
R12010 gnd.n3747 gnd.n1380 585
R12011 gnd.n4833 gnd.n1379 585
R12012 gnd.n3790 gnd.n1379 585
R12013 gnd.n3781 gnd.n1377 585
R12014 gnd.n3782 gnd.n3781 585
R12015 gnd.n4837 gnd.n1376 585
R12016 gnd.n2282 gnd.n1376 585
R12017 gnd.n4838 gnd.n1375 585
R12018 gnd.n2280 gnd.n1375 585
R12019 gnd.n4839 gnd.n1374 585
R12020 gnd.n2286 gnd.n1374 585
R12021 gnd.n2290 gnd.n1372 585
R12022 gnd.n2291 gnd.n2290 585
R12023 gnd.n4843 gnd.n1371 585
R12024 gnd.n2298 gnd.n1371 585
R12025 gnd.n4844 gnd.n1370 585
R12026 gnd.n3625 gnd.n1370 585
R12027 gnd.n4845 gnd.n1369 585
R12028 gnd.n2303 gnd.n1369 585
R12029 gnd.n3701 gnd.n1367 585
R12030 gnd.n3702 gnd.n3701 585
R12031 gnd.n4849 gnd.n1366 585
R12032 gnd.n3690 gnd.n1366 585
R12033 gnd.n4850 gnd.n1365 585
R12034 gnd.n2322 gnd.n1365 585
R12035 gnd.n4851 gnd.n1364 585
R12036 gnd.n2331 gnd.n1364 585
R12037 gnd.n2327 gnd.n1362 585
R12038 gnd.n2328 gnd.n2327 585
R12039 gnd.n4855 gnd.n1361 585
R12040 gnd.n3665 gnd.n1361 585
R12041 gnd.n4856 gnd.n1360 585
R12042 gnd.n3657 gnd.n1360 585
R12043 gnd.n4857 gnd.n1359 585
R12044 gnd.n2462 gnd.n1359 585
R12045 gnd.n3611 gnd.n1357 585
R12046 gnd.n3612 gnd.n3611 585
R12047 gnd.n4861 gnd.n1356 585
R12048 gnd.n3603 gnd.n1356 585
R12049 gnd.n4862 gnd.n1355 585
R12050 gnd.t245 gnd.n1355 585
R12051 gnd.n4863 gnd.n1354 585
R12052 gnd.n3582 gnd.n1354 585
R12053 gnd.n2369 gnd.n1352 585
R12054 gnd.n2370 gnd.n2369 585
R12055 gnd.n4867 gnd.n1351 585
R12056 gnd.n3573 gnd.n1351 585
R12057 gnd.n4868 gnd.n1350 585
R12058 gnd.n2421 gnd.n1350 585
R12059 gnd.n4869 gnd.n1349 585
R12060 gnd.n2387 gnd.n1349 585
R12061 gnd.n3398 gnd.n1347 585
R12062 gnd.n3399 gnd.n3398 585
R12063 gnd.n4873 gnd.n1346 585
R12064 gnd.n2684 gnd.n1346 585
R12065 gnd.n4874 gnd.n1345 585
R12066 gnd.n3387 gnd.n1345 585
R12067 gnd.n4875 gnd.n1344 585
R12068 gnd.n3385 gnd.n1344 585
R12069 gnd.n3382 gnd.n1342 585
R12070 gnd.n3383 gnd.n3382 585
R12071 gnd.n4879 gnd.n1341 585
R12072 gnd.n2690 gnd.n1341 585
R12073 gnd.n4880 gnd.n1340 585
R12074 gnd.n3371 gnd.n1340 585
R12075 gnd.n4881 gnd.n1339 585
R12076 gnd.n3369 gnd.n1339 585
R12077 gnd.n3366 gnd.n1337 585
R12078 gnd.n3367 gnd.n3366 585
R12079 gnd.n4885 gnd.n1336 585
R12080 gnd.n2696 gnd.n1336 585
R12081 gnd.n4886 gnd.n1335 585
R12082 gnd.n3355 gnd.n1335 585
R12083 gnd.n4887 gnd.n1334 585
R12084 gnd.n3353 gnd.n1334 585
R12085 gnd.n3350 gnd.n1332 585
R12086 gnd.n3351 gnd.n3350 585
R12087 gnd.n4891 gnd.n1331 585
R12088 gnd.n2702 gnd.n1331 585
R12089 gnd.n4892 gnd.n1330 585
R12090 gnd.n3339 gnd.n1330 585
R12091 gnd.n4893 gnd.n1329 585
R12092 gnd.n3337 gnd.n1329 585
R12093 gnd.n2838 gnd.n2837 585
R12094 gnd.n2836 gnd.n2724 585
R12095 gnd.n2726 gnd.n2723 585
R12096 gnd.n2840 gnd.n2723 585
R12097 gnd.n2829 gnd.n2739 585
R12098 gnd.n2828 gnd.n2740 585
R12099 gnd.n2742 gnd.n2741 585
R12100 gnd.n2821 gnd.n2750 585
R12101 gnd.n2820 gnd.n2751 585
R12102 gnd.n2761 gnd.n2752 585
R12103 gnd.n2813 gnd.n2762 585
R12104 gnd.n2812 gnd.n2763 585
R12105 gnd.n2765 gnd.n2764 585
R12106 gnd.n2805 gnd.n2773 585
R12107 gnd.n2804 gnd.n2774 585
R12108 gnd.n2786 gnd.n2775 585
R12109 gnd.n2797 gnd.n2787 585
R12110 gnd.n2796 gnd.n2789 585
R12111 gnd.n2788 gnd.n2647 585
R12112 gnd.n3443 gnd.n2648 585
R12113 gnd.n3442 gnd.n2649 585
R12114 gnd.n3441 gnd.n2650 585
R12115 gnd.n2717 gnd.n2651 585
R12116 gnd.n3437 gnd.n2653 585
R12117 gnd.n3436 gnd.n2654 585
R12118 gnd.n3435 gnd.n2655 585
R12119 gnd.n3432 gnd.n2660 585
R12120 gnd.n3431 gnd.n2661 585
R12121 gnd.n3430 gnd.n2662 585
R12122 gnd.n2721 gnd.n2663 585
R12123 gnd.n4456 gnd.n1457 585
R12124 gnd.n4740 gnd.n1457 585
R12125 gnd.n4455 gnd.n4454 585
R12126 gnd.n4454 gnd.n4453 585
R12127 gnd.n1802 gnd.n1801 585
R12128 gnd.n4440 gnd.n1802 585
R12129 gnd.n4438 gnd.n4437 585
R12130 gnd.n4442 gnd.n4438 585
R12131 gnd.n1810 gnd.n1809 585
R12132 gnd.n1809 gnd.n1808 585
R12133 gnd.n4432 gnd.n4431 585
R12134 gnd.n4431 gnd.n4430 585
R12135 gnd.n1813 gnd.n1812 585
R12136 gnd.n1815 gnd.n1813 585
R12137 gnd.n4417 gnd.n4416 585
R12138 gnd.n4419 gnd.n4417 585
R12139 gnd.n1823 gnd.n1822 585
R12140 gnd.n1822 gnd.n1821 585
R12141 gnd.n4412 gnd.n4411 585
R12142 gnd.n4411 gnd.n4410 585
R12143 gnd.n1826 gnd.n1825 585
R12144 gnd.n1828 gnd.n1826 585
R12145 gnd.n4397 gnd.n4396 585
R12146 gnd.n4399 gnd.n4397 585
R12147 gnd.n1836 gnd.n1835 585
R12148 gnd.n1835 gnd.n1834 585
R12149 gnd.n4392 gnd.n4391 585
R12150 gnd.n4391 gnd.n4390 585
R12151 gnd.n1839 gnd.n1838 585
R12152 gnd.n1841 gnd.n1839 585
R12153 gnd.n4377 gnd.n4376 585
R12154 gnd.n4379 gnd.n4377 585
R12155 gnd.n1848 gnd.n1847 585
R12156 gnd.n1870 gnd.n1847 585
R12157 gnd.n4372 gnd.n4371 585
R12158 gnd.n4371 gnd.n4370 585
R12159 gnd.n1851 gnd.n1850 585
R12160 gnd.n2037 gnd.n1851 585
R12161 gnd.n4148 gnd.n2044 585
R12162 gnd.n4207 gnd.n2044 585
R12163 gnd.n4147 gnd.n2052 585
R12164 gnd.n4194 gnd.n2052 585
R12165 gnd.n4152 gnd.n4146 585
R12166 gnd.n4146 gnd.n2056 585
R12167 gnd.n4153 gnd.n4145 585
R12168 gnd.n4145 gnd.n2066 585
R12169 gnd.n4154 gnd.n4144 585
R12170 gnd.n4144 gnd.n2061 585
R12171 gnd.n2083 gnd.n2073 585
R12172 gnd.n4168 gnd.n2073 585
R12173 gnd.n4159 gnd.n4158 585
R12174 gnd.n4160 gnd.n4159 585
R12175 gnd.n2082 gnd.n2081 585
R12176 gnd.n4069 gnd.n2081 585
R12177 gnd.n4140 gnd.n4139 585
R12178 gnd.n4139 gnd.n4138 585
R12179 gnd.n2086 gnd.n2085 585
R12180 gnd.n4130 gnd.n2086 585
R12181 gnd.n2110 gnd.n2108 585
R12182 gnd.n2108 gnd.n2101 585
R12183 gnd.n4107 gnd.n4106 585
R12184 gnd.n4109 gnd.n4107 585
R12185 gnd.n2109 gnd.n2107 585
R12186 gnd.n2115 gnd.n2107 585
R12187 gnd.n4101 gnd.n4100 585
R12188 gnd.n4100 gnd.n4099 585
R12189 gnd.n2113 gnd.n2112 585
R12190 gnd.n4047 gnd.n2113 585
R12191 gnd.n3981 gnd.n3979 585
R12192 gnd.n3979 gnd.n2123 585
R12193 gnd.n3982 gnd.n3978 585
R12194 gnd.n3978 gnd.n2129 585
R12195 gnd.n3983 gnd.n2138 585
R12196 gnd.n4040 gnd.n2138 585
R12197 gnd.n3976 gnd.n2145 585
R12198 gnd.n4029 gnd.n2145 585
R12199 gnd.n3987 gnd.n3975 585
R12200 gnd.n3975 gnd.n2150 585
R12201 gnd.n3988 gnd.n3974 585
R12202 gnd.n3974 gnd.n2159 585
R12203 gnd.n3989 gnd.n3973 585
R12204 gnd.n3973 gnd.n2155 585
R12205 gnd.n2175 gnd.n2166 585
R12206 gnd.n4004 gnd.n2166 585
R12207 gnd.n3994 gnd.n3993 585
R12208 gnd.n3996 gnd.n3994 585
R12209 gnd.n2174 gnd.n2173 585
R12210 gnd.n3925 gnd.n2173 585
R12211 gnd.n3969 gnd.n3968 585
R12212 gnd.n3968 gnd.n3967 585
R12213 gnd.n2178 gnd.n2177 585
R12214 gnd.n3959 gnd.n2178 585
R12215 gnd.n3810 gnd.n3809 585
R12216 gnd.n3809 gnd.n2195 585
R12217 gnd.n3813 gnd.n3808 585
R12218 gnd.n3808 gnd.n2192 585
R12219 gnd.n3814 gnd.n3807 585
R12220 gnd.n3807 gnd.n2199 585
R12221 gnd.n3815 gnd.n3806 585
R12222 gnd.n3806 gnd.n2203 585
R12223 gnd.n3805 gnd.n3803 585
R12224 gnd.n3805 gnd.n2212 585
R12225 gnd.n3819 gnd.n3802 585
R12226 gnd.n3802 gnd.n2209 585
R12227 gnd.n3820 gnd.n3801 585
R12228 gnd.n3801 gnd.n2217 585
R12229 gnd.n3821 gnd.n2226 585
R12230 gnd.n3879 gnd.n2226 585
R12231 gnd.n3799 gnd.n2233 585
R12232 gnd.n3868 gnd.n2233 585
R12233 gnd.n3825 gnd.n3798 585
R12234 gnd.n3798 gnd.n2237 585
R12235 gnd.n3826 gnd.n3797 585
R12236 gnd.n3797 gnd.n2246 585
R12237 gnd.n3827 gnd.n3796 585
R12238 gnd.n3796 gnd.n2242 585
R12239 gnd.n2262 gnd.n2253 585
R12240 gnd.n3842 gnd.n2253 585
R12241 gnd.n3832 gnd.n3831 585
R12242 gnd.n3833 gnd.n3832 585
R12243 gnd.n2261 gnd.n2260 585
R12244 gnd.n3747 gnd.n2260 585
R12245 gnd.n3792 gnd.n3791 585
R12246 gnd.n3791 gnd.n3790 585
R12247 gnd.n2265 gnd.n2264 585
R12248 gnd.n3782 gnd.n2265 585
R12249 gnd.n3634 gnd.n3633 585
R12250 gnd.n3633 gnd.n2282 585
R12251 gnd.n3637 gnd.n3632 585
R12252 gnd.n3632 gnd.n2280 585
R12253 gnd.n3638 gnd.n3631 585
R12254 gnd.n3631 gnd.n2286 585
R12255 gnd.n3639 gnd.n3630 585
R12256 gnd.n3630 gnd.n2291 585
R12257 gnd.n3629 gnd.n3627 585
R12258 gnd.n3629 gnd.n2298 585
R12259 gnd.n3643 gnd.n3626 585
R12260 gnd.n3626 gnd.n3625 585
R12261 gnd.n3644 gnd.n3623 585
R12262 gnd.n3623 gnd.n2303 585
R12263 gnd.n3645 gnd.n2311 585
R12264 gnd.n3702 gnd.n2311 585
R12265 gnd.n3621 gnd.n2318 585
R12266 gnd.n3690 gnd.n2318 585
R12267 gnd.n3649 gnd.n3620 585
R12268 gnd.n3620 gnd.n2322 585
R12269 gnd.n3650 gnd.n3619 585
R12270 gnd.n3619 gnd.n2331 585
R12271 gnd.n3651 gnd.n3618 585
R12272 gnd.n3618 gnd.n2328 585
R12273 gnd.n2347 gnd.n2338 585
R12274 gnd.n3665 gnd.n2338 585
R12275 gnd.n3656 gnd.n3655 585
R12276 gnd.n3657 gnd.n3656 585
R12277 gnd.n2346 gnd.n2345 585
R12278 gnd.n2462 gnd.n2345 585
R12279 gnd.n3614 gnd.n3613 585
R12280 gnd.n3613 gnd.n3612 585
R12281 gnd.n2350 gnd.n2349 585
R12282 gnd.n3603 gnd.n2350 585
R12283 gnd.n2376 gnd.n2374 585
R12284 gnd.n2374 gnd.t245 585
R12285 gnd.n3581 gnd.n3580 585
R12286 gnd.n3582 gnd.n3581 585
R12287 gnd.n2375 gnd.n2373 585
R12288 gnd.n2373 gnd.n2370 585
R12289 gnd.n3575 gnd.n3574 585
R12290 gnd.n3574 gnd.n3573 585
R12291 gnd.n2379 gnd.n2378 585
R12292 gnd.n2421 gnd.n2379 585
R12293 gnd.n3402 gnd.n3401 585
R12294 gnd.n3401 gnd.n2387 585
R12295 gnd.n3400 gnd.n2683 585
R12296 gnd.n3400 gnd.n3399 585
R12297 gnd.n3406 gnd.n2682 585
R12298 gnd.n2684 gnd.n2682 585
R12299 gnd.n3407 gnd.n2681 585
R12300 gnd.n3387 gnd.n2681 585
R12301 gnd.n3408 gnd.n2680 585
R12302 gnd.n3385 gnd.n2680 585
R12303 gnd.n3381 gnd.n2678 585
R12304 gnd.n3383 gnd.n3381 585
R12305 gnd.n3412 gnd.n2677 585
R12306 gnd.n2690 gnd.n2677 585
R12307 gnd.n3413 gnd.n2676 585
R12308 gnd.n3371 gnd.n2676 585
R12309 gnd.n3414 gnd.n2675 585
R12310 gnd.n3369 gnd.n2675 585
R12311 gnd.n3365 gnd.n2673 585
R12312 gnd.n3367 gnd.n3365 585
R12313 gnd.n3418 gnd.n2672 585
R12314 gnd.n2696 gnd.n2672 585
R12315 gnd.n3419 gnd.n2671 585
R12316 gnd.n3355 gnd.n2671 585
R12317 gnd.n3420 gnd.n2670 585
R12318 gnd.n3353 gnd.n2670 585
R12319 gnd.n3349 gnd.n2668 585
R12320 gnd.n3351 gnd.n3349 585
R12321 gnd.n3424 gnd.n2667 585
R12322 gnd.n2702 gnd.n2667 585
R12323 gnd.n3425 gnd.n2666 585
R12324 gnd.n3339 gnd.n2666 585
R12325 gnd.n3426 gnd.n2665 585
R12326 gnd.n3337 gnd.n2665 585
R12327 gnd.n1799 gnd.n1798 585
R12328 gnd.n1798 gnd.n1467 585
R12329 gnd.n4460 gnd.n1797 585
R12330 gnd.n4461 gnd.n1795 585
R12331 gnd.n4462 gnd.n1794 585
R12332 gnd.n1792 gnd.n1787 585
R12333 gnd.n4466 gnd.n1786 585
R12334 gnd.n4467 gnd.n1784 585
R12335 gnd.n4468 gnd.n1783 585
R12336 gnd.n1781 gnd.n1779 585
R12337 gnd.n4472 gnd.n1778 585
R12338 gnd.n4473 gnd.n1776 585
R12339 gnd.n4474 gnd.n1775 585
R12340 gnd.n1773 gnd.n1650 585
R12341 gnd.n1772 gnd.n1771 585
R12342 gnd.n1756 gnd.n1652 585
R12343 gnd.n1758 gnd.n1757 585
R12344 gnd.n1754 gnd.n1659 585
R12345 gnd.n1753 gnd.n1752 585
R12346 gnd.n1737 gnd.n1661 585
R12347 gnd.n1739 gnd.n1738 585
R12348 gnd.n1735 gnd.n1668 585
R12349 gnd.n1734 gnd.n1733 585
R12350 gnd.n1718 gnd.n1670 585
R12351 gnd.n1720 gnd.n1719 585
R12352 gnd.n1716 gnd.n1677 585
R12353 gnd.n1715 gnd.n1714 585
R12354 gnd.n1699 gnd.n1679 585
R12355 gnd.n1701 gnd.n1700 585
R12356 gnd.n1697 gnd.n1455 585
R12357 gnd.n4300 gnd.n2039 468.476
R12358 gnd.n4303 gnd.n4302 468.476
R12359 gnd.n2479 gnd.n2478 468.476
R12360 gnd.n3561 gnd.n2424 468.476
R12361 gnd.n6696 gnd.n6695 457.279
R12362 gnd.n2450 gnd.t266 389.64
R12363 gnd.n2032 gnd.t247 389.64
R12364 gnd.n2447 gnd.t213 389.64
R12365 gnd.n4231 gnd.t272 389.64
R12366 gnd.n2656 gnd.t240 371.625
R12367 gnd.n7613 gnd.t269 371.625
R12368 gnd.n1645 gnd.t260 371.625
R12369 gnd.n2782 gnd.t285 371.625
R12370 gnd.n1948 gnd.t234 371.625
R12371 gnd.n1977 gnd.t220 371.625
R12372 gnd.n180 gnd.t291 371.625
R12373 gnd.n7706 gnd.t209 371.625
R12374 gnd.n1031 gnd.t193 371.625
R12375 gnd.n1053 gnd.t282 371.625
R12376 gnd.n2634 gnd.t288 371.625
R12377 gnd.n2545 gnd.t201 371.625
R12378 gnd.n3041 gnd.t227 371.625
R12379 gnd.n1789 gnd.t197 371.625
R12380 gnd.n5707 gnd.t278 323.425
R12381 gnd.n5161 gnd.t205 323.425
R12382 gnd.n6375 gnd.n6349 289.615
R12383 gnd.n6343 gnd.n6317 289.615
R12384 gnd.n6311 gnd.n6285 289.615
R12385 gnd.n6280 gnd.n6254 289.615
R12386 gnd.n6248 gnd.n6222 289.615
R12387 gnd.n6216 gnd.n6190 289.615
R12388 gnd.n6184 gnd.n6158 289.615
R12389 gnd.n6153 gnd.n6127 289.615
R12390 gnd.n5557 gnd.t230 279.217
R12391 gnd.n5187 gnd.t186 279.217
R12392 gnd.n2431 gnd.t219 260.649
R12393 gnd.n4223 gnd.t253 260.649
R12394 gnd.n3563 gnd.n3562 256.663
R12395 gnd.n3563 gnd.n2388 256.663
R12396 gnd.n3563 gnd.n2389 256.663
R12397 gnd.n3563 gnd.n2390 256.663
R12398 gnd.n3563 gnd.n2391 256.663
R12399 gnd.n3563 gnd.n2392 256.663
R12400 gnd.n3563 gnd.n2393 256.663
R12401 gnd.n3563 gnd.n2394 256.663
R12402 gnd.n3563 gnd.n2395 256.663
R12403 gnd.n3563 gnd.n2396 256.663
R12404 gnd.n3563 gnd.n2397 256.663
R12405 gnd.n3563 gnd.n2398 256.663
R12406 gnd.n3563 gnd.n2399 256.663
R12407 gnd.n3563 gnd.n2400 256.663
R12408 gnd.n3563 gnd.n2401 256.663
R12409 gnd.n3563 gnd.n2402 256.663
R12410 gnd.n3499 gnd.n3496 256.663
R12411 gnd.n3563 gnd.n2403 256.663
R12412 gnd.n3563 gnd.n2404 256.663
R12413 gnd.n3563 gnd.n2405 256.663
R12414 gnd.n3563 gnd.n2406 256.663
R12415 gnd.n3563 gnd.n2407 256.663
R12416 gnd.n3563 gnd.n2408 256.663
R12417 gnd.n3563 gnd.n2409 256.663
R12418 gnd.n3563 gnd.n2410 256.663
R12419 gnd.n3563 gnd.n2411 256.663
R12420 gnd.n3563 gnd.n2412 256.663
R12421 gnd.n3563 gnd.n2413 256.663
R12422 gnd.n3563 gnd.n2414 256.663
R12423 gnd.n3563 gnd.n2415 256.663
R12424 gnd.n3563 gnd.n2416 256.663
R12425 gnd.n3563 gnd.n2417 256.663
R12426 gnd.n3563 gnd.n2418 256.663
R12427 gnd.n3563 gnd.n2419 256.663
R12428 gnd.n4369 gnd.n1872 256.663
R12429 gnd.n4369 gnd.n1873 256.663
R12430 gnd.n4369 gnd.n1874 256.663
R12431 gnd.n4369 gnd.n1875 256.663
R12432 gnd.n4369 gnd.n1876 256.663
R12433 gnd.n4369 gnd.n1877 256.663
R12434 gnd.n4369 gnd.n1878 256.663
R12435 gnd.n4369 gnd.n1879 256.663
R12436 gnd.n4369 gnd.n1880 256.663
R12437 gnd.n4369 gnd.n1881 256.663
R12438 gnd.n4369 gnd.n1882 256.663
R12439 gnd.n4369 gnd.n1883 256.663
R12440 gnd.n4369 gnd.n1884 256.663
R12441 gnd.n4369 gnd.n1885 256.663
R12442 gnd.n4369 gnd.n1886 256.663
R12443 gnd.n4369 gnd.n1887 256.663
R12444 gnd.n2031 gnd.n1888 256.663
R12445 gnd.n4369 gnd.n1869 256.663
R12446 gnd.n4369 gnd.n1868 256.663
R12447 gnd.n4369 gnd.n1867 256.663
R12448 gnd.n4369 gnd.n1866 256.663
R12449 gnd.n4369 gnd.n1865 256.663
R12450 gnd.n4369 gnd.n1864 256.663
R12451 gnd.n4369 gnd.n1863 256.663
R12452 gnd.n4369 gnd.n1862 256.663
R12453 gnd.n4369 gnd.n1861 256.663
R12454 gnd.n4369 gnd.n1860 256.663
R12455 gnd.n4369 gnd.n1859 256.663
R12456 gnd.n4369 gnd.n1858 256.663
R12457 gnd.n4369 gnd.n1857 256.663
R12458 gnd.n4369 gnd.n1856 256.663
R12459 gnd.n4369 gnd.n1855 256.663
R12460 gnd.n4369 gnd.n1854 256.663
R12461 gnd.n4369 gnd.n1853 256.663
R12462 gnd.n5138 gnd.n999 242.672
R12463 gnd.n5138 gnd.n1000 242.672
R12464 gnd.n5138 gnd.n1001 242.672
R12465 gnd.n5138 gnd.n1002 242.672
R12466 gnd.n5138 gnd.n1003 242.672
R12467 gnd.n5138 gnd.n1004 242.672
R12468 gnd.n5138 gnd.n1005 242.672
R12469 gnd.n5138 gnd.n1006 242.672
R12470 gnd.n5138 gnd.n1007 242.672
R12471 gnd.n2791 gnd.n2606 242.672
R12472 gnd.n2780 gnd.n2606 242.672
R12473 gnd.n2777 gnd.n2606 242.672
R12474 gnd.n2768 gnd.n2606 242.672
R12475 gnd.n2757 gnd.n2606 242.672
R12476 gnd.n2754 gnd.n2606 242.672
R12477 gnd.n2745 gnd.n2606 242.672
R12478 gnd.n2735 gnd.n2606 242.672
R12479 gnd.n2732 gnd.n2606 242.672
R12480 gnd.n1686 gnd.n1468 242.672
R12481 gnd.n1706 gnd.n1468 242.672
R12482 gnd.n1708 gnd.n1468 242.672
R12483 gnd.n1725 gnd.n1468 242.672
R12484 gnd.n1727 gnd.n1468 242.672
R12485 gnd.n1744 gnd.n1468 242.672
R12486 gnd.n1746 gnd.n1468 242.672
R12487 gnd.n1763 gnd.n1468 242.672
R12488 gnd.n1765 gnd.n1468 242.672
R12489 gnd.n7615 gnd.n117 242.672
R12490 gnd.n7611 gnd.n117 242.672
R12491 gnd.n7606 gnd.n117 242.672
R12492 gnd.n7603 gnd.n117 242.672
R12493 gnd.n7598 gnd.n117 242.672
R12494 gnd.n7595 gnd.n117 242.672
R12495 gnd.n7590 gnd.n117 242.672
R12496 gnd.n7587 gnd.n117 242.672
R12497 gnd.n7582 gnd.n117 242.672
R12498 gnd.n5612 gnd.n5521 242.672
R12499 gnd.n5525 gnd.n5521 242.672
R12500 gnd.n5605 gnd.n5521 242.672
R12501 gnd.n5599 gnd.n5521 242.672
R12502 gnd.n5597 gnd.n5521 242.672
R12503 gnd.n5591 gnd.n5521 242.672
R12504 gnd.n5589 gnd.n5521 242.672
R12505 gnd.n5583 gnd.n5521 242.672
R12506 gnd.n5581 gnd.n5521 242.672
R12507 gnd.n5575 gnd.n5521 242.672
R12508 gnd.n5573 gnd.n5521 242.672
R12509 gnd.n5566 gnd.n5521 242.672
R12510 gnd.n5564 gnd.n5521 242.672
R12511 gnd.n6490 gnd.n980 242.672
R12512 gnd.n6490 gnd.n979 242.672
R12513 gnd.n6490 gnd.n978 242.672
R12514 gnd.n6490 gnd.n977 242.672
R12515 gnd.n6490 gnd.n976 242.672
R12516 gnd.n6490 gnd.n975 242.672
R12517 gnd.n6490 gnd.n974 242.672
R12518 gnd.n6490 gnd.n973 242.672
R12519 gnd.n6490 gnd.n972 242.672
R12520 gnd.n6490 gnd.n971 242.672
R12521 gnd.n6490 gnd.n970 242.672
R12522 gnd.n6490 gnd.n969 242.672
R12523 gnd.n6490 gnd.n968 242.672
R12524 gnd.n5741 gnd.n5740 242.672
R12525 gnd.n5741 gnd.n5682 242.672
R12526 gnd.n5741 gnd.n5683 242.672
R12527 gnd.n5741 gnd.n5684 242.672
R12528 gnd.n5741 gnd.n5685 242.672
R12529 gnd.n5741 gnd.n5686 242.672
R12530 gnd.n5741 gnd.n5687 242.672
R12531 gnd.n5741 gnd.n5688 242.672
R12532 gnd.n6490 gnd.n5139 242.672
R12533 gnd.n6490 gnd.n5140 242.672
R12534 gnd.n6490 gnd.n5141 242.672
R12535 gnd.n6490 gnd.n5142 242.672
R12536 gnd.n6490 gnd.n5143 242.672
R12537 gnd.n6490 gnd.n5144 242.672
R12538 gnd.n6490 gnd.n5145 242.672
R12539 gnd.n6490 gnd.n6489 242.672
R12540 gnd.n5138 gnd.n5137 242.672
R12541 gnd.n5138 gnd.n981 242.672
R12542 gnd.n5138 gnd.n982 242.672
R12543 gnd.n5138 gnd.n983 242.672
R12544 gnd.n5138 gnd.n984 242.672
R12545 gnd.n5138 gnd.n985 242.672
R12546 gnd.n5138 gnd.n986 242.672
R12547 gnd.n5138 gnd.n987 242.672
R12548 gnd.n5138 gnd.n988 242.672
R12549 gnd.n5138 gnd.n989 242.672
R12550 gnd.n5138 gnd.n990 242.672
R12551 gnd.n5138 gnd.n991 242.672
R12552 gnd.n5138 gnd.n992 242.672
R12553 gnd.n5138 gnd.n993 242.672
R12554 gnd.n5138 gnd.n994 242.672
R12555 gnd.n5138 gnd.n995 242.672
R12556 gnd.n5138 gnd.n996 242.672
R12557 gnd.n5138 gnd.n997 242.672
R12558 gnd.n5138 gnd.n998 242.672
R12559 gnd.n3458 gnd.n2606 242.672
R12560 gnd.n2637 gnd.n2606 242.672
R12561 gnd.n3465 gnd.n2606 242.672
R12562 gnd.n2628 gnd.n2606 242.672
R12563 gnd.n3472 gnd.n2606 242.672
R12564 gnd.n2621 gnd.n2606 242.672
R12565 gnd.n3479 gnd.n2606 242.672
R12566 gnd.n2614 gnd.n2606 242.672
R12567 gnd.n3486 gnd.n2606 242.672
R12568 gnd.n3489 gnd.n2606 242.672
R12569 gnd.n2606 gnd.n2552 242.672
R12570 gnd.n3495 gnd.n2547 242.672
R12571 gnd.n2606 gnd.n2553 242.672
R12572 gnd.n2606 gnd.n2554 242.672
R12573 gnd.n2606 gnd.n2555 242.672
R12574 gnd.n2606 gnd.n2556 242.672
R12575 gnd.n2606 gnd.n2557 242.672
R12576 gnd.n2606 gnd.n2558 242.672
R12577 gnd.n2606 gnd.n2559 242.672
R12578 gnd.n2606 gnd.n2605 242.672
R12579 gnd.n1910 gnd.n1468 242.672
R12580 gnd.n1918 gnd.n1468 242.672
R12581 gnd.n1920 gnd.n1468 242.672
R12582 gnd.n1928 gnd.n1468 242.672
R12583 gnd.n1930 gnd.n1468 242.672
R12584 gnd.n1939 gnd.n1468 242.672
R12585 gnd.n1942 gnd.n1468 242.672
R12586 gnd.n1893 gnd.n1468 242.672
R12587 gnd.n2030 gnd.n1890 242.672
R12588 gnd.n2027 gnd.n1468 242.672
R12589 gnd.n2025 gnd.n1468 242.672
R12590 gnd.n2019 gnd.n1468 242.672
R12591 gnd.n2017 gnd.n1468 242.672
R12592 gnd.n2011 gnd.n1468 242.672
R12593 gnd.n2009 gnd.n1468 242.672
R12594 gnd.n2003 gnd.n1468 242.672
R12595 gnd.n2001 gnd.n1468 242.672
R12596 gnd.n1995 gnd.n1468 242.672
R12597 gnd.n1993 gnd.n1468 242.672
R12598 gnd.n1985 gnd.n1468 242.672
R12599 gnd.n177 gnd.n117 242.672
R12600 gnd.n7674 gnd.n117 242.672
R12601 gnd.n173 gnd.n117 242.672
R12602 gnd.n7681 gnd.n117 242.672
R12603 gnd.n166 gnd.n117 242.672
R12604 gnd.n7688 gnd.n117 242.672
R12605 gnd.n159 gnd.n117 242.672
R12606 gnd.n7695 gnd.n117 242.672
R12607 gnd.n152 gnd.n117 242.672
R12608 gnd.n7702 gnd.n117 242.672
R12609 gnd.n145 gnd.n117 242.672
R12610 gnd.n7712 gnd.n117 242.672
R12611 gnd.n138 gnd.n117 242.672
R12612 gnd.n7719 gnd.n117 242.672
R12613 gnd.n131 gnd.n117 242.672
R12614 gnd.n7726 gnd.n117 242.672
R12615 gnd.n124 gnd.n117 242.672
R12616 gnd.n7733 gnd.n117 242.672
R12617 gnd.n117 gnd.n116 242.672
R12618 gnd.n2840 gnd.n2839 242.672
R12619 gnd.n2840 gnd.n2708 242.672
R12620 gnd.n2840 gnd.n2709 242.672
R12621 gnd.n2840 gnd.n2710 242.672
R12622 gnd.n2840 gnd.n2711 242.672
R12623 gnd.n2840 gnd.n2712 242.672
R12624 gnd.n2840 gnd.n2713 242.672
R12625 gnd.n2840 gnd.n2714 242.672
R12626 gnd.n2840 gnd.n2715 242.672
R12627 gnd.n2840 gnd.n2716 242.672
R12628 gnd.n2840 gnd.n2718 242.672
R12629 gnd.n2840 gnd.n2719 242.672
R12630 gnd.n2840 gnd.n2720 242.672
R12631 gnd.n2840 gnd.n2722 242.672
R12632 gnd.n1796 gnd.n1467 242.672
R12633 gnd.n1793 gnd.n1467 242.672
R12634 gnd.n1785 gnd.n1467 242.672
R12635 gnd.n1782 gnd.n1467 242.672
R12636 gnd.n1777 gnd.n1467 242.672
R12637 gnd.n1774 gnd.n1467 242.672
R12638 gnd.n1651 gnd.n1467 242.672
R12639 gnd.n1755 gnd.n1467 242.672
R12640 gnd.n1660 gnd.n1467 242.672
R12641 gnd.n1736 gnd.n1467 242.672
R12642 gnd.n1669 gnd.n1467 242.672
R12643 gnd.n1717 gnd.n1467 242.672
R12644 gnd.n1678 gnd.n1467 242.672
R12645 gnd.n1698 gnd.n1467 242.672
R12646 gnd.n113 gnd.n109 240.244
R12647 gnd.n7735 gnd.n7734 240.244
R12648 gnd.n7732 gnd.n118 240.244
R12649 gnd.n7728 gnd.n7727 240.244
R12650 gnd.n7725 gnd.n125 240.244
R12651 gnd.n7721 gnd.n7720 240.244
R12652 gnd.n7718 gnd.n132 240.244
R12653 gnd.n7714 gnd.n7713 240.244
R12654 gnd.n7711 gnd.n139 240.244
R12655 gnd.n7704 gnd.n7703 240.244
R12656 gnd.n7701 gnd.n146 240.244
R12657 gnd.n7697 gnd.n7696 240.244
R12658 gnd.n7694 gnd.n153 240.244
R12659 gnd.n7690 gnd.n7689 240.244
R12660 gnd.n7687 gnd.n160 240.244
R12661 gnd.n7683 gnd.n7682 240.244
R12662 gnd.n7680 gnd.n167 240.244
R12663 gnd.n7676 gnd.n7675 240.244
R12664 gnd.n7673 gnd.n174 240.244
R12665 gnd.n1984 gnd.n1478 240.244
R12666 gnd.n4488 gnd.n1478 240.244
R12667 gnd.n4488 gnd.n1491 240.244
R12668 gnd.n1636 gnd.n1491 240.244
R12669 gnd.n4519 gnd.n1636 240.244
R12670 gnd.n4519 gnd.n1637 240.244
R12671 gnd.n1637 gnd.n1617 240.244
R12672 gnd.n1617 gnd.n1606 240.244
R12673 gnd.n4513 gnd.n1606 240.244
R12674 gnd.n4513 gnd.n1597 240.244
R12675 gnd.n4510 gnd.n1597 240.244
R12676 gnd.n4510 gnd.n1590 240.244
R12677 gnd.n1590 gnd.n1579 240.244
R12678 gnd.n4506 gnd.n1579 240.244
R12679 gnd.n4506 gnd.n1568 240.244
R12680 gnd.n1568 gnd.n1560 240.244
R12681 gnd.n4613 gnd.n1560 240.244
R12682 gnd.n4613 gnd.n1526 240.244
R12683 gnd.n4616 gnd.n1526 240.244
R12684 gnd.n4616 gnd.n1518 240.244
R12685 gnd.n4624 gnd.n1518 240.244
R12686 gnd.n4624 gnd.n278 240.244
R12687 gnd.n4638 gnd.n278 240.244
R12688 gnd.n4639 gnd.n4638 240.244
R12689 gnd.n4639 gnd.n1542 240.244
R12690 gnd.n4645 gnd.n1542 240.244
R12691 gnd.n4645 gnd.n298 240.244
R12692 gnd.n7479 gnd.n298 240.244
R12693 gnd.n7479 gnd.n295 240.244
R12694 gnd.n7475 gnd.n295 240.244
R12695 gnd.n7475 gnd.n263 240.244
R12696 gnd.n7407 gnd.n263 240.244
R12697 gnd.n7407 gnd.n256 240.244
R12698 gnd.n7414 gnd.n256 240.244
R12699 gnd.n7414 gnd.n248 240.244
R12700 gnd.n7418 gnd.n248 240.244
R12701 gnd.n7418 gnd.n240 240.244
R12702 gnd.n7455 gnd.n240 240.244
R12703 gnd.n7455 gnd.n232 240.244
R12704 gnd.n7451 gnd.n232 240.244
R12705 gnd.n7451 gnd.n226 240.244
R12706 gnd.n7447 gnd.n226 240.244
R12707 gnd.n7447 gnd.n219 240.244
R12708 gnd.n7444 gnd.n219 240.244
R12709 gnd.n7444 gnd.n209 240.244
R12710 gnd.n7441 gnd.n209 240.244
R12711 gnd.n7441 gnd.n202 240.244
R12712 gnd.n7438 gnd.n202 240.244
R12713 gnd.n7438 gnd.n194 240.244
R12714 gnd.n194 gnd.n184 240.244
R12715 gnd.n7664 gnd.n184 240.244
R12716 gnd.n7665 gnd.n7664 240.244
R12717 gnd.n7665 gnd.n105 240.244
R12718 gnd.n1911 gnd.n1904 240.244
R12719 gnd.n1917 gnd.n1904 240.244
R12720 gnd.n1921 gnd.n1919 240.244
R12721 gnd.n1927 gnd.n1900 240.244
R12722 gnd.n1931 gnd.n1929 240.244
R12723 gnd.n1938 gnd.n1896 240.244
R12724 gnd.n1941 gnd.n1940 240.244
R12725 gnd.n1943 gnd.n1894 240.244
R12726 gnd.n2028 gnd.n2026 240.244
R12727 gnd.n2024 gnd.n1952 240.244
R12728 gnd.n2020 gnd.n2018 240.244
R12729 gnd.n2016 gnd.n1958 240.244
R12730 gnd.n2012 gnd.n2010 240.244
R12731 gnd.n2008 gnd.n1964 240.244
R12732 gnd.n2004 gnd.n2002 240.244
R12733 gnd.n2000 gnd.n1970 240.244
R12734 gnd.n1996 gnd.n1994 240.244
R12735 gnd.n1992 gnd.n1976 240.244
R12736 gnd.n4723 gnd.n1482 240.244
R12737 gnd.n4723 gnd.n1483 240.244
R12738 gnd.n4719 gnd.n1483 240.244
R12739 gnd.n4719 gnd.n1489 240.244
R12740 gnd.n4527 gnd.n1489 240.244
R12741 gnd.n4527 gnd.n4521 240.244
R12742 gnd.n4521 gnd.n1604 240.244
R12743 gnd.n4551 gnd.n1604 240.244
R12744 gnd.n4551 gnd.n1599 240.244
R12745 gnd.n4559 gnd.n1599 240.244
R12746 gnd.n4559 gnd.n1600 240.244
R12747 gnd.n1600 gnd.n1577 240.244
R12748 gnd.n4590 gnd.n1577 240.244
R12749 gnd.n4590 gnd.n1570 240.244
R12750 gnd.n4598 gnd.n1570 240.244
R12751 gnd.n4598 gnd.n1573 240.244
R12752 gnd.n1573 gnd.n1525 240.244
R12753 gnd.n4680 gnd.n1525 240.244
R12754 gnd.n4680 gnd.n1521 240.244
R12755 gnd.n4686 gnd.n1521 240.244
R12756 gnd.n4686 gnd.n275 240.244
R12757 gnd.n7502 gnd.n275 240.244
R12758 gnd.n7502 gnd.n276 240.244
R12759 gnd.n1545 gnd.n276 240.244
R12760 gnd.n4663 gnd.n1545 240.244
R12761 gnd.n4663 gnd.n4661 240.244
R12762 gnd.n4661 gnd.n297 240.244
R12763 gnd.n7481 gnd.n297 240.244
R12764 gnd.n7484 gnd.n7481 240.244
R12765 gnd.n7484 gnd.n265 240.244
R12766 gnd.n7507 gnd.n265 240.244
R12767 gnd.n7507 gnd.n254 240.244
R12768 gnd.n7517 gnd.n254 240.244
R12769 gnd.n7517 gnd.n250 240.244
R12770 gnd.n7523 gnd.n250 240.244
R12771 gnd.n7523 gnd.n238 240.244
R12772 gnd.n7533 gnd.n238 240.244
R12773 gnd.n7533 gnd.n234 240.244
R12774 gnd.n7539 gnd.n234 240.244
R12775 gnd.n7539 gnd.n224 240.244
R12776 gnd.n7549 gnd.n224 240.244
R12777 gnd.n7549 gnd.n220 240.244
R12778 gnd.n7555 gnd.n220 240.244
R12779 gnd.n7555 gnd.n207 240.244
R12780 gnd.n7565 gnd.n207 240.244
R12781 gnd.n7565 gnd.n203 240.244
R12782 gnd.n7571 gnd.n203 240.244
R12783 gnd.n7571 gnd.n192 240.244
R12784 gnd.n7656 gnd.n192 240.244
R12785 gnd.n7656 gnd.n188 240.244
R12786 gnd.n7662 gnd.n188 240.244
R12787 gnd.n7662 gnd.n108 240.244
R12788 gnd.n7742 gnd.n108 240.244
R12789 gnd.n2560 gnd.n1319 240.244
R12790 gnd.n2604 gnd.n2561 240.244
R12791 gnd.n2600 gnd.n2599 240.244
R12792 gnd.n2596 gnd.n2595 240.244
R12793 gnd.n2592 gnd.n2591 240.244
R12794 gnd.n2588 gnd.n2587 240.244
R12795 gnd.n2584 gnd.n2583 240.244
R12796 gnd.n2580 gnd.n2579 240.244
R12797 gnd.n3490 gnd.n2551 240.244
R12798 gnd.n3488 gnd.n3487 240.244
R12799 gnd.n3485 gnd.n2608 240.244
R12800 gnd.n3481 gnd.n3480 240.244
R12801 gnd.n3478 gnd.n2615 240.244
R12802 gnd.n3474 gnd.n3473 240.244
R12803 gnd.n3471 gnd.n2622 240.244
R12804 gnd.n3467 gnd.n3466 240.244
R12805 gnd.n3464 gnd.n2629 240.244
R12806 gnd.n3460 gnd.n3459 240.244
R12807 gnd.n5059 gnd.n1057 240.244
R12808 gnd.n1061 gnd.n1057 240.244
R12809 gnd.n5052 gnd.n1061 240.244
R12810 gnd.n5052 gnd.n1062 240.244
R12811 gnd.n1075 gnd.n1062 240.244
R12812 gnd.n3126 gnd.n1075 240.244
R12813 gnd.n3126 gnd.n1086 240.244
R12814 gnd.n3131 gnd.n1086 240.244
R12815 gnd.n3131 gnd.n1096 240.244
R12816 gnd.n3134 gnd.n1096 240.244
R12817 gnd.n3134 gnd.n1106 240.244
R12818 gnd.n3140 gnd.n1106 240.244
R12819 gnd.n3140 gnd.n1117 240.244
R12820 gnd.n3150 gnd.n1117 240.244
R12821 gnd.n3150 gnd.n1128 240.244
R12822 gnd.n3156 gnd.n1128 240.244
R12823 gnd.n3156 gnd.n1139 240.244
R12824 gnd.n3166 gnd.n1139 240.244
R12825 gnd.n3166 gnd.n1149 240.244
R12826 gnd.n3172 gnd.n1149 240.244
R12827 gnd.n3172 gnd.n1159 240.244
R12828 gnd.n3182 gnd.n1159 240.244
R12829 gnd.n3182 gnd.n1170 240.244
R12830 gnd.n3188 gnd.n1170 240.244
R12831 gnd.n3188 gnd.n1179 240.244
R12832 gnd.n3199 gnd.n1179 240.244
R12833 gnd.n3199 gnd.n1189 240.244
R12834 gnd.n3206 gnd.n1189 240.244
R12835 gnd.n3206 gnd.n1196 240.244
R12836 gnd.n3216 gnd.n1196 240.244
R12837 gnd.n3216 gnd.n1207 240.244
R12838 gnd.n3222 gnd.n1207 240.244
R12839 gnd.n3222 gnd.n1217 240.244
R12840 gnd.n3232 gnd.n1217 240.244
R12841 gnd.n3232 gnd.n1227 240.244
R12842 gnd.n3238 gnd.n1227 240.244
R12843 gnd.n3238 gnd.n1237 240.244
R12844 gnd.n3248 gnd.n1237 240.244
R12845 gnd.n3248 gnd.n1248 240.244
R12846 gnd.n3255 gnd.n1248 240.244
R12847 gnd.n3255 gnd.n1259 240.244
R12848 gnd.n3265 gnd.n1259 240.244
R12849 gnd.n3265 gnd.n1269 240.244
R12850 gnd.n2858 gnd.n1269 240.244
R12851 gnd.n2858 gnd.n1279 240.244
R12852 gnd.n3273 gnd.n1279 240.244
R12853 gnd.n3273 gnd.n1290 240.244
R12854 gnd.n3277 gnd.n1290 240.244
R12855 gnd.n3277 gnd.n1301 240.244
R12856 gnd.n3284 gnd.n1301 240.244
R12857 gnd.n3284 gnd.n1312 240.244
R12858 gnd.n3451 gnd.n1312 240.244
R12859 gnd.n3451 gnd.n1321 240.244
R12860 gnd.n1011 gnd.n1010 240.244
R12861 gnd.n5131 gnd.n1010 240.244
R12862 gnd.n5129 gnd.n5128 240.244
R12863 gnd.n5125 gnd.n5124 240.244
R12864 gnd.n5121 gnd.n5120 240.244
R12865 gnd.n5117 gnd.n5116 240.244
R12866 gnd.n5113 gnd.n5112 240.244
R12867 gnd.n5109 gnd.n5108 240.244
R12868 gnd.n5105 gnd.n5104 240.244
R12869 gnd.n5100 gnd.n5099 240.244
R12870 gnd.n5096 gnd.n5095 240.244
R12871 gnd.n5092 gnd.n5091 240.244
R12872 gnd.n5088 gnd.n5087 240.244
R12873 gnd.n5084 gnd.n5083 240.244
R12874 gnd.n5080 gnd.n5079 240.244
R12875 gnd.n5076 gnd.n5075 240.244
R12876 gnd.n5072 gnd.n5071 240.244
R12877 gnd.n5068 gnd.n5067 240.244
R12878 gnd.n1052 gnd.n1051 240.244
R12879 gnd.n3099 gnd.n1012 240.244
R12880 gnd.n3099 gnd.n1067 240.244
R12881 gnd.n5050 gnd.n1067 240.244
R12882 gnd.n5050 gnd.n1068 240.244
R12883 gnd.n5046 gnd.n1068 240.244
R12884 gnd.n5046 gnd.n1074 240.244
R12885 gnd.n5038 gnd.n1074 240.244
R12886 gnd.n5038 gnd.n1089 240.244
R12887 gnd.n5034 gnd.n1089 240.244
R12888 gnd.n5034 gnd.n1095 240.244
R12889 gnd.n5026 gnd.n1095 240.244
R12890 gnd.n5026 gnd.n1109 240.244
R12891 gnd.n5022 gnd.n1109 240.244
R12892 gnd.n5022 gnd.n1115 240.244
R12893 gnd.n5014 gnd.n1115 240.244
R12894 gnd.n5014 gnd.n1131 240.244
R12895 gnd.n5010 gnd.n1131 240.244
R12896 gnd.n5010 gnd.n1137 240.244
R12897 gnd.n5002 gnd.n1137 240.244
R12898 gnd.n5002 gnd.n1151 240.244
R12899 gnd.n4998 gnd.n1151 240.244
R12900 gnd.n4998 gnd.n1157 240.244
R12901 gnd.n4990 gnd.n1157 240.244
R12902 gnd.n4990 gnd.n1173 240.244
R12903 gnd.n4986 gnd.n1173 240.244
R12904 gnd.n4986 gnd.n1177 240.244
R12905 gnd.n4978 gnd.n1177 240.244
R12906 gnd.n4978 gnd.n1191 240.244
R12907 gnd.n4973 gnd.n1191 240.244
R12908 gnd.n4973 gnd.n1194 240.244
R12909 gnd.n4965 gnd.n1194 240.244
R12910 gnd.n4965 gnd.n1210 240.244
R12911 gnd.n4961 gnd.n1210 240.244
R12912 gnd.n4961 gnd.n1215 240.244
R12913 gnd.n4953 gnd.n1215 240.244
R12914 gnd.n4953 gnd.n1229 240.244
R12915 gnd.n4949 gnd.n1229 240.244
R12916 gnd.n4949 gnd.n1235 240.244
R12917 gnd.n4941 gnd.n1235 240.244
R12918 gnd.n4941 gnd.n1251 240.244
R12919 gnd.n4937 gnd.n1251 240.244
R12920 gnd.n4937 gnd.n1257 240.244
R12921 gnd.n4929 gnd.n1257 240.244
R12922 gnd.n4929 gnd.n1271 240.244
R12923 gnd.n4925 gnd.n1271 240.244
R12924 gnd.n4925 gnd.n1277 240.244
R12925 gnd.n4917 gnd.n1277 240.244
R12926 gnd.n4917 gnd.n1293 240.244
R12927 gnd.n4913 gnd.n1293 240.244
R12928 gnd.n4913 gnd.n1299 240.244
R12929 gnd.n4905 gnd.n1299 240.244
R12930 gnd.n4905 gnd.n1314 240.244
R12931 gnd.n4901 gnd.n1314 240.244
R12932 gnd.n6491 gnd.n965 240.244
R12933 gnd.n6488 gnd.n5146 240.244
R12934 gnd.n6484 gnd.n6483 240.244
R12935 gnd.n6480 gnd.n6479 240.244
R12936 gnd.n6476 gnd.n6475 240.244
R12937 gnd.n6472 gnd.n6471 240.244
R12938 gnd.n6468 gnd.n6467 240.244
R12939 gnd.n6464 gnd.n6463 240.244
R12940 gnd.n5753 gnd.n5473 240.244
R12941 gnd.n5473 gnd.n5464 240.244
R12942 gnd.n5771 gnd.n5464 240.244
R12943 gnd.n5772 gnd.n5771 240.244
R12944 gnd.n5772 gnd.n5452 240.244
R12945 gnd.n5452 gnd.n5441 240.244
R12946 gnd.n5803 gnd.n5441 240.244
R12947 gnd.n5804 gnd.n5803 240.244
R12948 gnd.n5805 gnd.n5804 240.244
R12949 gnd.n5805 gnd.n5426 240.244
R12950 gnd.n5807 gnd.n5426 240.244
R12951 gnd.n5807 gnd.n5411 240.244
R12952 gnd.n5848 gnd.n5411 240.244
R12953 gnd.n5849 gnd.n5848 240.244
R12954 gnd.n5852 gnd.n5849 240.244
R12955 gnd.n5852 gnd.n5393 240.244
R12956 gnd.n5884 gnd.n5393 240.244
R12957 gnd.n5884 gnd.n5379 240.244
R12958 gnd.n5906 gnd.n5379 240.244
R12959 gnd.n5907 gnd.n5906 240.244
R12960 gnd.n5907 gnd.n5366 240.244
R12961 gnd.n5366 gnd.n5355 240.244
R12962 gnd.n5938 gnd.n5355 240.244
R12963 gnd.n5939 gnd.n5938 240.244
R12964 gnd.n5940 gnd.n5939 240.244
R12965 gnd.n5940 gnd.n5292 240.244
R12966 gnd.n5292 gnd.n5291 240.244
R12967 gnd.n5291 gnd.n5276 240.244
R12968 gnd.n5991 gnd.n5276 240.244
R12969 gnd.n5992 gnd.n5991 240.244
R12970 gnd.n5992 gnd.n5263 240.244
R12971 gnd.n5263 gnd.n5252 240.244
R12972 gnd.n6025 gnd.n5252 240.244
R12973 gnd.n6026 gnd.n6025 240.244
R12974 gnd.n6028 gnd.n6026 240.244
R12975 gnd.n6028 gnd.n6027 240.244
R12976 gnd.n6027 gnd.n5231 240.244
R12977 gnd.n6063 gnd.n5231 240.244
R12978 gnd.n6063 gnd.n5223 240.244
R12979 gnd.n5223 gnd.n5216 240.244
R12980 gnd.n6088 gnd.n5216 240.244
R12981 gnd.n6088 gnd.n908 240.244
R12982 gnd.n6101 gnd.n908 240.244
R12983 gnd.n6101 gnd.n918 240.244
R12984 gnd.n5204 gnd.n918 240.244
R12985 gnd.n6121 gnd.n5204 240.244
R12986 gnd.n6121 gnd.n930 240.244
R12987 gnd.n5199 gnd.n930 240.244
R12988 gnd.n5199 gnd.n943 240.244
R12989 gnd.n5197 gnd.n943 240.244
R12990 gnd.n6396 gnd.n5197 240.244
R12991 gnd.n6396 gnd.n955 240.244
R12992 gnd.n6392 gnd.n955 240.244
R12993 gnd.n5690 gnd.n5689 240.244
R12994 gnd.n5734 gnd.n5689 240.244
R12995 gnd.n5732 gnd.n5731 240.244
R12996 gnd.n5728 gnd.n5727 240.244
R12997 gnd.n5724 gnd.n5723 240.244
R12998 gnd.n5720 gnd.n5719 240.244
R12999 gnd.n5716 gnd.n5715 240.244
R13000 gnd.n5712 gnd.n5711 240.244
R13001 gnd.n5763 gnd.n5471 240.244
R13002 gnd.n5763 gnd.n5467 240.244
R13003 gnd.n5769 gnd.n5467 240.244
R13004 gnd.n5769 gnd.n5450 240.244
R13005 gnd.n5793 gnd.n5450 240.244
R13006 gnd.n5793 gnd.n5445 240.244
R13007 gnd.n5801 gnd.n5445 240.244
R13008 gnd.n5801 gnd.n5446 240.244
R13009 gnd.n5446 gnd.n5424 240.244
R13010 gnd.n5827 gnd.n5424 240.244
R13011 gnd.n5827 gnd.n5419 240.244
R13012 gnd.n5838 gnd.n5419 240.244
R13013 gnd.n5838 gnd.n5420 240.244
R13014 gnd.n5834 gnd.n5420 240.244
R13015 gnd.n5834 gnd.n5391 240.244
R13016 gnd.n5888 gnd.n5391 240.244
R13017 gnd.n5888 gnd.n5386 240.244
R13018 gnd.n5896 gnd.n5386 240.244
R13019 gnd.n5896 gnd.n5387 240.244
R13020 gnd.n5387 gnd.n5364 240.244
R13021 gnd.n5928 gnd.n5364 240.244
R13022 gnd.n5928 gnd.n5359 240.244
R13023 gnd.n5936 gnd.n5359 240.244
R13024 gnd.n5936 gnd.n5360 240.244
R13025 gnd.n5360 gnd.n5289 240.244
R13026 gnd.n5973 gnd.n5289 240.244
R13027 gnd.n5973 gnd.n5284 240.244
R13028 gnd.n5981 gnd.n5284 240.244
R13029 gnd.n5981 gnd.n5285 240.244
R13030 gnd.n5285 gnd.n5261 240.244
R13031 gnd.n6012 gnd.n5261 240.244
R13032 gnd.n6012 gnd.n5256 240.244
R13033 gnd.n6023 gnd.n5256 240.244
R13034 gnd.n6023 gnd.n5257 240.244
R13035 gnd.n6019 gnd.n5257 240.244
R13036 gnd.n6019 gnd.n5230 240.244
R13037 gnd.n6067 gnd.n5230 240.244
R13038 gnd.n6067 gnd.n5225 240.244
R13039 gnd.n6076 gnd.n5225 240.244
R13040 gnd.n6076 gnd.n5226 240.244
R13041 gnd.n5226 gnd.n910 240.244
R13042 gnd.n6525 gnd.n910 240.244
R13043 gnd.n6525 gnd.n911 240.244
R13044 gnd.n6521 gnd.n911 240.244
R13045 gnd.n6521 gnd.n917 240.244
R13046 gnd.n932 gnd.n917 240.244
R13047 gnd.n6511 gnd.n932 240.244
R13048 gnd.n6511 gnd.n933 240.244
R13049 gnd.n6507 gnd.n933 240.244
R13050 gnd.n6507 gnd.n941 240.244
R13051 gnd.n957 gnd.n941 240.244
R13052 gnd.n6497 gnd.n957 240.244
R13053 gnd.n6497 gnd.n958 240.244
R13054 gnd.n5165 gnd.n967 240.244
R13055 gnd.n6454 gnd.n6453 240.244
R13056 gnd.n6450 gnd.n6449 240.244
R13057 gnd.n6446 gnd.n6445 240.244
R13058 gnd.n6442 gnd.n6441 240.244
R13059 gnd.n6438 gnd.n6437 240.244
R13060 gnd.n6434 gnd.n6433 240.244
R13061 gnd.n6430 gnd.n6429 240.244
R13062 gnd.n6426 gnd.n6425 240.244
R13063 gnd.n6422 gnd.n6421 240.244
R13064 gnd.n6418 gnd.n6417 240.244
R13065 gnd.n6414 gnd.n6413 240.244
R13066 gnd.n6410 gnd.n6409 240.244
R13067 gnd.n5621 gnd.n5517 240.244
R13068 gnd.n5627 gnd.n5517 240.244
R13069 gnd.n5627 gnd.n5509 240.244
R13070 gnd.n5637 gnd.n5509 240.244
R13071 gnd.n5637 gnd.n5505 240.244
R13072 gnd.n5643 gnd.n5505 240.244
R13073 gnd.n5643 gnd.n5496 240.244
R13074 gnd.n5653 gnd.n5496 240.244
R13075 gnd.n5653 gnd.n5491 240.244
R13076 gnd.n5681 gnd.n5491 240.244
R13077 gnd.n5681 gnd.n5492 240.244
R13078 gnd.n5492 gnd.n5484 240.244
R13079 gnd.n5676 gnd.n5484 240.244
R13080 gnd.n5676 gnd.n5474 240.244
R13081 gnd.n5673 gnd.n5474 240.244
R13082 gnd.n5673 gnd.n5463 240.244
R13083 gnd.n5670 gnd.n5463 240.244
R13084 gnd.n5670 gnd.n5453 240.244
R13085 gnd.n5667 gnd.n5453 240.244
R13086 gnd.n5667 gnd.n5431 240.244
R13087 gnd.n5816 gnd.n5431 240.244
R13088 gnd.n5816 gnd.n5427 240.244
R13089 gnd.n5824 gnd.n5427 240.244
R13090 gnd.n5824 gnd.n5417 240.244
R13091 gnd.n5417 gnd.n5398 240.244
R13092 gnd.n5863 gnd.n5398 240.244
R13093 gnd.n5863 gnd.n5399 240.244
R13094 gnd.n5399 gnd.n5394 240.244
R13095 gnd.n5883 gnd.n5394 240.244
R13096 gnd.n5883 gnd.n5384 240.244
R13097 gnd.n5878 gnd.n5384 240.244
R13098 gnd.n5878 gnd.n5378 240.244
R13099 gnd.n5874 gnd.n5378 240.244
R13100 gnd.n5874 gnd.n5367 240.244
R13101 gnd.n5870 gnd.n5367 240.244
R13102 gnd.n5870 gnd.n5345 240.244
R13103 gnd.n5949 gnd.n5345 240.244
R13104 gnd.n5949 gnd.n5293 240.244
R13105 gnd.n5970 gnd.n5293 240.244
R13106 gnd.n5970 gnd.n5282 240.244
R13107 gnd.n5966 gnd.n5282 240.244
R13108 gnd.n5966 gnd.n5275 240.244
R13109 gnd.n5963 gnd.n5275 240.244
R13110 gnd.n5963 gnd.n5264 240.244
R13111 gnd.n5960 gnd.n5264 240.244
R13112 gnd.n5960 gnd.n5242 240.244
R13113 gnd.n6035 gnd.n5242 240.244
R13114 gnd.n6035 gnd.n5238 240.244
R13115 gnd.n6053 gnd.n5238 240.244
R13116 gnd.n6053 gnd.n5232 240.244
R13117 gnd.n5232 gnd.n5222 240.244
R13118 gnd.n6048 gnd.n5222 240.244
R13119 gnd.n6048 gnd.n5215 240.244
R13120 gnd.n6045 gnd.n5215 240.244
R13121 gnd.n6045 gnd.n5208 240.244
R13122 gnd.n6104 gnd.n5208 240.244
R13123 gnd.n6104 gnd.n919 240.244
R13124 gnd.n6118 gnd.n919 240.244
R13125 gnd.n6118 gnd.n929 240.244
R13126 gnd.n6114 gnd.n929 240.244
R13127 gnd.n6114 gnd.n6113 240.244
R13128 gnd.n6113 gnd.n944 240.244
R13129 gnd.n6399 gnd.n944 240.244
R13130 gnd.n6399 gnd.n954 240.244
R13131 gnd.n6405 gnd.n954 240.244
R13132 gnd.n5613 gnd.n5611 240.244
R13133 gnd.n5611 gnd.n5610 240.244
R13134 gnd.n5607 gnd.n5606 240.244
R13135 gnd.n5604 gnd.n5530 240.244
R13136 gnd.n5600 gnd.n5598 240.244
R13137 gnd.n5596 gnd.n5536 240.244
R13138 gnd.n5592 gnd.n5590 240.244
R13139 gnd.n5588 gnd.n5542 240.244
R13140 gnd.n5584 gnd.n5582 240.244
R13141 gnd.n5580 gnd.n5548 240.244
R13142 gnd.n5576 gnd.n5574 240.244
R13143 gnd.n5572 gnd.n5554 240.244
R13144 gnd.n5567 gnd.n5565 240.244
R13145 gnd.n5619 gnd.n5515 240.244
R13146 gnd.n5629 gnd.n5515 240.244
R13147 gnd.n5629 gnd.n5511 240.244
R13148 gnd.n5635 gnd.n5511 240.244
R13149 gnd.n5635 gnd.n5503 240.244
R13150 gnd.n5645 gnd.n5503 240.244
R13151 gnd.n5645 gnd.n5499 240.244
R13152 gnd.n5651 gnd.n5499 240.244
R13153 gnd.n5651 gnd.n5490 240.244
R13154 gnd.n5743 gnd.n5490 240.244
R13155 gnd.n5743 gnd.n5485 240.244
R13156 gnd.n5750 gnd.n5485 240.244
R13157 gnd.n5750 gnd.n5476 240.244
R13158 gnd.n5760 gnd.n5476 240.244
R13159 gnd.n5760 gnd.n5462 240.244
R13160 gnd.n5775 gnd.n5462 240.244
R13161 gnd.n5775 gnd.n5455 240.244
R13162 gnd.n5790 gnd.n5455 240.244
R13163 gnd.n5790 gnd.n5456 240.244
R13164 gnd.n5456 gnd.n5434 240.244
R13165 gnd.n5814 gnd.n5434 240.244
R13166 gnd.n5814 gnd.n5435 240.244
R13167 gnd.n5435 gnd.n5415 240.244
R13168 gnd.n5841 gnd.n5415 240.244
R13169 gnd.n5841 gnd.n5402 240.244
R13170 gnd.n5861 gnd.n5402 240.244
R13171 gnd.n5861 gnd.n5403 240.244
R13172 gnd.n5857 gnd.n5403 240.244
R13173 gnd.n5857 gnd.n5383 240.244
R13174 gnd.n5899 gnd.n5383 240.244
R13175 gnd.n5899 gnd.n5376 240.244
R13176 gnd.n5910 gnd.n5376 240.244
R13177 gnd.n5910 gnd.n5369 240.244
R13178 gnd.n5925 gnd.n5369 240.244
R13179 gnd.n5925 gnd.n5370 240.244
R13180 gnd.n5370 gnd.n5348 240.244
R13181 gnd.n5947 gnd.n5348 240.244
R13182 gnd.n5947 gnd.n5349 240.244
R13183 gnd.n5349 gnd.n5280 240.244
R13184 gnd.n5984 gnd.n5280 240.244
R13185 gnd.n5984 gnd.n5273 240.244
R13186 gnd.n5995 gnd.n5273 240.244
R13187 gnd.n5995 gnd.n5266 240.244
R13188 gnd.n6009 gnd.n5266 240.244
R13189 gnd.n6009 gnd.n5267 240.244
R13190 gnd.n5267 gnd.n5246 240.244
R13191 gnd.n6033 gnd.n5246 240.244
R13192 gnd.n6033 gnd.n5236 240.244
R13193 gnd.n6055 gnd.n5236 240.244
R13194 gnd.n6055 gnd.n5221 240.244
R13195 gnd.n6079 gnd.n5221 240.244
R13196 gnd.n6079 gnd.n5212 240.244
R13197 gnd.n6091 gnd.n5212 240.244
R13198 gnd.n6092 gnd.n6091 240.244
R13199 gnd.n6093 gnd.n6092 240.244
R13200 gnd.n6093 gnd.n921 240.244
R13201 gnd.n6518 gnd.n921 240.244
R13202 gnd.n6518 gnd.n922 240.244
R13203 gnd.n6514 gnd.n922 240.244
R13204 gnd.n6514 gnd.n928 240.244
R13205 gnd.n946 gnd.n928 240.244
R13206 gnd.n6504 gnd.n946 240.244
R13207 gnd.n6504 gnd.n947 240.244
R13208 gnd.n6500 gnd.n947 240.244
R13209 gnd.n6500 gnd.n953 240.244
R13210 gnd.n7581 gnd.n7580 240.244
R13211 gnd.n7586 gnd.n7583 240.244
R13212 gnd.n7589 gnd.n7588 240.244
R13213 gnd.n7594 gnd.n7591 240.244
R13214 gnd.n7597 gnd.n7596 240.244
R13215 gnd.n7602 gnd.n7599 240.244
R13216 gnd.n7605 gnd.n7604 240.244
R13217 gnd.n7610 gnd.n7607 240.244
R13218 gnd.n7616 gnd.n7612 240.244
R13219 gnd.n4479 gnd.n1479 240.244
R13220 gnd.n4486 gnd.n1479 240.244
R13221 gnd.n4486 gnd.n1492 240.244
R13222 gnd.n1623 gnd.n1492 240.244
R13223 gnd.n4529 gnd.n1623 240.244
R13224 gnd.n4529 gnd.n1618 240.244
R13225 gnd.n4536 gnd.n1618 240.244
R13226 gnd.n4536 gnd.n1607 240.244
R13227 gnd.n1607 gnd.n1596 240.244
R13228 gnd.n4561 gnd.n1596 240.244
R13229 gnd.n4561 gnd.n1591 240.244
R13230 gnd.n4568 gnd.n1591 240.244
R13231 gnd.n4568 gnd.n1580 240.244
R13232 gnd.n1580 gnd.n1567 240.244
R13233 gnd.n4600 gnd.n1567 240.244
R13234 gnd.n4600 gnd.n1562 240.244
R13235 gnd.n4610 gnd.n1562 240.244
R13236 gnd.n4610 gnd.n1527 240.244
R13237 gnd.n4604 gnd.n1527 240.244
R13238 gnd.n4604 gnd.n1519 240.244
R13239 gnd.n4626 gnd.n1519 240.244
R13240 gnd.n4626 gnd.n279 240.244
R13241 gnd.n4635 gnd.n279 240.244
R13242 gnd.n4635 gnd.n1551 240.244
R13243 gnd.n1551 gnd.n1543 240.244
R13244 gnd.n4646 gnd.n1543 240.244
R13245 gnd.n4646 gnd.n70 240.244
R13246 gnd.n71 gnd.n70 240.244
R13247 gnd.n72 gnd.n71 240.244
R13248 gnd.n305 gnd.n72 240.244
R13249 gnd.n305 gnd.n75 240.244
R13250 gnd.n76 gnd.n75 240.244
R13251 gnd.n77 gnd.n76 240.244
R13252 gnd.n7412 gnd.n77 240.244
R13253 gnd.n7412 gnd.n80 240.244
R13254 gnd.n81 gnd.n80 240.244
R13255 gnd.n82 gnd.n81 240.244
R13256 gnd.n7456 gnd.n82 240.244
R13257 gnd.n7456 gnd.n85 240.244
R13258 gnd.n86 gnd.n85 240.244
R13259 gnd.n87 gnd.n86 240.244
R13260 gnd.n217 gnd.n87 240.244
R13261 gnd.n217 gnd.n90 240.244
R13262 gnd.n91 gnd.n90 240.244
R13263 gnd.n92 gnd.n91 240.244
R13264 gnd.n210 gnd.n92 240.244
R13265 gnd.n210 gnd.n95 240.244
R13266 gnd.n96 gnd.n95 240.244
R13267 gnd.n97 gnd.n96 240.244
R13268 gnd.n185 gnd.n97 240.244
R13269 gnd.n185 gnd.n100 240.244
R13270 gnd.n101 gnd.n100 240.244
R13271 gnd.n7744 gnd.n101 240.244
R13272 gnd.n1705 gnd.n1682 240.244
R13273 gnd.n1709 gnd.n1707 240.244
R13274 gnd.n1724 gnd.n1673 240.244
R13275 gnd.n1728 gnd.n1726 240.244
R13276 gnd.n1743 gnd.n1664 240.244
R13277 gnd.n1747 gnd.n1745 240.244
R13278 gnd.n1762 gnd.n1655 240.244
R13279 gnd.n1766 gnd.n1764 240.244
R13280 gnd.n4478 gnd.n1644 240.244
R13281 gnd.n1688 gnd.n1481 240.244
R13282 gnd.n1494 gnd.n1481 240.244
R13283 gnd.n4717 gnd.n1494 240.244
R13284 gnd.n4717 gnd.n1495 240.244
R13285 gnd.n1500 gnd.n1495 240.244
R13286 gnd.n1501 gnd.n1500 240.244
R13287 gnd.n1502 gnd.n1501 240.244
R13288 gnd.n4549 gnd.n1502 240.244
R13289 gnd.n4549 gnd.n1505 240.244
R13290 gnd.n1506 gnd.n1505 240.244
R13291 gnd.n1507 gnd.n1506 240.244
R13292 gnd.n4569 gnd.n1507 240.244
R13293 gnd.n4569 gnd.n1510 240.244
R13294 gnd.n1511 gnd.n1510 240.244
R13295 gnd.n1512 gnd.n1511 240.244
R13296 gnd.n1571 gnd.n1512 240.244
R13297 gnd.n1571 gnd.n1515 240.244
R13298 gnd.n1516 gnd.n1515 240.244
R13299 gnd.n1517 gnd.n1516 240.244
R13300 gnd.n4688 gnd.n1517 240.244
R13301 gnd.n4688 gnd.n281 240.244
R13302 gnd.n7500 gnd.n281 240.244
R13303 gnd.n7500 gnd.n282 240.244
R13304 gnd.n287 gnd.n282 240.244
R13305 gnd.n288 gnd.n287 240.244
R13306 gnd.n289 gnd.n288 240.244
R13307 gnd.n4647 gnd.n289 240.244
R13308 gnd.n4647 gnd.n293 240.244
R13309 gnd.n7486 gnd.n293 240.244
R13310 gnd.n7486 gnd.n262 240.244
R13311 gnd.n7509 gnd.n262 240.244
R13312 gnd.n7509 gnd.n258 240.244
R13313 gnd.n7515 gnd.n258 240.244
R13314 gnd.n7515 gnd.n246 240.244
R13315 gnd.n7525 gnd.n246 240.244
R13316 gnd.n7525 gnd.n242 240.244
R13317 gnd.n7531 gnd.n242 240.244
R13318 gnd.n7531 gnd.n231 240.244
R13319 gnd.n7541 gnd.n231 240.244
R13320 gnd.n7541 gnd.n227 240.244
R13321 gnd.n7547 gnd.n227 240.244
R13322 gnd.n7547 gnd.n216 240.244
R13323 gnd.n7557 gnd.n216 240.244
R13324 gnd.n7557 gnd.n212 240.244
R13325 gnd.n7563 gnd.n212 240.244
R13326 gnd.n7563 gnd.n201 240.244
R13327 gnd.n7573 gnd.n201 240.244
R13328 gnd.n7573 gnd.n195 240.244
R13329 gnd.n7654 gnd.n195 240.244
R13330 gnd.n7654 gnd.n196 240.244
R13331 gnd.n196 gnd.n187 240.244
R13332 gnd.n7578 gnd.n187 240.244
R13333 gnd.n7578 gnd.n107 240.244
R13334 gnd.n2731 gnd.n1324 240.244
R13335 gnd.n2734 gnd.n2733 240.244
R13336 gnd.n2744 gnd.n2736 240.244
R13337 gnd.n2747 gnd.n2746 240.244
R13338 gnd.n2756 gnd.n2755 240.244
R13339 gnd.n2767 gnd.n2758 240.244
R13340 gnd.n2770 gnd.n2769 240.244
R13341 gnd.n2779 gnd.n2778 240.244
R13342 gnd.n2790 gnd.n2781 240.244
R13343 gnd.n3101 gnd.n3020 240.244
R13344 gnd.n3102 gnd.n3101 240.244
R13345 gnd.n3102 gnd.n1064 240.244
R13346 gnd.n3105 gnd.n1064 240.244
R13347 gnd.n3105 gnd.n1076 240.244
R13348 gnd.n3110 gnd.n1076 240.244
R13349 gnd.n3110 gnd.n1087 240.244
R13350 gnd.n3113 gnd.n1087 240.244
R13351 gnd.n3113 gnd.n1097 240.244
R13352 gnd.n3118 gnd.n1097 240.244
R13353 gnd.n3118 gnd.n1107 240.244
R13354 gnd.n3142 gnd.n1107 240.244
R13355 gnd.n3142 gnd.n1118 240.244
R13356 gnd.n3148 gnd.n1118 240.244
R13357 gnd.n3148 gnd.n1129 240.244
R13358 gnd.n3158 gnd.n1129 240.244
R13359 gnd.n3158 gnd.n1140 240.244
R13360 gnd.n3164 gnd.n1140 240.244
R13361 gnd.n3164 gnd.n1150 240.244
R13362 gnd.n3174 gnd.n1150 240.244
R13363 gnd.n3174 gnd.n1160 240.244
R13364 gnd.n3180 gnd.n1160 240.244
R13365 gnd.n3180 gnd.n1171 240.244
R13366 gnd.n3190 gnd.n1171 240.244
R13367 gnd.n3190 gnd.n1180 240.244
R13368 gnd.n3197 gnd.n1180 240.244
R13369 gnd.n3197 gnd.n1190 240.244
R13370 gnd.n3208 gnd.n1190 240.244
R13371 gnd.n3208 gnd.n1197 240.244
R13372 gnd.n3214 gnd.n1197 240.244
R13373 gnd.n3214 gnd.n1208 240.244
R13374 gnd.n3224 gnd.n1208 240.244
R13375 gnd.n3224 gnd.n1218 240.244
R13376 gnd.n3230 gnd.n1218 240.244
R13377 gnd.n3230 gnd.n1228 240.244
R13378 gnd.n3240 gnd.n1228 240.244
R13379 gnd.n3240 gnd.n1238 240.244
R13380 gnd.n3246 gnd.n1238 240.244
R13381 gnd.n3246 gnd.n1249 240.244
R13382 gnd.n3257 gnd.n1249 240.244
R13383 gnd.n3257 gnd.n1260 240.244
R13384 gnd.n3263 gnd.n1260 240.244
R13385 gnd.n3263 gnd.n1270 240.244
R13386 gnd.n3298 gnd.n1270 240.244
R13387 gnd.n3298 gnd.n1280 240.244
R13388 gnd.n2863 gnd.n1280 240.244
R13389 gnd.n2863 gnd.n1291 240.244
R13390 gnd.n2864 gnd.n1291 240.244
R13391 gnd.n2864 gnd.n1302 240.244
R13392 gnd.n3286 gnd.n1302 240.244
R13393 gnd.n3286 gnd.n1313 240.244
R13394 gnd.n3449 gnd.n1313 240.244
R13395 gnd.n3449 gnd.n1322 240.244
R13396 gnd.n3081 gnd.n3080 240.244
R13397 gnd.n3077 gnd.n3076 240.244
R13398 gnd.n3073 gnd.n3072 240.244
R13399 gnd.n3069 gnd.n3068 240.244
R13400 gnd.n3065 gnd.n3064 240.244
R13401 gnd.n3061 gnd.n3060 240.244
R13402 gnd.n3057 gnd.n3056 240.244
R13403 gnd.n3053 gnd.n3052 240.244
R13404 gnd.n3040 gnd.n1008 240.244
R13405 gnd.n3093 gnd.n3021 240.244
R13406 gnd.n3093 gnd.n3022 240.244
R13407 gnd.n3022 gnd.n1066 240.244
R13408 gnd.n1078 gnd.n1066 240.244
R13409 gnd.n5044 gnd.n1078 240.244
R13410 gnd.n5044 gnd.n1079 240.244
R13411 gnd.n5040 gnd.n1079 240.244
R13412 gnd.n5040 gnd.n1085 240.244
R13413 gnd.n5032 gnd.n1085 240.244
R13414 gnd.n5032 gnd.n1098 240.244
R13415 gnd.n5028 gnd.n1098 240.244
R13416 gnd.n5028 gnd.n1104 240.244
R13417 gnd.n5020 gnd.n1104 240.244
R13418 gnd.n5020 gnd.n1120 240.244
R13419 gnd.n5016 gnd.n1120 240.244
R13420 gnd.n5016 gnd.n1126 240.244
R13421 gnd.n5008 gnd.n1126 240.244
R13422 gnd.n5008 gnd.n1141 240.244
R13423 gnd.n5004 gnd.n1141 240.244
R13424 gnd.n5004 gnd.n1147 240.244
R13425 gnd.n4996 gnd.n1147 240.244
R13426 gnd.n4996 gnd.n1162 240.244
R13427 gnd.n4992 gnd.n1162 240.244
R13428 gnd.n4992 gnd.n1168 240.244
R13429 gnd.n4984 gnd.n1168 240.244
R13430 gnd.n4984 gnd.n1181 240.244
R13431 gnd.n4980 gnd.n1181 240.244
R13432 gnd.n4980 gnd.n1187 240.244
R13433 gnd.n4971 gnd.n1187 240.244
R13434 gnd.n4971 gnd.n1199 240.244
R13435 gnd.n4967 gnd.n1199 240.244
R13436 gnd.n4967 gnd.n1205 240.244
R13437 gnd.n4959 gnd.n1205 240.244
R13438 gnd.n4959 gnd.n1219 240.244
R13439 gnd.n4955 gnd.n1219 240.244
R13440 gnd.n4955 gnd.n1225 240.244
R13441 gnd.n4947 gnd.n1225 240.244
R13442 gnd.n4947 gnd.n1240 240.244
R13443 gnd.n4943 gnd.n1240 240.244
R13444 gnd.n4943 gnd.n1246 240.244
R13445 gnd.n4935 gnd.n1246 240.244
R13446 gnd.n4935 gnd.n1261 240.244
R13447 gnd.n4931 gnd.n1261 240.244
R13448 gnd.n4931 gnd.n1267 240.244
R13449 gnd.n4923 gnd.n1267 240.244
R13450 gnd.n4923 gnd.n1282 240.244
R13451 gnd.n4919 gnd.n1282 240.244
R13452 gnd.n4919 gnd.n1288 240.244
R13453 gnd.n4911 gnd.n1288 240.244
R13454 gnd.n4911 gnd.n1304 240.244
R13455 gnd.n4907 gnd.n1304 240.244
R13456 gnd.n4907 gnd.n1310 240.244
R13457 gnd.n4899 gnd.n1310 240.244
R13458 gnd.n6698 gnd.n739 240.244
R13459 gnd.n6698 gnd.n735 240.244
R13460 gnd.n6704 gnd.n735 240.244
R13461 gnd.n6704 gnd.n733 240.244
R13462 gnd.n6708 gnd.n733 240.244
R13463 gnd.n6708 gnd.n729 240.244
R13464 gnd.n6714 gnd.n729 240.244
R13465 gnd.n6714 gnd.n727 240.244
R13466 gnd.n6718 gnd.n727 240.244
R13467 gnd.n6718 gnd.n723 240.244
R13468 gnd.n6724 gnd.n723 240.244
R13469 gnd.n6724 gnd.n721 240.244
R13470 gnd.n6728 gnd.n721 240.244
R13471 gnd.n6728 gnd.n717 240.244
R13472 gnd.n6734 gnd.n717 240.244
R13473 gnd.n6734 gnd.n715 240.244
R13474 gnd.n6738 gnd.n715 240.244
R13475 gnd.n6738 gnd.n711 240.244
R13476 gnd.n6744 gnd.n711 240.244
R13477 gnd.n6744 gnd.n709 240.244
R13478 gnd.n6748 gnd.n709 240.244
R13479 gnd.n6748 gnd.n705 240.244
R13480 gnd.n6754 gnd.n705 240.244
R13481 gnd.n6754 gnd.n703 240.244
R13482 gnd.n6758 gnd.n703 240.244
R13483 gnd.n6758 gnd.n699 240.244
R13484 gnd.n6764 gnd.n699 240.244
R13485 gnd.n6764 gnd.n697 240.244
R13486 gnd.n6768 gnd.n697 240.244
R13487 gnd.n6768 gnd.n693 240.244
R13488 gnd.n6774 gnd.n693 240.244
R13489 gnd.n6774 gnd.n691 240.244
R13490 gnd.n6778 gnd.n691 240.244
R13491 gnd.n6778 gnd.n687 240.244
R13492 gnd.n6784 gnd.n687 240.244
R13493 gnd.n6784 gnd.n685 240.244
R13494 gnd.n6788 gnd.n685 240.244
R13495 gnd.n6788 gnd.n681 240.244
R13496 gnd.n6794 gnd.n681 240.244
R13497 gnd.n6794 gnd.n679 240.244
R13498 gnd.n6798 gnd.n679 240.244
R13499 gnd.n6798 gnd.n675 240.244
R13500 gnd.n6804 gnd.n675 240.244
R13501 gnd.n6804 gnd.n673 240.244
R13502 gnd.n6808 gnd.n673 240.244
R13503 gnd.n6808 gnd.n669 240.244
R13504 gnd.n6814 gnd.n669 240.244
R13505 gnd.n6814 gnd.n667 240.244
R13506 gnd.n6818 gnd.n667 240.244
R13507 gnd.n6818 gnd.n663 240.244
R13508 gnd.n6824 gnd.n663 240.244
R13509 gnd.n6824 gnd.n661 240.244
R13510 gnd.n6828 gnd.n661 240.244
R13511 gnd.n6828 gnd.n657 240.244
R13512 gnd.n6834 gnd.n657 240.244
R13513 gnd.n6834 gnd.n655 240.244
R13514 gnd.n6838 gnd.n655 240.244
R13515 gnd.n6838 gnd.n651 240.244
R13516 gnd.n6844 gnd.n651 240.244
R13517 gnd.n6844 gnd.n649 240.244
R13518 gnd.n6848 gnd.n649 240.244
R13519 gnd.n6848 gnd.n645 240.244
R13520 gnd.n6854 gnd.n645 240.244
R13521 gnd.n6854 gnd.n643 240.244
R13522 gnd.n6858 gnd.n643 240.244
R13523 gnd.n6858 gnd.n639 240.244
R13524 gnd.n6864 gnd.n639 240.244
R13525 gnd.n6864 gnd.n637 240.244
R13526 gnd.n6868 gnd.n637 240.244
R13527 gnd.n6868 gnd.n633 240.244
R13528 gnd.n6874 gnd.n633 240.244
R13529 gnd.n6874 gnd.n631 240.244
R13530 gnd.n6878 gnd.n631 240.244
R13531 gnd.n6878 gnd.n627 240.244
R13532 gnd.n6884 gnd.n627 240.244
R13533 gnd.n6884 gnd.n625 240.244
R13534 gnd.n6888 gnd.n625 240.244
R13535 gnd.n6888 gnd.n621 240.244
R13536 gnd.n6894 gnd.n621 240.244
R13537 gnd.n6894 gnd.n619 240.244
R13538 gnd.n6898 gnd.n619 240.244
R13539 gnd.n6898 gnd.n615 240.244
R13540 gnd.n6904 gnd.n615 240.244
R13541 gnd.n6904 gnd.n613 240.244
R13542 gnd.n6908 gnd.n613 240.244
R13543 gnd.n6908 gnd.n609 240.244
R13544 gnd.n6914 gnd.n609 240.244
R13545 gnd.n6914 gnd.n607 240.244
R13546 gnd.n6918 gnd.n607 240.244
R13547 gnd.n6918 gnd.n603 240.244
R13548 gnd.n6924 gnd.n603 240.244
R13549 gnd.n6924 gnd.n601 240.244
R13550 gnd.n6928 gnd.n601 240.244
R13551 gnd.n6928 gnd.n597 240.244
R13552 gnd.n6934 gnd.n597 240.244
R13553 gnd.n6934 gnd.n595 240.244
R13554 gnd.n6938 gnd.n595 240.244
R13555 gnd.n6938 gnd.n591 240.244
R13556 gnd.n6944 gnd.n591 240.244
R13557 gnd.n6944 gnd.n589 240.244
R13558 gnd.n6948 gnd.n589 240.244
R13559 gnd.n6948 gnd.n585 240.244
R13560 gnd.n6954 gnd.n585 240.244
R13561 gnd.n6954 gnd.n583 240.244
R13562 gnd.n6958 gnd.n583 240.244
R13563 gnd.n6958 gnd.n579 240.244
R13564 gnd.n6964 gnd.n579 240.244
R13565 gnd.n6964 gnd.n577 240.244
R13566 gnd.n6968 gnd.n577 240.244
R13567 gnd.n6968 gnd.n573 240.244
R13568 gnd.n6974 gnd.n573 240.244
R13569 gnd.n6974 gnd.n571 240.244
R13570 gnd.n6978 gnd.n571 240.244
R13571 gnd.n6978 gnd.n567 240.244
R13572 gnd.n6984 gnd.n567 240.244
R13573 gnd.n6984 gnd.n565 240.244
R13574 gnd.n6988 gnd.n565 240.244
R13575 gnd.n6988 gnd.n561 240.244
R13576 gnd.n6994 gnd.n561 240.244
R13577 gnd.n6994 gnd.n559 240.244
R13578 gnd.n6998 gnd.n559 240.244
R13579 gnd.n6998 gnd.n555 240.244
R13580 gnd.n7004 gnd.n555 240.244
R13581 gnd.n7004 gnd.n553 240.244
R13582 gnd.n7008 gnd.n553 240.244
R13583 gnd.n7008 gnd.n549 240.244
R13584 gnd.n7014 gnd.n549 240.244
R13585 gnd.n7014 gnd.n547 240.244
R13586 gnd.n7018 gnd.n547 240.244
R13587 gnd.n7018 gnd.n543 240.244
R13588 gnd.n7024 gnd.n543 240.244
R13589 gnd.n7024 gnd.n541 240.244
R13590 gnd.n7028 gnd.n541 240.244
R13591 gnd.n7028 gnd.n537 240.244
R13592 gnd.n7034 gnd.n537 240.244
R13593 gnd.n7034 gnd.n535 240.244
R13594 gnd.n7038 gnd.n535 240.244
R13595 gnd.n7038 gnd.n531 240.244
R13596 gnd.n7044 gnd.n531 240.244
R13597 gnd.n7044 gnd.n529 240.244
R13598 gnd.n7048 gnd.n529 240.244
R13599 gnd.n7048 gnd.n525 240.244
R13600 gnd.n7054 gnd.n525 240.244
R13601 gnd.n7054 gnd.n523 240.244
R13602 gnd.n7058 gnd.n523 240.244
R13603 gnd.n7058 gnd.n519 240.244
R13604 gnd.n7064 gnd.n519 240.244
R13605 gnd.n7064 gnd.n517 240.244
R13606 gnd.n7068 gnd.n517 240.244
R13607 gnd.n7068 gnd.n513 240.244
R13608 gnd.n7074 gnd.n513 240.244
R13609 gnd.n7074 gnd.n511 240.244
R13610 gnd.n7078 gnd.n511 240.244
R13611 gnd.n7078 gnd.n507 240.244
R13612 gnd.n7084 gnd.n507 240.244
R13613 gnd.n7084 gnd.n505 240.244
R13614 gnd.n7088 gnd.n505 240.244
R13615 gnd.n7088 gnd.n501 240.244
R13616 gnd.n7094 gnd.n501 240.244
R13617 gnd.n7094 gnd.n499 240.244
R13618 gnd.n7098 gnd.n499 240.244
R13619 gnd.n7098 gnd.n495 240.244
R13620 gnd.n7104 gnd.n495 240.244
R13621 gnd.n7104 gnd.n493 240.244
R13622 gnd.n7108 gnd.n493 240.244
R13623 gnd.n7108 gnd.n489 240.244
R13624 gnd.n7114 gnd.n489 240.244
R13625 gnd.n7114 gnd.n487 240.244
R13626 gnd.n7118 gnd.n487 240.244
R13627 gnd.n7118 gnd.n483 240.244
R13628 gnd.n7124 gnd.n483 240.244
R13629 gnd.n7124 gnd.n481 240.244
R13630 gnd.n7128 gnd.n481 240.244
R13631 gnd.n7128 gnd.n477 240.244
R13632 gnd.n7134 gnd.n477 240.244
R13633 gnd.n7134 gnd.n475 240.244
R13634 gnd.n7138 gnd.n475 240.244
R13635 gnd.n7138 gnd.n471 240.244
R13636 gnd.n7144 gnd.n471 240.244
R13637 gnd.n7144 gnd.n469 240.244
R13638 gnd.n7148 gnd.n469 240.244
R13639 gnd.n7148 gnd.n465 240.244
R13640 gnd.n7154 gnd.n465 240.244
R13641 gnd.n7154 gnd.n463 240.244
R13642 gnd.n7158 gnd.n463 240.244
R13643 gnd.n7158 gnd.n459 240.244
R13644 gnd.n7164 gnd.n459 240.244
R13645 gnd.n7164 gnd.n457 240.244
R13646 gnd.n7168 gnd.n457 240.244
R13647 gnd.n7168 gnd.n453 240.244
R13648 gnd.n7175 gnd.n453 240.244
R13649 gnd.n7175 gnd.n451 240.244
R13650 gnd.n7179 gnd.n451 240.244
R13651 gnd.n7179 gnd.n448 240.244
R13652 gnd.n7185 gnd.n446 240.244
R13653 gnd.n7189 gnd.n446 240.244
R13654 gnd.n7189 gnd.n442 240.244
R13655 gnd.n7195 gnd.n442 240.244
R13656 gnd.n7195 gnd.n440 240.244
R13657 gnd.n7199 gnd.n440 240.244
R13658 gnd.n7199 gnd.n436 240.244
R13659 gnd.n7205 gnd.n436 240.244
R13660 gnd.n7205 gnd.n434 240.244
R13661 gnd.n7209 gnd.n434 240.244
R13662 gnd.n7209 gnd.n430 240.244
R13663 gnd.n7215 gnd.n430 240.244
R13664 gnd.n7215 gnd.n428 240.244
R13665 gnd.n7219 gnd.n428 240.244
R13666 gnd.n7219 gnd.n424 240.244
R13667 gnd.n7225 gnd.n424 240.244
R13668 gnd.n7225 gnd.n422 240.244
R13669 gnd.n7229 gnd.n422 240.244
R13670 gnd.n7229 gnd.n418 240.244
R13671 gnd.n7235 gnd.n418 240.244
R13672 gnd.n7235 gnd.n416 240.244
R13673 gnd.n7239 gnd.n416 240.244
R13674 gnd.n7239 gnd.n412 240.244
R13675 gnd.n7245 gnd.n412 240.244
R13676 gnd.n7245 gnd.n410 240.244
R13677 gnd.n7249 gnd.n410 240.244
R13678 gnd.n7249 gnd.n406 240.244
R13679 gnd.n7255 gnd.n406 240.244
R13680 gnd.n7255 gnd.n404 240.244
R13681 gnd.n7259 gnd.n404 240.244
R13682 gnd.n7259 gnd.n400 240.244
R13683 gnd.n7265 gnd.n400 240.244
R13684 gnd.n7265 gnd.n398 240.244
R13685 gnd.n7269 gnd.n398 240.244
R13686 gnd.n7269 gnd.n394 240.244
R13687 gnd.n7275 gnd.n394 240.244
R13688 gnd.n7275 gnd.n392 240.244
R13689 gnd.n7279 gnd.n392 240.244
R13690 gnd.n7279 gnd.n388 240.244
R13691 gnd.n7285 gnd.n388 240.244
R13692 gnd.n7285 gnd.n386 240.244
R13693 gnd.n7289 gnd.n386 240.244
R13694 gnd.n7289 gnd.n382 240.244
R13695 gnd.n7295 gnd.n382 240.244
R13696 gnd.n7295 gnd.n380 240.244
R13697 gnd.n7299 gnd.n380 240.244
R13698 gnd.n7299 gnd.n376 240.244
R13699 gnd.n7305 gnd.n376 240.244
R13700 gnd.n7305 gnd.n374 240.244
R13701 gnd.n7309 gnd.n374 240.244
R13702 gnd.n7309 gnd.n370 240.244
R13703 gnd.n7315 gnd.n370 240.244
R13704 gnd.n7315 gnd.n368 240.244
R13705 gnd.n7319 gnd.n368 240.244
R13706 gnd.n7319 gnd.n364 240.244
R13707 gnd.n7325 gnd.n364 240.244
R13708 gnd.n7325 gnd.n362 240.244
R13709 gnd.n7329 gnd.n362 240.244
R13710 gnd.n7329 gnd.n358 240.244
R13711 gnd.n7335 gnd.n358 240.244
R13712 gnd.n7335 gnd.n356 240.244
R13713 gnd.n7339 gnd.n356 240.244
R13714 gnd.n7339 gnd.n352 240.244
R13715 gnd.n7345 gnd.n352 240.244
R13716 gnd.n7345 gnd.n350 240.244
R13717 gnd.n7349 gnd.n350 240.244
R13718 gnd.n7349 gnd.n346 240.244
R13719 gnd.n7355 gnd.n346 240.244
R13720 gnd.n7355 gnd.n344 240.244
R13721 gnd.n7359 gnd.n344 240.244
R13722 gnd.n7359 gnd.n340 240.244
R13723 gnd.n7365 gnd.n340 240.244
R13724 gnd.n7365 gnd.n338 240.244
R13725 gnd.n7369 gnd.n338 240.244
R13726 gnd.n7369 gnd.n334 240.244
R13727 gnd.n7375 gnd.n334 240.244
R13728 gnd.n7375 gnd.n332 240.244
R13729 gnd.n7379 gnd.n332 240.244
R13730 gnd.n7379 gnd.n328 240.244
R13731 gnd.n7385 gnd.n328 240.244
R13732 gnd.n7385 gnd.n326 240.244
R13733 gnd.n7390 gnd.n326 240.244
R13734 gnd.n7390 gnd.n322 240.244
R13735 gnd.n7397 gnd.n322 240.244
R13736 gnd.n2929 gnd.n2920 240.244
R13737 gnd.n2930 gnd.n2929 240.244
R13738 gnd.n2931 gnd.n2930 240.244
R13739 gnd.n2931 gnd.n2915 240.244
R13740 gnd.n3004 gnd.n2915 240.244
R13741 gnd.n3004 gnd.n2916 240.244
R13742 gnd.n3000 gnd.n2916 240.244
R13743 gnd.n3000 gnd.n2999 240.244
R13744 gnd.n2999 gnd.n2998 240.244
R13745 gnd.n2998 gnd.n2939 240.244
R13746 gnd.n2991 gnd.n2939 240.244
R13747 gnd.n2991 gnd.n2990 240.244
R13748 gnd.n2990 gnd.n2989 240.244
R13749 gnd.n2989 gnd.n2987 240.244
R13750 gnd.n2987 gnd.n2984 240.244
R13751 gnd.n2984 gnd.n2983 240.244
R13752 gnd.n2983 gnd.n2980 240.244
R13753 gnd.n2980 gnd.n2979 240.244
R13754 gnd.n2979 gnd.n2946 240.244
R13755 gnd.n2975 gnd.n2946 240.244
R13756 gnd.n2975 gnd.n2974 240.244
R13757 gnd.n2974 gnd.n2973 240.244
R13758 gnd.n2973 gnd.n2949 240.244
R13759 gnd.n2969 gnd.n2949 240.244
R13760 gnd.n2969 gnd.n2968 240.244
R13761 gnd.n2968 gnd.n2967 240.244
R13762 gnd.n2967 gnd.n2955 240.244
R13763 gnd.n2963 gnd.n2955 240.244
R13764 gnd.n2963 gnd.n2962 240.244
R13765 gnd.n2962 gnd.n2857 240.244
R13766 gnd.n3301 gnd.n2857 240.244
R13767 gnd.n3301 gnd.n2853 240.244
R13768 gnd.n3307 gnd.n2853 240.244
R13769 gnd.n3308 gnd.n3307 240.244
R13770 gnd.n3309 gnd.n3308 240.244
R13771 gnd.n3309 gnd.n2849 240.244
R13772 gnd.n3315 gnd.n2849 240.244
R13773 gnd.n3316 gnd.n3315 240.244
R13774 gnd.n3317 gnd.n3316 240.244
R13775 gnd.n3317 gnd.n2845 240.244
R13776 gnd.n3323 gnd.n2845 240.244
R13777 gnd.n3324 gnd.n3323 240.244
R13778 gnd.n3328 gnd.n3324 240.244
R13779 gnd.n3328 gnd.n2841 240.244
R13780 gnd.n3334 gnd.n2841 240.244
R13781 gnd.n3334 gnd.n2707 240.244
R13782 gnd.n3341 gnd.n2707 240.244
R13783 gnd.n3341 gnd.n2703 240.244
R13784 gnd.n3347 gnd.n2703 240.244
R13785 gnd.n3347 gnd.n2701 240.244
R13786 gnd.n3357 gnd.n2701 240.244
R13787 gnd.n3357 gnd.n2697 240.244
R13788 gnd.n3363 gnd.n2697 240.244
R13789 gnd.n3363 gnd.n2695 240.244
R13790 gnd.n3373 gnd.n2695 240.244
R13791 gnd.n3373 gnd.n2691 240.244
R13792 gnd.n3379 gnd.n2691 240.244
R13793 gnd.n3379 gnd.n2689 240.244
R13794 gnd.n3389 gnd.n2689 240.244
R13795 gnd.n3389 gnd.n2685 240.244
R13796 gnd.n3395 gnd.n2685 240.244
R13797 gnd.n3395 gnd.n2386 240.244
R13798 gnd.n3565 gnd.n2386 240.244
R13799 gnd.n3565 gnd.n2382 240.244
R13800 gnd.n3571 gnd.n2382 240.244
R13801 gnd.n3571 gnd.n2364 240.244
R13802 gnd.n3593 gnd.n2364 240.244
R13803 gnd.n3593 gnd.n2359 240.244
R13804 gnd.n3601 gnd.n2359 240.244
R13805 gnd.n3601 gnd.n2360 240.244
R13806 gnd.n2360 gnd.n2336 240.244
R13807 gnd.n3667 gnd.n2336 240.244
R13808 gnd.n3667 gnd.n2332 240.244
R13809 gnd.n3673 gnd.n2332 240.244
R13810 gnd.n3673 gnd.n2316 240.244
R13811 gnd.n3692 gnd.n2316 240.244
R13812 gnd.n3692 gnd.n2312 240.244
R13813 gnd.n3698 gnd.n2312 240.244
R13814 gnd.n3698 gnd.n2296 240.244
R13815 gnd.n3726 gnd.n2296 240.244
R13816 gnd.n3726 gnd.n2292 240.244
R13817 gnd.n3732 gnd.n2292 240.244
R13818 gnd.n3732 gnd.n2279 240.244
R13819 gnd.n3771 gnd.n2279 240.244
R13820 gnd.n3771 gnd.n2274 240.244
R13821 gnd.n3779 gnd.n2274 240.244
R13822 gnd.n3779 gnd.n2275 240.244
R13823 gnd.n2275 gnd.n2251 240.244
R13824 gnd.n3844 gnd.n2251 240.244
R13825 gnd.n3844 gnd.n2247 240.244
R13826 gnd.n3850 gnd.n2247 240.244
R13827 gnd.n3850 gnd.n2231 240.244
R13828 gnd.n3870 gnd.n2231 240.244
R13829 gnd.n3870 gnd.n2227 240.244
R13830 gnd.n3876 gnd.n2227 240.244
R13831 gnd.n3876 gnd.n2208 240.244
R13832 gnd.n3903 gnd.n2208 240.244
R13833 gnd.n3903 gnd.n2204 240.244
R13834 gnd.n3909 gnd.n2204 240.244
R13835 gnd.n3909 gnd.n2191 240.244
R13836 gnd.n3949 gnd.n2191 240.244
R13837 gnd.n3949 gnd.n2186 240.244
R13838 gnd.n3957 gnd.n2186 240.244
R13839 gnd.n3957 gnd.n2187 240.244
R13840 gnd.n2187 gnd.n2164 240.244
R13841 gnd.n4006 gnd.n2164 240.244
R13842 gnd.n4006 gnd.n2160 240.244
R13843 gnd.n4012 gnd.n2160 240.244
R13844 gnd.n4012 gnd.n2143 240.244
R13845 gnd.n4031 gnd.n2143 240.244
R13846 gnd.n4031 gnd.n2139 240.244
R13847 gnd.n4037 gnd.n2139 240.244
R13848 gnd.n4037 gnd.n2121 240.244
R13849 gnd.n4091 gnd.n2121 240.244
R13850 gnd.n4091 gnd.n2117 240.244
R13851 gnd.n4097 gnd.n2117 240.244
R13852 gnd.n4097 gnd.n2099 240.244
R13853 gnd.n4120 gnd.n2099 240.244
R13854 gnd.n4120 gnd.n2094 240.244
R13855 gnd.n4128 gnd.n2094 240.244
R13856 gnd.n4128 gnd.n2095 240.244
R13857 gnd.n2095 gnd.n2071 240.244
R13858 gnd.n4170 gnd.n2071 240.244
R13859 gnd.n4170 gnd.n2067 240.244
R13860 gnd.n4176 gnd.n2067 240.244
R13861 gnd.n4176 gnd.n2050 240.244
R13862 gnd.n4196 gnd.n2050 240.244
R13863 gnd.n4196 gnd.n2045 240.244
R13864 gnd.n4204 gnd.n2045 240.244
R13865 gnd.n4204 gnd.n2046 240.244
R13866 gnd.n2046 gnd.n1846 240.244
R13867 gnd.n4381 gnd.n1846 240.244
R13868 gnd.n4381 gnd.n1842 240.244
R13869 gnd.n4387 gnd.n1842 240.244
R13870 gnd.n4387 gnd.n1833 240.244
R13871 gnd.n4401 gnd.n1833 240.244
R13872 gnd.n4401 gnd.n1829 240.244
R13873 gnd.n4407 gnd.n1829 240.244
R13874 gnd.n4407 gnd.n1820 240.244
R13875 gnd.n4421 gnd.n1820 240.244
R13876 gnd.n4421 gnd.n1816 240.244
R13877 gnd.n4427 gnd.n1816 240.244
R13878 gnd.n4427 gnd.n1807 240.244
R13879 gnd.n4444 gnd.n1807 240.244
R13880 gnd.n4444 gnd.n1803 240.244
R13881 gnd.n4451 gnd.n1803 240.244
R13882 gnd.n4451 gnd.n1459 240.244
R13883 gnd.n4738 gnd.n1459 240.244
R13884 gnd.n4738 gnd.n1460 240.244
R13885 gnd.n4734 gnd.n1460 240.244
R13886 gnd.n4734 gnd.n1466 240.244
R13887 gnd.n4730 gnd.n1466 240.244
R13888 gnd.n4730 gnd.n1469 240.244
R13889 gnd.n4726 gnd.n1469 240.244
R13890 gnd.n4726 gnd.n1475 240.244
R13891 gnd.n1627 gnd.n1475 240.244
R13892 gnd.n1627 gnd.n1624 240.244
R13893 gnd.n1633 gnd.n1624 240.244
R13894 gnd.n1633 gnd.n1615 240.244
R13895 gnd.n4539 gnd.n1615 240.244
R13896 gnd.n4539 gnd.n1609 240.244
R13897 gnd.n4547 gnd.n1609 240.244
R13898 gnd.n4547 gnd.n1611 240.244
R13899 gnd.n1611 gnd.n1588 240.244
R13900 gnd.n4572 gnd.n1588 240.244
R13901 gnd.n4572 gnd.n1582 240.244
R13902 gnd.n4587 gnd.n1582 240.244
R13903 gnd.n4587 gnd.n1584 240.244
R13904 gnd.n4583 gnd.n1584 240.244
R13905 gnd.n4583 gnd.n4582 240.244
R13906 gnd.n4582 gnd.n1529 240.244
R13907 gnd.n4677 gnd.n1529 240.244
R13908 gnd.n4677 gnd.n1531 240.244
R13909 gnd.n4673 gnd.n1531 240.244
R13910 gnd.n4673 gnd.n4672 240.244
R13911 gnd.n4672 gnd.n4671 240.244
R13912 gnd.n4671 gnd.n1538 240.244
R13913 gnd.n4666 gnd.n1538 240.244
R13914 gnd.n4666 gnd.n1540 240.244
R13915 gnd.n4658 gnd.n1540 240.244
R13916 gnd.n4658 gnd.n4650 240.244
R13917 gnd.n4653 gnd.n4650 240.244
R13918 gnd.n4653 gnd.n306 240.244
R13919 gnd.n7472 gnd.n306 240.244
R13920 gnd.n7472 gnd.n307 240.244
R13921 gnd.n7467 gnd.n307 240.244
R13922 gnd.n7467 gnd.n7466 240.244
R13923 gnd.n7466 gnd.n7465 240.244
R13924 gnd.n7465 gnd.n311 240.244
R13925 gnd.n7461 gnd.n311 240.244
R13926 gnd.n7461 gnd.n7460 240.244
R13927 gnd.n7460 gnd.n7459 240.244
R13928 gnd.n7459 gnd.n317 240.244
R13929 gnd.n7398 gnd.n317 240.244
R13930 gnd.n6694 gnd.n741 240.244
R13931 gnd.n6690 gnd.n741 240.244
R13932 gnd.n6690 gnd.n746 240.244
R13933 gnd.n6686 gnd.n746 240.244
R13934 gnd.n6686 gnd.n748 240.244
R13935 gnd.n6682 gnd.n748 240.244
R13936 gnd.n6682 gnd.n754 240.244
R13937 gnd.n6678 gnd.n754 240.244
R13938 gnd.n6678 gnd.n756 240.244
R13939 gnd.n6674 gnd.n756 240.244
R13940 gnd.n6674 gnd.n762 240.244
R13941 gnd.n6670 gnd.n762 240.244
R13942 gnd.n6670 gnd.n764 240.244
R13943 gnd.n6666 gnd.n764 240.244
R13944 gnd.n6666 gnd.n770 240.244
R13945 gnd.n6662 gnd.n770 240.244
R13946 gnd.n6662 gnd.n772 240.244
R13947 gnd.n6658 gnd.n772 240.244
R13948 gnd.n6658 gnd.n778 240.244
R13949 gnd.n6654 gnd.n778 240.244
R13950 gnd.n6654 gnd.n780 240.244
R13951 gnd.n6650 gnd.n780 240.244
R13952 gnd.n6650 gnd.n786 240.244
R13953 gnd.n6646 gnd.n786 240.244
R13954 gnd.n6646 gnd.n788 240.244
R13955 gnd.n6642 gnd.n788 240.244
R13956 gnd.n6642 gnd.n794 240.244
R13957 gnd.n6638 gnd.n794 240.244
R13958 gnd.n6638 gnd.n796 240.244
R13959 gnd.n6634 gnd.n796 240.244
R13960 gnd.n6634 gnd.n802 240.244
R13961 gnd.n6630 gnd.n802 240.244
R13962 gnd.n6630 gnd.n804 240.244
R13963 gnd.n6626 gnd.n804 240.244
R13964 gnd.n6626 gnd.n810 240.244
R13965 gnd.n6622 gnd.n810 240.244
R13966 gnd.n6622 gnd.n812 240.244
R13967 gnd.n6618 gnd.n812 240.244
R13968 gnd.n6618 gnd.n818 240.244
R13969 gnd.n6614 gnd.n818 240.244
R13970 gnd.n6614 gnd.n820 240.244
R13971 gnd.n6610 gnd.n820 240.244
R13972 gnd.n6610 gnd.n826 240.244
R13973 gnd.n6606 gnd.n826 240.244
R13974 gnd.n6606 gnd.n828 240.244
R13975 gnd.n6602 gnd.n828 240.244
R13976 gnd.n6602 gnd.n834 240.244
R13977 gnd.n6598 gnd.n834 240.244
R13978 gnd.n6598 gnd.n836 240.244
R13979 gnd.n6594 gnd.n836 240.244
R13980 gnd.n6594 gnd.n842 240.244
R13981 gnd.n6590 gnd.n842 240.244
R13982 gnd.n6590 gnd.n844 240.244
R13983 gnd.n6586 gnd.n844 240.244
R13984 gnd.n6586 gnd.n850 240.244
R13985 gnd.n6582 gnd.n850 240.244
R13986 gnd.n6582 gnd.n852 240.244
R13987 gnd.n6578 gnd.n852 240.244
R13988 gnd.n6578 gnd.n858 240.244
R13989 gnd.n6574 gnd.n858 240.244
R13990 gnd.n6574 gnd.n860 240.244
R13991 gnd.n6570 gnd.n860 240.244
R13992 gnd.n6570 gnd.n866 240.244
R13993 gnd.n6566 gnd.n866 240.244
R13994 gnd.n6566 gnd.n868 240.244
R13995 gnd.n6562 gnd.n868 240.244
R13996 gnd.n6562 gnd.n874 240.244
R13997 gnd.n6558 gnd.n874 240.244
R13998 gnd.n6558 gnd.n876 240.244
R13999 gnd.n6554 gnd.n876 240.244
R14000 gnd.n6554 gnd.n882 240.244
R14001 gnd.n6550 gnd.n882 240.244
R14002 gnd.n6550 gnd.n884 240.244
R14003 gnd.n6546 gnd.n884 240.244
R14004 gnd.n6546 gnd.n890 240.244
R14005 gnd.n6542 gnd.n890 240.244
R14006 gnd.n6542 gnd.n892 240.244
R14007 gnd.n6538 gnd.n892 240.244
R14008 gnd.n6538 gnd.n898 240.244
R14009 gnd.n6534 gnd.n898 240.244
R14010 gnd.n6534 gnd.n900 240.244
R14011 gnd.n6530 gnd.n900 240.244
R14012 gnd.n6530 gnd.n906 240.244
R14013 gnd.n2923 gnd.n906 240.244
R14014 gnd.n1330 gnd.n1329 240.244
R14015 gnd.n1331 gnd.n1330 240.244
R14016 gnd.n3350 gnd.n1331 240.244
R14017 gnd.n3350 gnd.n1334 240.244
R14018 gnd.n1335 gnd.n1334 240.244
R14019 gnd.n1336 gnd.n1335 240.244
R14020 gnd.n3366 gnd.n1336 240.244
R14021 gnd.n3366 gnd.n1339 240.244
R14022 gnd.n1340 gnd.n1339 240.244
R14023 gnd.n1341 gnd.n1340 240.244
R14024 gnd.n3382 gnd.n1341 240.244
R14025 gnd.n3382 gnd.n1344 240.244
R14026 gnd.n1345 gnd.n1344 240.244
R14027 gnd.n1346 gnd.n1345 240.244
R14028 gnd.n3398 gnd.n1346 240.244
R14029 gnd.n3398 gnd.n1349 240.244
R14030 gnd.n1350 gnd.n1349 240.244
R14031 gnd.n1351 gnd.n1350 240.244
R14032 gnd.n2369 gnd.n1351 240.244
R14033 gnd.n2369 gnd.n1354 240.244
R14034 gnd.n1355 gnd.n1354 240.244
R14035 gnd.n1356 gnd.n1355 240.244
R14036 gnd.n3611 gnd.n1356 240.244
R14037 gnd.n3611 gnd.n1359 240.244
R14038 gnd.n1360 gnd.n1359 240.244
R14039 gnd.n1361 gnd.n1360 240.244
R14040 gnd.n2327 gnd.n1361 240.244
R14041 gnd.n2327 gnd.n1364 240.244
R14042 gnd.n1365 gnd.n1364 240.244
R14043 gnd.n1366 gnd.n1365 240.244
R14044 gnd.n3701 gnd.n1366 240.244
R14045 gnd.n3701 gnd.n1369 240.244
R14046 gnd.n1370 gnd.n1369 240.244
R14047 gnd.n1371 gnd.n1370 240.244
R14048 gnd.n2290 gnd.n1371 240.244
R14049 gnd.n2290 gnd.n1374 240.244
R14050 gnd.n1375 gnd.n1374 240.244
R14051 gnd.n1376 gnd.n1375 240.244
R14052 gnd.n3781 gnd.n1376 240.244
R14053 gnd.n3781 gnd.n1379 240.244
R14054 gnd.n1380 gnd.n1379 240.244
R14055 gnd.n1381 gnd.n1380 240.244
R14056 gnd.n3841 gnd.n1381 240.244
R14057 gnd.n3841 gnd.n1384 240.244
R14058 gnd.n1385 gnd.n1384 240.244
R14059 gnd.n1386 gnd.n1385 240.244
R14060 gnd.n3867 gnd.n1386 240.244
R14061 gnd.n3867 gnd.n1389 240.244
R14062 gnd.n1390 gnd.n1389 240.244
R14063 gnd.n1391 gnd.n1390 240.244
R14064 gnd.n2211 gnd.n1391 240.244
R14065 gnd.n2211 gnd.n1394 240.244
R14066 gnd.n1395 gnd.n1394 240.244
R14067 gnd.n1396 gnd.n1395 240.244
R14068 gnd.n2194 gnd.n1396 240.244
R14069 gnd.n2194 gnd.n1399 240.244
R14070 gnd.n1400 gnd.n1399 240.244
R14071 gnd.n1401 gnd.n1400 240.244
R14072 gnd.n3995 gnd.n1401 240.244
R14073 gnd.n3995 gnd.n1404 240.244
R14074 gnd.n1405 gnd.n1404 240.244
R14075 gnd.n1406 gnd.n1405 240.244
R14076 gnd.n2149 gnd.n1406 240.244
R14077 gnd.n2149 gnd.n1409 240.244
R14078 gnd.n1410 gnd.n1409 240.244
R14079 gnd.n1411 gnd.n1410 240.244
R14080 gnd.n2122 gnd.n1411 240.244
R14081 gnd.n2122 gnd.n1414 240.244
R14082 gnd.n1415 gnd.n1414 240.244
R14083 gnd.n1416 gnd.n1415 240.244
R14084 gnd.n4108 gnd.n1416 240.244
R14085 gnd.n4108 gnd.n1419 240.244
R14086 gnd.n1420 gnd.n1419 240.244
R14087 gnd.n1421 gnd.n1420 240.244
R14088 gnd.n4068 gnd.n1421 240.244
R14089 gnd.n4068 gnd.n1424 240.244
R14090 gnd.n1425 gnd.n1424 240.244
R14091 gnd.n1426 gnd.n1425 240.244
R14092 gnd.n2065 gnd.n1426 240.244
R14093 gnd.n2065 gnd.n1429 240.244
R14094 gnd.n1430 gnd.n1429 240.244
R14095 gnd.n1431 gnd.n1430 240.244
R14096 gnd.n2036 gnd.n1431 240.244
R14097 gnd.n2036 gnd.n1434 240.244
R14098 gnd.n1435 gnd.n1434 240.244
R14099 gnd.n1436 gnd.n1435 240.244
R14100 gnd.n1840 gnd.n1436 240.244
R14101 gnd.n1840 gnd.n1439 240.244
R14102 gnd.n1440 gnd.n1439 240.244
R14103 gnd.n1441 gnd.n1440 240.244
R14104 gnd.n1827 gnd.n1441 240.244
R14105 gnd.n1827 gnd.n1444 240.244
R14106 gnd.n1445 gnd.n1444 240.244
R14107 gnd.n1446 gnd.n1445 240.244
R14108 gnd.n1814 gnd.n1446 240.244
R14109 gnd.n1814 gnd.n1449 240.244
R14110 gnd.n1450 gnd.n1449 240.244
R14111 gnd.n1451 gnd.n1450 240.244
R14112 gnd.n4439 gnd.n1451 240.244
R14113 gnd.n4439 gnd.n1454 240.244
R14114 gnd.n4741 gnd.n1454 240.244
R14115 gnd.n2724 gnd.n2723 240.244
R14116 gnd.n2739 gnd.n2723 240.244
R14117 gnd.n2741 gnd.n2740 240.244
R14118 gnd.n2751 gnd.n2750 240.244
R14119 gnd.n2762 gnd.n2761 240.244
R14120 gnd.n2764 gnd.n2763 240.244
R14121 gnd.n2774 gnd.n2773 240.244
R14122 gnd.n2787 gnd.n2786 240.244
R14123 gnd.n2789 gnd.n2788 240.244
R14124 gnd.n2649 gnd.n2648 240.244
R14125 gnd.n2717 gnd.n2650 240.244
R14126 gnd.n2654 gnd.n2653 240.244
R14127 gnd.n2660 gnd.n2655 240.244
R14128 gnd.n2662 gnd.n2661 240.244
R14129 gnd.n2666 gnd.n2665 240.244
R14130 gnd.n2667 gnd.n2666 240.244
R14131 gnd.n3349 gnd.n2667 240.244
R14132 gnd.n3349 gnd.n2670 240.244
R14133 gnd.n2671 gnd.n2670 240.244
R14134 gnd.n2672 gnd.n2671 240.244
R14135 gnd.n3365 gnd.n2672 240.244
R14136 gnd.n3365 gnd.n2675 240.244
R14137 gnd.n2676 gnd.n2675 240.244
R14138 gnd.n2677 gnd.n2676 240.244
R14139 gnd.n3381 gnd.n2677 240.244
R14140 gnd.n3381 gnd.n2680 240.244
R14141 gnd.n2681 gnd.n2680 240.244
R14142 gnd.n2682 gnd.n2681 240.244
R14143 gnd.n3400 gnd.n2682 240.244
R14144 gnd.n3401 gnd.n3400 240.244
R14145 gnd.n3401 gnd.n2379 240.244
R14146 gnd.n3574 gnd.n2379 240.244
R14147 gnd.n3574 gnd.n2373 240.244
R14148 gnd.n3581 gnd.n2373 240.244
R14149 gnd.n3581 gnd.n2374 240.244
R14150 gnd.n2374 gnd.n2350 240.244
R14151 gnd.n3613 gnd.n2350 240.244
R14152 gnd.n3613 gnd.n2345 240.244
R14153 gnd.n3656 gnd.n2345 240.244
R14154 gnd.n3656 gnd.n2338 240.244
R14155 gnd.n3618 gnd.n2338 240.244
R14156 gnd.n3619 gnd.n3618 240.244
R14157 gnd.n3620 gnd.n3619 240.244
R14158 gnd.n3620 gnd.n2318 240.244
R14159 gnd.n2318 gnd.n2311 240.244
R14160 gnd.n3623 gnd.n2311 240.244
R14161 gnd.n3626 gnd.n3623 240.244
R14162 gnd.n3629 gnd.n3626 240.244
R14163 gnd.n3630 gnd.n3629 240.244
R14164 gnd.n3631 gnd.n3630 240.244
R14165 gnd.n3632 gnd.n3631 240.244
R14166 gnd.n3633 gnd.n3632 240.244
R14167 gnd.n3633 gnd.n2265 240.244
R14168 gnd.n3791 gnd.n2265 240.244
R14169 gnd.n3791 gnd.n2260 240.244
R14170 gnd.n3832 gnd.n2260 240.244
R14171 gnd.n3832 gnd.n2253 240.244
R14172 gnd.n3796 gnd.n2253 240.244
R14173 gnd.n3797 gnd.n3796 240.244
R14174 gnd.n3798 gnd.n3797 240.244
R14175 gnd.n3798 gnd.n2233 240.244
R14176 gnd.n2233 gnd.n2226 240.244
R14177 gnd.n3801 gnd.n2226 240.244
R14178 gnd.n3802 gnd.n3801 240.244
R14179 gnd.n3805 gnd.n3802 240.244
R14180 gnd.n3806 gnd.n3805 240.244
R14181 gnd.n3807 gnd.n3806 240.244
R14182 gnd.n3808 gnd.n3807 240.244
R14183 gnd.n3809 gnd.n3808 240.244
R14184 gnd.n3809 gnd.n2178 240.244
R14185 gnd.n3968 gnd.n2178 240.244
R14186 gnd.n3968 gnd.n2173 240.244
R14187 gnd.n3994 gnd.n2173 240.244
R14188 gnd.n3994 gnd.n2166 240.244
R14189 gnd.n3973 gnd.n2166 240.244
R14190 gnd.n3974 gnd.n3973 240.244
R14191 gnd.n3975 gnd.n3974 240.244
R14192 gnd.n3975 gnd.n2145 240.244
R14193 gnd.n2145 gnd.n2138 240.244
R14194 gnd.n3978 gnd.n2138 240.244
R14195 gnd.n3979 gnd.n3978 240.244
R14196 gnd.n3979 gnd.n2113 240.244
R14197 gnd.n4100 gnd.n2113 240.244
R14198 gnd.n4100 gnd.n2107 240.244
R14199 gnd.n4107 gnd.n2107 240.244
R14200 gnd.n4107 gnd.n2108 240.244
R14201 gnd.n2108 gnd.n2086 240.244
R14202 gnd.n4139 gnd.n2086 240.244
R14203 gnd.n4139 gnd.n2081 240.244
R14204 gnd.n4159 gnd.n2081 240.244
R14205 gnd.n4159 gnd.n2073 240.244
R14206 gnd.n4144 gnd.n2073 240.244
R14207 gnd.n4145 gnd.n4144 240.244
R14208 gnd.n4146 gnd.n4145 240.244
R14209 gnd.n4146 gnd.n2052 240.244
R14210 gnd.n2052 gnd.n2044 240.244
R14211 gnd.n2044 gnd.n1851 240.244
R14212 gnd.n4371 gnd.n1851 240.244
R14213 gnd.n4371 gnd.n1847 240.244
R14214 gnd.n4377 gnd.n1847 240.244
R14215 gnd.n4377 gnd.n1839 240.244
R14216 gnd.n4391 gnd.n1839 240.244
R14217 gnd.n4391 gnd.n1835 240.244
R14218 gnd.n4397 gnd.n1835 240.244
R14219 gnd.n4397 gnd.n1826 240.244
R14220 gnd.n4411 gnd.n1826 240.244
R14221 gnd.n4411 gnd.n1822 240.244
R14222 gnd.n4417 gnd.n1822 240.244
R14223 gnd.n4417 gnd.n1813 240.244
R14224 gnd.n4431 gnd.n1813 240.244
R14225 gnd.n4431 gnd.n1809 240.244
R14226 gnd.n4438 gnd.n1809 240.244
R14227 gnd.n4438 gnd.n1802 240.244
R14228 gnd.n4454 gnd.n1802 240.244
R14229 gnd.n4454 gnd.n1457 240.244
R14230 gnd.n1700 gnd.n1699 240.244
R14231 gnd.n1716 gnd.n1715 240.244
R14232 gnd.n1719 gnd.n1718 240.244
R14233 gnd.n1735 gnd.n1734 240.244
R14234 gnd.n1738 gnd.n1737 240.244
R14235 gnd.n1754 gnd.n1753 240.244
R14236 gnd.n1757 gnd.n1756 240.244
R14237 gnd.n1773 gnd.n1772 240.244
R14238 gnd.n1776 gnd.n1775 240.244
R14239 gnd.n1781 gnd.n1778 240.244
R14240 gnd.n1784 gnd.n1783 240.244
R14241 gnd.n1792 gnd.n1786 240.244
R14242 gnd.n1795 gnd.n1794 240.244
R14243 gnd.n1798 gnd.n1797 240.244
R14244 gnd.n2431 gnd.n2430 240.132
R14245 gnd.n4223 gnd.n4222 240.132
R14246 gnd.n6697 gnd.n6696 225.874
R14247 gnd.n6697 gnd.n734 225.874
R14248 gnd.n6705 gnd.n734 225.874
R14249 gnd.n6706 gnd.n6705 225.874
R14250 gnd.n6707 gnd.n6706 225.874
R14251 gnd.n6707 gnd.n728 225.874
R14252 gnd.n6715 gnd.n728 225.874
R14253 gnd.n6716 gnd.n6715 225.874
R14254 gnd.n6717 gnd.n6716 225.874
R14255 gnd.n6717 gnd.n722 225.874
R14256 gnd.n6725 gnd.n722 225.874
R14257 gnd.n6726 gnd.n6725 225.874
R14258 gnd.n6727 gnd.n6726 225.874
R14259 gnd.n6727 gnd.n716 225.874
R14260 gnd.n6735 gnd.n716 225.874
R14261 gnd.n6736 gnd.n6735 225.874
R14262 gnd.n6737 gnd.n6736 225.874
R14263 gnd.n6737 gnd.n710 225.874
R14264 gnd.n6745 gnd.n710 225.874
R14265 gnd.n6746 gnd.n6745 225.874
R14266 gnd.n6747 gnd.n6746 225.874
R14267 gnd.n6747 gnd.n704 225.874
R14268 gnd.n6755 gnd.n704 225.874
R14269 gnd.n6756 gnd.n6755 225.874
R14270 gnd.n6757 gnd.n6756 225.874
R14271 gnd.n6757 gnd.n698 225.874
R14272 gnd.n6765 gnd.n698 225.874
R14273 gnd.n6766 gnd.n6765 225.874
R14274 gnd.n6767 gnd.n6766 225.874
R14275 gnd.n6767 gnd.n692 225.874
R14276 gnd.n6775 gnd.n692 225.874
R14277 gnd.n6776 gnd.n6775 225.874
R14278 gnd.n6777 gnd.n6776 225.874
R14279 gnd.n6777 gnd.n686 225.874
R14280 gnd.n6785 gnd.n686 225.874
R14281 gnd.n6786 gnd.n6785 225.874
R14282 gnd.n6787 gnd.n6786 225.874
R14283 gnd.n6787 gnd.n680 225.874
R14284 gnd.n6795 gnd.n680 225.874
R14285 gnd.n6796 gnd.n6795 225.874
R14286 gnd.n6797 gnd.n6796 225.874
R14287 gnd.n6797 gnd.n674 225.874
R14288 gnd.n6805 gnd.n674 225.874
R14289 gnd.n6806 gnd.n6805 225.874
R14290 gnd.n6807 gnd.n6806 225.874
R14291 gnd.n6807 gnd.n668 225.874
R14292 gnd.n6815 gnd.n668 225.874
R14293 gnd.n6816 gnd.n6815 225.874
R14294 gnd.n6817 gnd.n6816 225.874
R14295 gnd.n6817 gnd.n662 225.874
R14296 gnd.n6825 gnd.n662 225.874
R14297 gnd.n6826 gnd.n6825 225.874
R14298 gnd.n6827 gnd.n6826 225.874
R14299 gnd.n6827 gnd.n656 225.874
R14300 gnd.n6835 gnd.n656 225.874
R14301 gnd.n6836 gnd.n6835 225.874
R14302 gnd.n6837 gnd.n6836 225.874
R14303 gnd.n6837 gnd.n650 225.874
R14304 gnd.n6845 gnd.n650 225.874
R14305 gnd.n6846 gnd.n6845 225.874
R14306 gnd.n6847 gnd.n6846 225.874
R14307 gnd.n6847 gnd.n644 225.874
R14308 gnd.n6855 gnd.n644 225.874
R14309 gnd.n6856 gnd.n6855 225.874
R14310 gnd.n6857 gnd.n6856 225.874
R14311 gnd.n6857 gnd.n638 225.874
R14312 gnd.n6865 gnd.n638 225.874
R14313 gnd.n6866 gnd.n6865 225.874
R14314 gnd.n6867 gnd.n6866 225.874
R14315 gnd.n6867 gnd.n632 225.874
R14316 gnd.n6875 gnd.n632 225.874
R14317 gnd.n6876 gnd.n6875 225.874
R14318 gnd.n6877 gnd.n6876 225.874
R14319 gnd.n6877 gnd.n626 225.874
R14320 gnd.n6885 gnd.n626 225.874
R14321 gnd.n6886 gnd.n6885 225.874
R14322 gnd.n6887 gnd.n6886 225.874
R14323 gnd.n6887 gnd.n620 225.874
R14324 gnd.n6895 gnd.n620 225.874
R14325 gnd.n6896 gnd.n6895 225.874
R14326 gnd.n6897 gnd.n6896 225.874
R14327 gnd.n6897 gnd.n614 225.874
R14328 gnd.n6905 gnd.n614 225.874
R14329 gnd.n6906 gnd.n6905 225.874
R14330 gnd.n6907 gnd.n6906 225.874
R14331 gnd.n6907 gnd.n608 225.874
R14332 gnd.n6915 gnd.n608 225.874
R14333 gnd.n6916 gnd.n6915 225.874
R14334 gnd.n6917 gnd.n6916 225.874
R14335 gnd.n6917 gnd.n602 225.874
R14336 gnd.n6925 gnd.n602 225.874
R14337 gnd.n6926 gnd.n6925 225.874
R14338 gnd.n6927 gnd.n6926 225.874
R14339 gnd.n6927 gnd.n596 225.874
R14340 gnd.n6935 gnd.n596 225.874
R14341 gnd.n6936 gnd.n6935 225.874
R14342 gnd.n6937 gnd.n6936 225.874
R14343 gnd.n6937 gnd.n590 225.874
R14344 gnd.n6945 gnd.n590 225.874
R14345 gnd.n6946 gnd.n6945 225.874
R14346 gnd.n6947 gnd.n6946 225.874
R14347 gnd.n6947 gnd.n584 225.874
R14348 gnd.n6955 gnd.n584 225.874
R14349 gnd.n6956 gnd.n6955 225.874
R14350 gnd.n6957 gnd.n6956 225.874
R14351 gnd.n6957 gnd.n578 225.874
R14352 gnd.n6965 gnd.n578 225.874
R14353 gnd.n6966 gnd.n6965 225.874
R14354 gnd.n6967 gnd.n6966 225.874
R14355 gnd.n6967 gnd.n572 225.874
R14356 gnd.n6975 gnd.n572 225.874
R14357 gnd.n6976 gnd.n6975 225.874
R14358 gnd.n6977 gnd.n6976 225.874
R14359 gnd.n6977 gnd.n566 225.874
R14360 gnd.n6985 gnd.n566 225.874
R14361 gnd.n6986 gnd.n6985 225.874
R14362 gnd.n6987 gnd.n6986 225.874
R14363 gnd.n6987 gnd.n560 225.874
R14364 gnd.n6995 gnd.n560 225.874
R14365 gnd.n6996 gnd.n6995 225.874
R14366 gnd.n6997 gnd.n6996 225.874
R14367 gnd.n6997 gnd.n554 225.874
R14368 gnd.n7005 gnd.n554 225.874
R14369 gnd.n7006 gnd.n7005 225.874
R14370 gnd.n7007 gnd.n7006 225.874
R14371 gnd.n7007 gnd.n548 225.874
R14372 gnd.n7015 gnd.n548 225.874
R14373 gnd.n7016 gnd.n7015 225.874
R14374 gnd.n7017 gnd.n7016 225.874
R14375 gnd.n7017 gnd.n542 225.874
R14376 gnd.n7025 gnd.n542 225.874
R14377 gnd.n7026 gnd.n7025 225.874
R14378 gnd.n7027 gnd.n7026 225.874
R14379 gnd.n7027 gnd.n536 225.874
R14380 gnd.n7035 gnd.n536 225.874
R14381 gnd.n7036 gnd.n7035 225.874
R14382 gnd.n7037 gnd.n7036 225.874
R14383 gnd.n7037 gnd.n530 225.874
R14384 gnd.n7045 gnd.n530 225.874
R14385 gnd.n7046 gnd.n7045 225.874
R14386 gnd.n7047 gnd.n7046 225.874
R14387 gnd.n7047 gnd.n524 225.874
R14388 gnd.n7055 gnd.n524 225.874
R14389 gnd.n7056 gnd.n7055 225.874
R14390 gnd.n7057 gnd.n7056 225.874
R14391 gnd.n7057 gnd.n518 225.874
R14392 gnd.n7065 gnd.n518 225.874
R14393 gnd.n7066 gnd.n7065 225.874
R14394 gnd.n7067 gnd.n7066 225.874
R14395 gnd.n7067 gnd.n512 225.874
R14396 gnd.n7075 gnd.n512 225.874
R14397 gnd.n7076 gnd.n7075 225.874
R14398 gnd.n7077 gnd.n7076 225.874
R14399 gnd.n7077 gnd.n506 225.874
R14400 gnd.n7085 gnd.n506 225.874
R14401 gnd.n7086 gnd.n7085 225.874
R14402 gnd.n7087 gnd.n7086 225.874
R14403 gnd.n7087 gnd.n500 225.874
R14404 gnd.n7095 gnd.n500 225.874
R14405 gnd.n7096 gnd.n7095 225.874
R14406 gnd.n7097 gnd.n7096 225.874
R14407 gnd.n7097 gnd.n494 225.874
R14408 gnd.n7105 gnd.n494 225.874
R14409 gnd.n7106 gnd.n7105 225.874
R14410 gnd.n7107 gnd.n7106 225.874
R14411 gnd.n7107 gnd.n488 225.874
R14412 gnd.n7115 gnd.n488 225.874
R14413 gnd.n7116 gnd.n7115 225.874
R14414 gnd.n7117 gnd.n7116 225.874
R14415 gnd.n7117 gnd.n482 225.874
R14416 gnd.n7125 gnd.n482 225.874
R14417 gnd.n7126 gnd.n7125 225.874
R14418 gnd.n7127 gnd.n7126 225.874
R14419 gnd.n7127 gnd.n476 225.874
R14420 gnd.n7135 gnd.n476 225.874
R14421 gnd.n7136 gnd.n7135 225.874
R14422 gnd.n7137 gnd.n7136 225.874
R14423 gnd.n7137 gnd.n470 225.874
R14424 gnd.n7145 gnd.n470 225.874
R14425 gnd.n7146 gnd.n7145 225.874
R14426 gnd.n7147 gnd.n7146 225.874
R14427 gnd.n7147 gnd.n464 225.874
R14428 gnd.n7155 gnd.n464 225.874
R14429 gnd.n7156 gnd.n7155 225.874
R14430 gnd.n7157 gnd.n7156 225.874
R14431 gnd.n7157 gnd.n458 225.874
R14432 gnd.n7165 gnd.n458 225.874
R14433 gnd.n7166 gnd.n7165 225.874
R14434 gnd.n7167 gnd.n7166 225.874
R14435 gnd.n7167 gnd.n452 225.874
R14436 gnd.n7176 gnd.n452 225.874
R14437 gnd.n7177 gnd.n7176 225.874
R14438 gnd.n7178 gnd.n7177 225.874
R14439 gnd.n7178 gnd.n447 225.874
R14440 gnd.n5557 gnd.t233 224.174
R14441 gnd.n5187 gnd.t188 224.174
R14442 gnd.n1893 gnd.n1890 199.319
R14443 gnd.n2027 gnd.n1890 199.319
R14444 gnd.n2553 gnd.n2547 199.319
R14445 gnd.n2552 gnd.n2547 199.319
R14446 gnd.n2432 gnd.n2429 186.49
R14447 gnd.n4224 gnd.n4221 186.49
R14448 gnd.n6376 gnd.n6375 185
R14449 gnd.n6374 gnd.n6373 185
R14450 gnd.n6353 gnd.n6352 185
R14451 gnd.n6368 gnd.n6367 185
R14452 gnd.n6366 gnd.n6365 185
R14453 gnd.n6357 gnd.n6356 185
R14454 gnd.n6360 gnd.n6359 185
R14455 gnd.n6344 gnd.n6343 185
R14456 gnd.n6342 gnd.n6341 185
R14457 gnd.n6321 gnd.n6320 185
R14458 gnd.n6336 gnd.n6335 185
R14459 gnd.n6334 gnd.n6333 185
R14460 gnd.n6325 gnd.n6324 185
R14461 gnd.n6328 gnd.n6327 185
R14462 gnd.n6312 gnd.n6311 185
R14463 gnd.n6310 gnd.n6309 185
R14464 gnd.n6289 gnd.n6288 185
R14465 gnd.n6304 gnd.n6303 185
R14466 gnd.n6302 gnd.n6301 185
R14467 gnd.n6293 gnd.n6292 185
R14468 gnd.n6296 gnd.n6295 185
R14469 gnd.n6281 gnd.n6280 185
R14470 gnd.n6279 gnd.n6278 185
R14471 gnd.n6258 gnd.n6257 185
R14472 gnd.n6273 gnd.n6272 185
R14473 gnd.n6271 gnd.n6270 185
R14474 gnd.n6262 gnd.n6261 185
R14475 gnd.n6265 gnd.n6264 185
R14476 gnd.n6249 gnd.n6248 185
R14477 gnd.n6247 gnd.n6246 185
R14478 gnd.n6226 gnd.n6225 185
R14479 gnd.n6241 gnd.n6240 185
R14480 gnd.n6239 gnd.n6238 185
R14481 gnd.n6230 gnd.n6229 185
R14482 gnd.n6233 gnd.n6232 185
R14483 gnd.n6217 gnd.n6216 185
R14484 gnd.n6215 gnd.n6214 185
R14485 gnd.n6194 gnd.n6193 185
R14486 gnd.n6209 gnd.n6208 185
R14487 gnd.n6207 gnd.n6206 185
R14488 gnd.n6198 gnd.n6197 185
R14489 gnd.n6201 gnd.n6200 185
R14490 gnd.n6185 gnd.n6184 185
R14491 gnd.n6183 gnd.n6182 185
R14492 gnd.n6162 gnd.n6161 185
R14493 gnd.n6177 gnd.n6176 185
R14494 gnd.n6175 gnd.n6174 185
R14495 gnd.n6166 gnd.n6165 185
R14496 gnd.n6169 gnd.n6168 185
R14497 gnd.n6154 gnd.n6153 185
R14498 gnd.n6152 gnd.n6151 185
R14499 gnd.n6131 gnd.n6130 185
R14500 gnd.n6146 gnd.n6145 185
R14501 gnd.n6144 gnd.n6143 185
R14502 gnd.n6135 gnd.n6134 185
R14503 gnd.n6138 gnd.n6137 185
R14504 gnd.n5558 gnd.t232 178.987
R14505 gnd.n5188 gnd.t189 178.987
R14506 gnd.n1 gnd.t160 170.774
R14507 gnd.n9 gnd.t129 170.103
R14508 gnd.n8 gnd.t98 170.103
R14509 gnd.n7 gnd.t69 170.103
R14510 gnd.n6 gnd.t307 170.103
R14511 gnd.n5 gnd.t121 170.103
R14512 gnd.n4 gnd.t322 170.103
R14513 gnd.n3 gnd.t60 170.103
R14514 gnd.n2 gnd.t58 170.103
R14515 gnd.n1 gnd.t56 170.103
R14516 gnd.n4295 gnd.n4294 163.367
R14517 gnd.n4291 gnd.n4290 163.367
R14518 gnd.n4287 gnd.n4286 163.367
R14519 gnd.n4283 gnd.n4282 163.367
R14520 gnd.n4279 gnd.n4278 163.367
R14521 gnd.n4275 gnd.n4274 163.367
R14522 gnd.n4271 gnd.n4270 163.367
R14523 gnd.n4267 gnd.n4266 163.367
R14524 gnd.n4263 gnd.n4262 163.367
R14525 gnd.n4259 gnd.n4258 163.367
R14526 gnd.n4255 gnd.n4254 163.367
R14527 gnd.n4251 gnd.n4250 163.367
R14528 gnd.n4247 gnd.n4246 163.367
R14529 gnd.n4243 gnd.n4242 163.367
R14530 gnd.n4238 gnd.n4237 163.367
R14531 gnd.n4234 gnd.n4233 163.367
R14532 gnd.n4368 gnd.n4367 163.367
R14533 gnd.n4364 gnd.n4363 163.367
R14534 gnd.n4359 gnd.n4358 163.367
R14535 gnd.n4355 gnd.n4354 163.367
R14536 gnd.n4351 gnd.n4350 163.367
R14537 gnd.n4347 gnd.n4346 163.367
R14538 gnd.n4343 gnd.n4342 163.367
R14539 gnd.n4339 gnd.n4338 163.367
R14540 gnd.n4335 gnd.n4334 163.367
R14541 gnd.n4331 gnd.n4330 163.367
R14542 gnd.n4327 gnd.n4326 163.367
R14543 gnd.n4323 gnd.n4322 163.367
R14544 gnd.n4319 gnd.n4318 163.367
R14545 gnd.n4315 gnd.n4314 163.367
R14546 gnd.n4311 gnd.n4310 163.367
R14547 gnd.n4307 gnd.n4306 163.367
R14548 gnd.n2478 gnd.n2477 163.367
R14549 gnd.n2477 gnd.n2371 163.367
R14550 gnd.n2372 gnd.n2371 163.367
R14551 gnd.n2372 gnd.n2365 163.367
R14552 gnd.n2471 gnd.n2365 163.367
R14553 gnd.n2471 gnd.n2357 163.367
R14554 gnd.n2467 gnd.n2357 163.367
R14555 gnd.n2467 gnd.n2351 163.367
R14556 gnd.n2464 gnd.n2351 163.367
R14557 gnd.n2464 gnd.n2344 163.367
R14558 gnd.n2459 gnd.n2344 163.367
R14559 gnd.n2459 gnd.n2339 163.367
R14560 gnd.n2456 gnd.n2339 163.367
R14561 gnd.n2456 gnd.n2329 163.367
R14562 gnd.n2329 gnd.n2321 163.367
R14563 gnd.n3683 gnd.n2321 163.367
R14564 gnd.n3683 gnd.n2319 163.367
R14565 gnd.n3688 gnd.n2319 163.367
R14566 gnd.n3688 gnd.n2310 163.367
R14567 gnd.n2310 gnd.n2302 163.367
R14568 gnd.n3719 gnd.n2302 163.367
R14569 gnd.n3719 gnd.n2299 163.367
R14570 gnd.n3724 gnd.n2299 163.367
R14571 gnd.n3724 gnd.n2300 163.367
R14572 gnd.n2300 gnd.n2289 163.367
R14573 gnd.n3735 gnd.n2289 163.367
R14574 gnd.n3735 gnd.n2287 163.367
R14575 gnd.n3760 gnd.n2287 163.367
R14576 gnd.n3760 gnd.n2281 163.367
R14577 gnd.n3756 gnd.n2281 163.367
R14578 gnd.n3756 gnd.n2273 163.367
R14579 gnd.n3752 gnd.n2273 163.367
R14580 gnd.n3752 gnd.n2267 163.367
R14581 gnd.n3749 gnd.n2267 163.367
R14582 gnd.n3749 gnd.n2259 163.367
R14583 gnd.n3744 gnd.n2259 163.367
R14584 gnd.n3744 gnd.n2254 163.367
R14585 gnd.n3741 gnd.n2254 163.367
R14586 gnd.n3741 gnd.n2243 163.367
R14587 gnd.n2243 gnd.n2236 163.367
R14588 gnd.n3860 gnd.n2236 163.367
R14589 gnd.n3860 gnd.n2234 163.367
R14590 gnd.n3865 gnd.n2234 163.367
R14591 gnd.n3865 gnd.n2225 163.367
R14592 gnd.n2225 gnd.n2216 163.367
R14593 gnd.n3896 gnd.n2216 163.367
R14594 gnd.n3896 gnd.n2213 163.367
R14595 gnd.n3901 gnd.n2213 163.367
R14596 gnd.n3901 gnd.n2214 163.367
R14597 gnd.n2214 gnd.n2202 163.367
R14598 gnd.n3912 gnd.n2202 163.367
R14599 gnd.n3912 gnd.n2200 163.367
R14600 gnd.n3938 gnd.n2200 163.367
R14601 gnd.n3938 gnd.n2193 163.367
R14602 gnd.n3934 gnd.n2193 163.367
R14603 gnd.n3934 gnd.n2185 163.367
R14604 gnd.n3930 gnd.n2185 163.367
R14605 gnd.n3930 gnd.n2180 163.367
R14606 gnd.n3927 gnd.n2180 163.367
R14607 gnd.n3927 gnd.n2172 163.367
R14608 gnd.n3921 gnd.n2172 163.367
R14609 gnd.n3921 gnd.n2167 163.367
R14610 gnd.n3918 gnd.n2167 163.367
R14611 gnd.n3918 gnd.n2156 163.367
R14612 gnd.n2156 gnd.n2148 163.367
R14613 gnd.n4022 gnd.n2148 163.367
R14614 gnd.n4022 gnd.n2146 163.367
R14615 gnd.n4027 gnd.n2146 163.367
R14616 gnd.n4027 gnd.n2137 163.367
R14617 gnd.n2137 gnd.n2128 163.367
R14618 gnd.n4057 gnd.n2128 163.367
R14619 gnd.n4057 gnd.n2125 163.367
R14620 gnd.n4089 gnd.n2125 163.367
R14621 gnd.n4089 gnd.n2126 163.367
R14622 gnd.n4085 gnd.n2126 163.367
R14623 gnd.n4085 gnd.n4084 163.367
R14624 gnd.n4084 gnd.n2105 163.367
R14625 gnd.n2106 gnd.n2105 163.367
R14626 gnd.n2106 gnd.n2100 163.367
R14627 gnd.n4078 gnd.n2100 163.367
R14628 gnd.n4078 gnd.n2093 163.367
R14629 gnd.n4074 gnd.n2093 163.367
R14630 gnd.n4074 gnd.n2088 163.367
R14631 gnd.n4071 gnd.n2088 163.367
R14632 gnd.n4071 gnd.n2080 163.367
R14633 gnd.n4065 gnd.n2080 163.367
R14634 gnd.n4065 gnd.n2074 163.367
R14635 gnd.n4062 gnd.n2074 163.367
R14636 gnd.n4062 gnd.n2062 163.367
R14637 gnd.n2062 gnd.n2055 163.367
R14638 gnd.n4186 gnd.n2055 163.367
R14639 gnd.n4186 gnd.n2053 163.367
R14640 gnd.n4192 gnd.n2053 163.367
R14641 gnd.n4192 gnd.n2043 163.367
R14642 gnd.n2043 gnd.n2035 163.367
R14643 gnd.n4302 gnd.n2035 163.367
R14644 gnd.n2423 gnd.n2422 163.367
R14645 gnd.n3556 gnd.n2422 163.367
R14646 gnd.n3554 gnd.n3553 163.367
R14647 gnd.n3550 gnd.n3549 163.367
R14648 gnd.n3546 gnd.n3545 163.367
R14649 gnd.n3542 gnd.n3541 163.367
R14650 gnd.n3538 gnd.n3537 163.367
R14651 gnd.n3534 gnd.n3533 163.367
R14652 gnd.n3530 gnd.n3529 163.367
R14653 gnd.n3526 gnd.n3525 163.367
R14654 gnd.n3522 gnd.n3521 163.367
R14655 gnd.n3518 gnd.n3517 163.367
R14656 gnd.n3514 gnd.n3513 163.367
R14657 gnd.n3510 gnd.n3509 163.367
R14658 gnd.n3506 gnd.n3505 163.367
R14659 gnd.n3502 gnd.n3501 163.367
R14660 gnd.n3498 gnd.n3497 163.367
R14661 gnd.n2540 gnd.n2539 163.367
R14662 gnd.n2535 gnd.n2534 163.367
R14663 gnd.n2531 gnd.n2530 163.367
R14664 gnd.n2527 gnd.n2526 163.367
R14665 gnd.n2523 gnd.n2522 163.367
R14666 gnd.n2519 gnd.n2518 163.367
R14667 gnd.n2515 gnd.n2514 163.367
R14668 gnd.n2511 gnd.n2510 163.367
R14669 gnd.n2507 gnd.n2506 163.367
R14670 gnd.n2503 gnd.n2502 163.367
R14671 gnd.n2499 gnd.n2498 163.367
R14672 gnd.n2495 gnd.n2494 163.367
R14673 gnd.n2491 gnd.n2490 163.367
R14674 gnd.n2487 gnd.n2486 163.367
R14675 gnd.n2483 gnd.n2482 163.367
R14676 gnd.n2424 gnd.n2368 163.367
R14677 gnd.n3586 gnd.n2368 163.367
R14678 gnd.n3586 gnd.n2366 163.367
R14679 gnd.n3590 gnd.n2366 163.367
R14680 gnd.n3590 gnd.n2355 163.367
R14681 gnd.n3605 gnd.n2355 163.367
R14682 gnd.n3605 gnd.n2353 163.367
R14683 gnd.n3609 gnd.n2353 163.367
R14684 gnd.n3609 gnd.n2342 163.367
R14685 gnd.n3659 gnd.n2342 163.367
R14686 gnd.n3659 gnd.n2340 163.367
R14687 gnd.n3663 gnd.n2340 163.367
R14688 gnd.n3663 gnd.n2326 163.367
R14689 gnd.n3676 gnd.n2326 163.367
R14690 gnd.n3676 gnd.n2323 163.367
R14691 gnd.n3681 gnd.n2323 163.367
R14692 gnd.n3681 gnd.n2324 163.367
R14693 gnd.n2324 gnd.n2308 163.367
R14694 gnd.n3704 gnd.n2308 163.367
R14695 gnd.n3704 gnd.n2305 163.367
R14696 gnd.n3717 gnd.n2305 163.367
R14697 gnd.n3717 gnd.n2306 163.367
R14698 gnd.n2306 gnd.n2297 163.367
R14699 gnd.n3712 gnd.n2297 163.367
R14700 gnd.n3712 gnd.n3708 163.367
R14701 gnd.n3708 gnd.n2285 163.367
R14702 gnd.n3764 gnd.n2285 163.367
R14703 gnd.n3764 gnd.n2283 163.367
R14704 gnd.n3768 gnd.n2283 163.367
R14705 gnd.n3768 gnd.n2271 163.367
R14706 gnd.n3784 gnd.n2271 163.367
R14707 gnd.n3784 gnd.n2269 163.367
R14708 gnd.n3788 gnd.n2269 163.367
R14709 gnd.n3788 gnd.n2257 163.367
R14710 gnd.n3835 gnd.n2257 163.367
R14711 gnd.n3835 gnd.n2255 163.367
R14712 gnd.n3839 gnd.n2255 163.367
R14713 gnd.n3839 gnd.n2241 163.367
R14714 gnd.n3853 gnd.n2241 163.367
R14715 gnd.n3853 gnd.n2238 163.367
R14716 gnd.n3858 gnd.n2238 163.367
R14717 gnd.n3858 gnd.n2239 163.367
R14718 gnd.n2239 gnd.n2223 163.367
R14719 gnd.n3881 gnd.n2223 163.367
R14720 gnd.n3881 gnd.n2219 163.367
R14721 gnd.n3894 gnd.n2219 163.367
R14722 gnd.n3894 gnd.n2221 163.367
R14723 gnd.n2221 gnd.n2210 163.367
R14724 gnd.n3889 gnd.n2210 163.367
R14725 gnd.n3889 gnd.n3885 163.367
R14726 gnd.n3885 gnd.n2198 163.367
R14727 gnd.n3942 gnd.n2198 163.367
R14728 gnd.n3942 gnd.n2196 163.367
R14729 gnd.n3946 gnd.n2196 163.367
R14730 gnd.n3946 gnd.n2183 163.367
R14731 gnd.n3961 gnd.n2183 163.367
R14732 gnd.n3961 gnd.n2181 163.367
R14733 gnd.n3965 gnd.n2181 163.367
R14734 gnd.n3965 gnd.n2170 163.367
R14735 gnd.n3998 gnd.n2170 163.367
R14736 gnd.n3998 gnd.n2168 163.367
R14737 gnd.n4002 gnd.n2168 163.367
R14738 gnd.n4002 gnd.n2154 163.367
R14739 gnd.n4015 gnd.n2154 163.367
R14740 gnd.n4015 gnd.n2151 163.367
R14741 gnd.n4020 gnd.n2151 163.367
R14742 gnd.n4020 gnd.n2152 163.367
R14743 gnd.n2152 gnd.n2135 163.367
R14744 gnd.n4042 gnd.n2135 163.367
R14745 gnd.n4042 gnd.n2131 163.367
R14746 gnd.n4055 gnd.n2131 163.367
R14747 gnd.n4055 gnd.n2133 163.367
R14748 gnd.n2133 gnd.n2124 163.367
R14749 gnd.n4050 gnd.n2124 163.367
R14750 gnd.n4050 gnd.n4046 163.367
R14751 gnd.n4046 gnd.n2104 163.367
R14752 gnd.n4113 gnd.n2104 163.367
R14753 gnd.n4113 gnd.n2102 163.367
R14754 gnd.n4117 gnd.n2102 163.367
R14755 gnd.n4117 gnd.n2092 163.367
R14756 gnd.n4132 gnd.n2092 163.367
R14757 gnd.n4132 gnd.n2090 163.367
R14758 gnd.n4136 gnd.n2090 163.367
R14759 gnd.n4136 gnd.n2078 163.367
R14760 gnd.n4162 gnd.n2078 163.367
R14761 gnd.n4162 gnd.n2076 163.367
R14762 gnd.n4166 gnd.n2076 163.367
R14763 gnd.n4166 gnd.n2060 163.367
R14764 gnd.n4179 gnd.n2060 163.367
R14765 gnd.n4179 gnd.n2057 163.367
R14766 gnd.n4184 gnd.n2057 163.367
R14767 gnd.n4184 gnd.n2058 163.367
R14768 gnd.n2058 gnd.n2041 163.367
R14769 gnd.n4209 gnd.n2041 163.367
R14770 gnd.n4209 gnd.n2038 163.367
R14771 gnd.n4300 gnd.n2038 163.367
R14772 gnd.n7187 gnd.n7186 157.537
R14773 gnd.n7188 gnd.n7187 157.537
R14774 gnd.n7188 gnd.n441 157.537
R14775 gnd.n7196 gnd.n441 157.537
R14776 gnd.n7197 gnd.n7196 157.537
R14777 gnd.n7198 gnd.n7197 157.537
R14778 gnd.n7198 gnd.n435 157.537
R14779 gnd.n7206 gnd.n435 157.537
R14780 gnd.n7207 gnd.n7206 157.537
R14781 gnd.n7208 gnd.n7207 157.537
R14782 gnd.n7208 gnd.n429 157.537
R14783 gnd.n7216 gnd.n429 157.537
R14784 gnd.n7217 gnd.n7216 157.537
R14785 gnd.n7218 gnd.n7217 157.537
R14786 gnd.n7218 gnd.n423 157.537
R14787 gnd.n7226 gnd.n423 157.537
R14788 gnd.n7227 gnd.n7226 157.537
R14789 gnd.n7228 gnd.n7227 157.537
R14790 gnd.n7228 gnd.n417 157.537
R14791 gnd.n7236 gnd.n417 157.537
R14792 gnd.n7237 gnd.n7236 157.537
R14793 gnd.n7238 gnd.n7237 157.537
R14794 gnd.n7238 gnd.n411 157.537
R14795 gnd.n7246 gnd.n411 157.537
R14796 gnd.n7247 gnd.n7246 157.537
R14797 gnd.n7248 gnd.n7247 157.537
R14798 gnd.n7248 gnd.n405 157.537
R14799 gnd.n7256 gnd.n405 157.537
R14800 gnd.n7257 gnd.n7256 157.537
R14801 gnd.n7258 gnd.n7257 157.537
R14802 gnd.n7258 gnd.n399 157.537
R14803 gnd.n7266 gnd.n399 157.537
R14804 gnd.n7267 gnd.n7266 157.537
R14805 gnd.n7268 gnd.n7267 157.537
R14806 gnd.n7268 gnd.n393 157.537
R14807 gnd.n7276 gnd.n393 157.537
R14808 gnd.n7277 gnd.n7276 157.537
R14809 gnd.n7278 gnd.n7277 157.537
R14810 gnd.n7278 gnd.n387 157.537
R14811 gnd.n7286 gnd.n387 157.537
R14812 gnd.n7287 gnd.n7286 157.537
R14813 gnd.n7288 gnd.n7287 157.537
R14814 gnd.n7288 gnd.n381 157.537
R14815 gnd.n7296 gnd.n381 157.537
R14816 gnd.n7297 gnd.n7296 157.537
R14817 gnd.n7298 gnd.n7297 157.537
R14818 gnd.n7298 gnd.n375 157.537
R14819 gnd.n7306 gnd.n375 157.537
R14820 gnd.n7307 gnd.n7306 157.537
R14821 gnd.n7308 gnd.n7307 157.537
R14822 gnd.n7308 gnd.n369 157.537
R14823 gnd.n7316 gnd.n369 157.537
R14824 gnd.n7317 gnd.n7316 157.537
R14825 gnd.n7318 gnd.n7317 157.537
R14826 gnd.n7318 gnd.n363 157.537
R14827 gnd.n7326 gnd.n363 157.537
R14828 gnd.n7327 gnd.n7326 157.537
R14829 gnd.n7328 gnd.n7327 157.537
R14830 gnd.n7328 gnd.n357 157.537
R14831 gnd.n7336 gnd.n357 157.537
R14832 gnd.n7337 gnd.n7336 157.537
R14833 gnd.n7338 gnd.n7337 157.537
R14834 gnd.n7338 gnd.n351 157.537
R14835 gnd.n7346 gnd.n351 157.537
R14836 gnd.n7347 gnd.n7346 157.537
R14837 gnd.n7348 gnd.n7347 157.537
R14838 gnd.n7348 gnd.n345 157.537
R14839 gnd.n7356 gnd.n345 157.537
R14840 gnd.n7357 gnd.n7356 157.537
R14841 gnd.n7358 gnd.n7357 157.537
R14842 gnd.n7358 gnd.n339 157.537
R14843 gnd.n7366 gnd.n339 157.537
R14844 gnd.n7367 gnd.n7366 157.537
R14845 gnd.n7368 gnd.n7367 157.537
R14846 gnd.n7368 gnd.n333 157.537
R14847 gnd.n7376 gnd.n333 157.537
R14848 gnd.n7377 gnd.n7376 157.537
R14849 gnd.n7378 gnd.n7377 157.537
R14850 gnd.n7378 gnd.n327 157.537
R14851 gnd.n7386 gnd.n327 157.537
R14852 gnd.n7387 gnd.n7386 157.537
R14853 gnd.n7389 gnd.n7387 157.537
R14854 gnd.n7389 gnd.n7388 157.537
R14855 gnd.n4230 gnd.n4229 156.462
R14856 gnd.n6316 gnd.n6284 153.042
R14857 gnd.n6380 gnd.n6379 152.079
R14858 gnd.n6348 gnd.n6347 152.079
R14859 gnd.n6316 gnd.n6315 152.079
R14860 gnd.n2437 gnd.n2436 152
R14861 gnd.n2438 gnd.n2427 152
R14862 gnd.n2440 gnd.n2439 152
R14863 gnd.n2442 gnd.n2425 152
R14864 gnd.n2444 gnd.n2443 152
R14865 gnd.n4228 gnd.n4212 152
R14866 gnd.n4220 gnd.n4213 152
R14867 gnd.n4219 gnd.n4218 152
R14868 gnd.n4217 gnd.n4214 152
R14869 gnd.n4215 gnd.t251 150.546
R14870 gnd.t168 gnd.n6358 147.661
R14871 gnd.t164 gnd.n6326 147.661
R14872 gnd.t119 gnd.n6294 147.661
R14873 gnd.t1 gnd.n6263 147.661
R14874 gnd.t327 gnd.n6231 147.661
R14875 gnd.t3 gnd.n6199 147.661
R14876 gnd.t317 gnd.n6167 147.661
R14877 gnd.t15 gnd.n6136 147.661
R14878 gnd.n1888 gnd.n1869 143.351
R14879 gnd.n3496 gnd.n2402 143.351
R14880 gnd.n3496 gnd.n2403 143.351
R14881 gnd.n2031 gnd.n2030 136.385
R14882 gnd.n3499 gnd.n3495 136.385
R14883 gnd.n2434 gnd.t224 130.484
R14884 gnd.n2443 gnd.t217 126.766
R14885 gnd.n2441 gnd.t257 126.766
R14886 gnd.n2427 gnd.t244 126.766
R14887 gnd.n2435 gnd.t275 126.766
R14888 gnd.n4216 gnd.t237 126.766
R14889 gnd.n4218 gnd.t254 126.766
R14890 gnd.n4227 gnd.t190 126.766
R14891 gnd.n4229 gnd.t263 126.766
R14892 gnd.n6375 gnd.n6374 104.615
R14893 gnd.n6374 gnd.n6352 104.615
R14894 gnd.n6367 gnd.n6352 104.615
R14895 gnd.n6367 gnd.n6366 104.615
R14896 gnd.n6366 gnd.n6356 104.615
R14897 gnd.n6359 gnd.n6356 104.615
R14898 gnd.n6343 gnd.n6342 104.615
R14899 gnd.n6342 gnd.n6320 104.615
R14900 gnd.n6335 gnd.n6320 104.615
R14901 gnd.n6335 gnd.n6334 104.615
R14902 gnd.n6334 gnd.n6324 104.615
R14903 gnd.n6327 gnd.n6324 104.615
R14904 gnd.n6311 gnd.n6310 104.615
R14905 gnd.n6310 gnd.n6288 104.615
R14906 gnd.n6303 gnd.n6288 104.615
R14907 gnd.n6303 gnd.n6302 104.615
R14908 gnd.n6302 gnd.n6292 104.615
R14909 gnd.n6295 gnd.n6292 104.615
R14910 gnd.n6280 gnd.n6279 104.615
R14911 gnd.n6279 gnd.n6257 104.615
R14912 gnd.n6272 gnd.n6257 104.615
R14913 gnd.n6272 gnd.n6271 104.615
R14914 gnd.n6271 gnd.n6261 104.615
R14915 gnd.n6264 gnd.n6261 104.615
R14916 gnd.n6248 gnd.n6247 104.615
R14917 gnd.n6247 gnd.n6225 104.615
R14918 gnd.n6240 gnd.n6225 104.615
R14919 gnd.n6240 gnd.n6239 104.615
R14920 gnd.n6239 gnd.n6229 104.615
R14921 gnd.n6232 gnd.n6229 104.615
R14922 gnd.n6216 gnd.n6215 104.615
R14923 gnd.n6215 gnd.n6193 104.615
R14924 gnd.n6208 gnd.n6193 104.615
R14925 gnd.n6208 gnd.n6207 104.615
R14926 gnd.n6207 gnd.n6197 104.615
R14927 gnd.n6200 gnd.n6197 104.615
R14928 gnd.n6184 gnd.n6183 104.615
R14929 gnd.n6183 gnd.n6161 104.615
R14930 gnd.n6176 gnd.n6161 104.615
R14931 gnd.n6176 gnd.n6175 104.615
R14932 gnd.n6175 gnd.n6165 104.615
R14933 gnd.n6168 gnd.n6165 104.615
R14934 gnd.n6153 gnd.n6152 104.615
R14935 gnd.n6152 gnd.n6130 104.615
R14936 gnd.n6145 gnd.n6130 104.615
R14937 gnd.n6145 gnd.n6144 104.615
R14938 gnd.n6144 gnd.n6134 104.615
R14939 gnd.n6137 gnd.n6134 104.615
R14940 gnd.n5707 gnd.t281 100.632
R14941 gnd.n5161 gnd.t207 100.632
R14942 gnd.n7735 gnd.n116 99.6594
R14943 gnd.n7733 gnd.n7732 99.6594
R14944 gnd.n7728 gnd.n124 99.6594
R14945 gnd.n7726 gnd.n7725 99.6594
R14946 gnd.n7721 gnd.n131 99.6594
R14947 gnd.n7719 gnd.n7718 99.6594
R14948 gnd.n7714 gnd.n138 99.6594
R14949 gnd.n7712 gnd.n7711 99.6594
R14950 gnd.n7704 gnd.n145 99.6594
R14951 gnd.n7702 gnd.n7701 99.6594
R14952 gnd.n7697 gnd.n152 99.6594
R14953 gnd.n7695 gnd.n7694 99.6594
R14954 gnd.n7690 gnd.n159 99.6594
R14955 gnd.n7688 gnd.n7687 99.6594
R14956 gnd.n7683 gnd.n166 99.6594
R14957 gnd.n7681 gnd.n7680 99.6594
R14958 gnd.n7676 gnd.n173 99.6594
R14959 gnd.n7674 gnd.n7673 99.6594
R14960 gnd.n178 gnd.n177 99.6594
R14961 gnd.n1910 gnd.n1909 99.6594
R14962 gnd.n1918 gnd.n1917 99.6594
R14963 gnd.n1921 gnd.n1920 99.6594
R14964 gnd.n1928 gnd.n1927 99.6594
R14965 gnd.n1931 gnd.n1930 99.6594
R14966 gnd.n1939 gnd.n1938 99.6594
R14967 gnd.n1942 gnd.n1941 99.6594
R14968 gnd.n1894 gnd.n1893 99.6594
R14969 gnd.n2026 gnd.n2025 99.6594
R14970 gnd.n2019 gnd.n1952 99.6594
R14971 gnd.n2018 gnd.n2017 99.6594
R14972 gnd.n2011 gnd.n1958 99.6594
R14973 gnd.n2010 gnd.n2009 99.6594
R14974 gnd.n2003 gnd.n1964 99.6594
R14975 gnd.n2002 gnd.n2001 99.6594
R14976 gnd.n1995 gnd.n1970 99.6594
R14977 gnd.n1994 gnd.n1993 99.6594
R14978 gnd.n1985 gnd.n1976 99.6594
R14979 gnd.n2605 gnd.n2604 99.6594
R14980 gnd.n2600 gnd.n2559 99.6594
R14981 gnd.n2596 gnd.n2558 99.6594
R14982 gnd.n2592 gnd.n2557 99.6594
R14983 gnd.n2588 gnd.n2556 99.6594
R14984 gnd.n2584 gnd.n2555 99.6594
R14985 gnd.n2580 gnd.n2554 99.6594
R14986 gnd.n2552 gnd.n2551 99.6594
R14987 gnd.n3489 gnd.n3488 99.6594
R14988 gnd.n3486 gnd.n3485 99.6594
R14989 gnd.n3481 gnd.n2614 99.6594
R14990 gnd.n3479 gnd.n3478 99.6594
R14991 gnd.n3474 gnd.n2621 99.6594
R14992 gnd.n3472 gnd.n3471 99.6594
R14993 gnd.n3467 gnd.n2628 99.6594
R14994 gnd.n3465 gnd.n3464 99.6594
R14995 gnd.n3460 gnd.n2637 99.6594
R14996 gnd.n3458 gnd.n3457 99.6594
R14997 gnd.n5137 gnd.n5136 99.6594
R14998 gnd.n5131 gnd.n981 99.6594
R14999 gnd.n5128 gnd.n982 99.6594
R15000 gnd.n5124 gnd.n983 99.6594
R15001 gnd.n5120 gnd.n984 99.6594
R15002 gnd.n5116 gnd.n985 99.6594
R15003 gnd.n5112 gnd.n986 99.6594
R15004 gnd.n5108 gnd.n987 99.6594
R15005 gnd.n5104 gnd.n988 99.6594
R15006 gnd.n5099 gnd.n989 99.6594
R15007 gnd.n5095 gnd.n990 99.6594
R15008 gnd.n5091 gnd.n991 99.6594
R15009 gnd.n5087 gnd.n992 99.6594
R15010 gnd.n5083 gnd.n993 99.6594
R15011 gnd.n5079 gnd.n994 99.6594
R15012 gnd.n5075 gnd.n995 99.6594
R15013 gnd.n5071 gnd.n996 99.6594
R15014 gnd.n5067 gnd.n997 99.6594
R15015 gnd.n1052 gnd.n998 99.6594
R15016 gnd.n6489 gnd.n6488 99.6594
R15017 gnd.n6484 gnd.n5145 99.6594
R15018 gnd.n6480 gnd.n5144 99.6594
R15019 gnd.n6476 gnd.n5143 99.6594
R15020 gnd.n6472 gnd.n5142 99.6594
R15021 gnd.n6468 gnd.n5141 99.6594
R15022 gnd.n6464 gnd.n5140 99.6594
R15023 gnd.n6391 gnd.n5139 99.6594
R15024 gnd.n5740 gnd.n5739 99.6594
R15025 gnd.n5734 gnd.n5682 99.6594
R15026 gnd.n5731 gnd.n5683 99.6594
R15027 gnd.n5727 gnd.n5684 99.6594
R15028 gnd.n5723 gnd.n5685 99.6594
R15029 gnd.n5719 gnd.n5686 99.6594
R15030 gnd.n5715 gnd.n5687 99.6594
R15031 gnd.n5711 gnd.n5688 99.6594
R15032 gnd.n6454 gnd.n968 99.6594
R15033 gnd.n6450 gnd.n969 99.6594
R15034 gnd.n6446 gnd.n970 99.6594
R15035 gnd.n6442 gnd.n971 99.6594
R15036 gnd.n6438 gnd.n972 99.6594
R15037 gnd.n6434 gnd.n973 99.6594
R15038 gnd.n6430 gnd.n974 99.6594
R15039 gnd.n6426 gnd.n975 99.6594
R15040 gnd.n6422 gnd.n976 99.6594
R15041 gnd.n6418 gnd.n977 99.6594
R15042 gnd.n6414 gnd.n978 99.6594
R15043 gnd.n6410 gnd.n979 99.6594
R15044 gnd.n6406 gnd.n980 99.6594
R15045 gnd.n5612 gnd.n5522 99.6594
R15046 gnd.n5610 gnd.n5525 99.6594
R15047 gnd.n5606 gnd.n5605 99.6594
R15048 gnd.n5599 gnd.n5530 99.6594
R15049 gnd.n5598 gnd.n5597 99.6594
R15050 gnd.n5591 gnd.n5536 99.6594
R15051 gnd.n5590 gnd.n5589 99.6594
R15052 gnd.n5583 gnd.n5542 99.6594
R15053 gnd.n5582 gnd.n5581 99.6594
R15054 gnd.n5575 gnd.n5548 99.6594
R15055 gnd.n5574 gnd.n5573 99.6594
R15056 gnd.n5566 gnd.n5554 99.6594
R15057 gnd.n5565 gnd.n5564 99.6594
R15058 gnd.n7583 gnd.n7582 99.6594
R15059 gnd.n7588 gnd.n7587 99.6594
R15060 gnd.n7591 gnd.n7590 99.6594
R15061 gnd.n7596 gnd.n7595 99.6594
R15062 gnd.n7599 gnd.n7598 99.6594
R15063 gnd.n7604 gnd.n7603 99.6594
R15064 gnd.n7607 gnd.n7606 99.6594
R15065 gnd.n7612 gnd.n7611 99.6594
R15066 gnd.n7615 gnd.n103 99.6594
R15067 gnd.n1687 gnd.n1686 99.6594
R15068 gnd.n1706 gnd.n1705 99.6594
R15069 gnd.n1709 gnd.n1708 99.6594
R15070 gnd.n1725 gnd.n1724 99.6594
R15071 gnd.n1728 gnd.n1727 99.6594
R15072 gnd.n1744 gnd.n1743 99.6594
R15073 gnd.n1747 gnd.n1746 99.6594
R15074 gnd.n1763 gnd.n1762 99.6594
R15075 gnd.n1766 gnd.n1765 99.6594
R15076 gnd.n2733 gnd.n2732 99.6594
R15077 gnd.n2736 gnd.n2735 99.6594
R15078 gnd.n2746 gnd.n2745 99.6594
R15079 gnd.n2755 gnd.n2754 99.6594
R15080 gnd.n2758 gnd.n2757 99.6594
R15081 gnd.n2769 gnd.n2768 99.6594
R15082 gnd.n2778 gnd.n2777 99.6594
R15083 gnd.n2781 gnd.n2780 99.6594
R15084 gnd.n2792 gnd.n2791 99.6594
R15085 gnd.n3083 gnd.n999 99.6594
R15086 gnd.n3080 gnd.n1000 99.6594
R15087 gnd.n3076 gnd.n1001 99.6594
R15088 gnd.n3072 gnd.n1002 99.6594
R15089 gnd.n3068 gnd.n1003 99.6594
R15090 gnd.n3064 gnd.n1004 99.6594
R15091 gnd.n3060 gnd.n1005 99.6594
R15092 gnd.n3056 gnd.n1006 99.6594
R15093 gnd.n3052 gnd.n1007 99.6594
R15094 gnd.n3081 gnd.n999 99.6594
R15095 gnd.n3077 gnd.n1000 99.6594
R15096 gnd.n3073 gnd.n1001 99.6594
R15097 gnd.n3069 gnd.n1002 99.6594
R15098 gnd.n3065 gnd.n1003 99.6594
R15099 gnd.n3061 gnd.n1004 99.6594
R15100 gnd.n3057 gnd.n1005 99.6594
R15101 gnd.n3053 gnd.n1006 99.6594
R15102 gnd.n3040 gnd.n1007 99.6594
R15103 gnd.n2791 gnd.n2790 99.6594
R15104 gnd.n2780 gnd.n2779 99.6594
R15105 gnd.n2777 gnd.n2770 99.6594
R15106 gnd.n2768 gnd.n2767 99.6594
R15107 gnd.n2757 gnd.n2756 99.6594
R15108 gnd.n2754 gnd.n2747 99.6594
R15109 gnd.n2745 gnd.n2744 99.6594
R15110 gnd.n2735 gnd.n2734 99.6594
R15111 gnd.n2732 gnd.n2731 99.6594
R15112 gnd.n1686 gnd.n1682 99.6594
R15113 gnd.n1707 gnd.n1706 99.6594
R15114 gnd.n1708 gnd.n1673 99.6594
R15115 gnd.n1726 gnd.n1725 99.6594
R15116 gnd.n1727 gnd.n1664 99.6594
R15117 gnd.n1745 gnd.n1744 99.6594
R15118 gnd.n1746 gnd.n1655 99.6594
R15119 gnd.n1764 gnd.n1763 99.6594
R15120 gnd.n1765 gnd.n1644 99.6594
R15121 gnd.n7616 gnd.n7615 99.6594
R15122 gnd.n7611 gnd.n7610 99.6594
R15123 gnd.n7606 gnd.n7605 99.6594
R15124 gnd.n7603 gnd.n7602 99.6594
R15125 gnd.n7598 gnd.n7597 99.6594
R15126 gnd.n7595 gnd.n7594 99.6594
R15127 gnd.n7590 gnd.n7589 99.6594
R15128 gnd.n7587 gnd.n7586 99.6594
R15129 gnd.n7582 gnd.n7581 99.6594
R15130 gnd.n5613 gnd.n5612 99.6594
R15131 gnd.n5607 gnd.n5525 99.6594
R15132 gnd.n5605 gnd.n5604 99.6594
R15133 gnd.n5600 gnd.n5599 99.6594
R15134 gnd.n5597 gnd.n5596 99.6594
R15135 gnd.n5592 gnd.n5591 99.6594
R15136 gnd.n5589 gnd.n5588 99.6594
R15137 gnd.n5584 gnd.n5583 99.6594
R15138 gnd.n5581 gnd.n5580 99.6594
R15139 gnd.n5576 gnd.n5575 99.6594
R15140 gnd.n5573 gnd.n5572 99.6594
R15141 gnd.n5567 gnd.n5566 99.6594
R15142 gnd.n5564 gnd.n5520 99.6594
R15143 gnd.n6409 gnd.n980 99.6594
R15144 gnd.n6413 gnd.n979 99.6594
R15145 gnd.n6417 gnd.n978 99.6594
R15146 gnd.n6421 gnd.n977 99.6594
R15147 gnd.n6425 gnd.n976 99.6594
R15148 gnd.n6429 gnd.n975 99.6594
R15149 gnd.n6433 gnd.n974 99.6594
R15150 gnd.n6437 gnd.n973 99.6594
R15151 gnd.n6441 gnd.n972 99.6594
R15152 gnd.n6445 gnd.n971 99.6594
R15153 gnd.n6449 gnd.n970 99.6594
R15154 gnd.n6453 gnd.n969 99.6594
R15155 gnd.n5165 gnd.n968 99.6594
R15156 gnd.n5740 gnd.n5690 99.6594
R15157 gnd.n5732 gnd.n5682 99.6594
R15158 gnd.n5728 gnd.n5683 99.6594
R15159 gnd.n5724 gnd.n5684 99.6594
R15160 gnd.n5720 gnd.n5685 99.6594
R15161 gnd.n5716 gnd.n5686 99.6594
R15162 gnd.n5712 gnd.n5687 99.6594
R15163 gnd.n5688 gnd.n5482 99.6594
R15164 gnd.n6463 gnd.n5139 99.6594
R15165 gnd.n6467 gnd.n5140 99.6594
R15166 gnd.n6471 gnd.n5141 99.6594
R15167 gnd.n6475 gnd.n5142 99.6594
R15168 gnd.n6479 gnd.n5143 99.6594
R15169 gnd.n6483 gnd.n5144 99.6594
R15170 gnd.n5146 gnd.n5145 99.6594
R15171 gnd.n6489 gnd.n965 99.6594
R15172 gnd.n5137 gnd.n1011 99.6594
R15173 gnd.n5129 gnd.n981 99.6594
R15174 gnd.n5125 gnd.n982 99.6594
R15175 gnd.n5121 gnd.n983 99.6594
R15176 gnd.n5117 gnd.n984 99.6594
R15177 gnd.n5113 gnd.n985 99.6594
R15178 gnd.n5109 gnd.n986 99.6594
R15179 gnd.n5105 gnd.n987 99.6594
R15180 gnd.n5100 gnd.n988 99.6594
R15181 gnd.n5096 gnd.n989 99.6594
R15182 gnd.n5092 gnd.n990 99.6594
R15183 gnd.n5088 gnd.n991 99.6594
R15184 gnd.n5084 gnd.n992 99.6594
R15185 gnd.n5080 gnd.n993 99.6594
R15186 gnd.n5076 gnd.n994 99.6594
R15187 gnd.n5072 gnd.n995 99.6594
R15188 gnd.n5068 gnd.n996 99.6594
R15189 gnd.n1051 gnd.n997 99.6594
R15190 gnd.n5060 gnd.n998 99.6594
R15191 gnd.n3459 gnd.n3458 99.6594
R15192 gnd.n2637 gnd.n2629 99.6594
R15193 gnd.n3466 gnd.n3465 99.6594
R15194 gnd.n2628 gnd.n2622 99.6594
R15195 gnd.n3473 gnd.n3472 99.6594
R15196 gnd.n2621 gnd.n2615 99.6594
R15197 gnd.n3480 gnd.n3479 99.6594
R15198 gnd.n2614 gnd.n2608 99.6594
R15199 gnd.n3487 gnd.n3486 99.6594
R15200 gnd.n3490 gnd.n3489 99.6594
R15201 gnd.n2579 gnd.n2553 99.6594
R15202 gnd.n2583 gnd.n2554 99.6594
R15203 gnd.n2587 gnd.n2555 99.6594
R15204 gnd.n2591 gnd.n2556 99.6594
R15205 gnd.n2595 gnd.n2557 99.6594
R15206 gnd.n2599 gnd.n2558 99.6594
R15207 gnd.n2561 gnd.n2559 99.6594
R15208 gnd.n2605 gnd.n2560 99.6594
R15209 gnd.n1911 gnd.n1910 99.6594
R15210 gnd.n1919 gnd.n1918 99.6594
R15211 gnd.n1920 gnd.n1900 99.6594
R15212 gnd.n1929 gnd.n1928 99.6594
R15213 gnd.n1930 gnd.n1896 99.6594
R15214 gnd.n1940 gnd.n1939 99.6594
R15215 gnd.n1943 gnd.n1942 99.6594
R15216 gnd.n2028 gnd.n2027 99.6594
R15217 gnd.n2025 gnd.n2024 99.6594
R15218 gnd.n2020 gnd.n2019 99.6594
R15219 gnd.n2017 gnd.n2016 99.6594
R15220 gnd.n2012 gnd.n2011 99.6594
R15221 gnd.n2009 gnd.n2008 99.6594
R15222 gnd.n2004 gnd.n2003 99.6594
R15223 gnd.n2001 gnd.n2000 99.6594
R15224 gnd.n1996 gnd.n1995 99.6594
R15225 gnd.n1993 gnd.n1992 99.6594
R15226 gnd.n1986 gnd.n1985 99.6594
R15227 gnd.n177 gnd.n174 99.6594
R15228 gnd.n7675 gnd.n7674 99.6594
R15229 gnd.n173 gnd.n167 99.6594
R15230 gnd.n7682 gnd.n7681 99.6594
R15231 gnd.n166 gnd.n160 99.6594
R15232 gnd.n7689 gnd.n7688 99.6594
R15233 gnd.n159 gnd.n153 99.6594
R15234 gnd.n7696 gnd.n7695 99.6594
R15235 gnd.n152 gnd.n146 99.6594
R15236 gnd.n7703 gnd.n7702 99.6594
R15237 gnd.n145 gnd.n139 99.6594
R15238 gnd.n7713 gnd.n7712 99.6594
R15239 gnd.n138 gnd.n132 99.6594
R15240 gnd.n7720 gnd.n7719 99.6594
R15241 gnd.n131 gnd.n125 99.6594
R15242 gnd.n7727 gnd.n7726 99.6594
R15243 gnd.n124 gnd.n118 99.6594
R15244 gnd.n7734 gnd.n7733 99.6594
R15245 gnd.n116 gnd.n113 99.6594
R15246 gnd.n2839 gnd.n2838 99.6594
R15247 gnd.n2739 gnd.n2708 99.6594
R15248 gnd.n2741 gnd.n2709 99.6594
R15249 gnd.n2751 gnd.n2710 99.6594
R15250 gnd.n2762 gnd.n2711 99.6594
R15251 gnd.n2764 gnd.n2712 99.6594
R15252 gnd.n2774 gnd.n2713 99.6594
R15253 gnd.n2787 gnd.n2714 99.6594
R15254 gnd.n2788 gnd.n2715 99.6594
R15255 gnd.n2716 gnd.n2649 99.6594
R15256 gnd.n2718 gnd.n2717 99.6594
R15257 gnd.n2719 gnd.n2654 99.6594
R15258 gnd.n2720 gnd.n2660 99.6594
R15259 gnd.n2722 gnd.n2662 99.6594
R15260 gnd.n2839 gnd.n2724 99.6594
R15261 gnd.n2740 gnd.n2708 99.6594
R15262 gnd.n2750 gnd.n2709 99.6594
R15263 gnd.n2761 gnd.n2710 99.6594
R15264 gnd.n2763 gnd.n2711 99.6594
R15265 gnd.n2773 gnd.n2712 99.6594
R15266 gnd.n2786 gnd.n2713 99.6594
R15267 gnd.n2789 gnd.n2714 99.6594
R15268 gnd.n2715 gnd.n2648 99.6594
R15269 gnd.n2716 gnd.n2650 99.6594
R15270 gnd.n2718 gnd.n2653 99.6594
R15271 gnd.n2719 gnd.n2655 99.6594
R15272 gnd.n2720 gnd.n2661 99.6594
R15273 gnd.n2722 gnd.n2721 99.6594
R15274 gnd.n1700 gnd.n1698 99.6594
R15275 gnd.n1715 gnd.n1678 99.6594
R15276 gnd.n1719 gnd.n1717 99.6594
R15277 gnd.n1734 gnd.n1669 99.6594
R15278 gnd.n1738 gnd.n1736 99.6594
R15279 gnd.n1753 gnd.n1660 99.6594
R15280 gnd.n1757 gnd.n1755 99.6594
R15281 gnd.n1772 gnd.n1651 99.6594
R15282 gnd.n1775 gnd.n1774 99.6594
R15283 gnd.n1778 gnd.n1777 99.6594
R15284 gnd.n1783 gnd.n1782 99.6594
R15285 gnd.n1786 gnd.n1785 99.6594
R15286 gnd.n1794 gnd.n1793 99.6594
R15287 gnd.n1797 gnd.n1796 99.6594
R15288 gnd.n1796 gnd.n1795 99.6594
R15289 gnd.n1793 gnd.n1792 99.6594
R15290 gnd.n1785 gnd.n1784 99.6594
R15291 gnd.n1782 gnd.n1781 99.6594
R15292 gnd.n1777 gnd.n1776 99.6594
R15293 gnd.n1774 gnd.n1773 99.6594
R15294 gnd.n1756 gnd.n1651 99.6594
R15295 gnd.n1755 gnd.n1754 99.6594
R15296 gnd.n1737 gnd.n1660 99.6594
R15297 gnd.n1736 gnd.n1735 99.6594
R15298 gnd.n1718 gnd.n1669 99.6594
R15299 gnd.n1717 gnd.n1716 99.6594
R15300 gnd.n1699 gnd.n1678 99.6594
R15301 gnd.n1698 gnd.n1455 99.6594
R15302 gnd.n2656 gnd.t243 98.63
R15303 gnd.n7613 gnd.t270 98.63
R15304 gnd.n1645 gnd.t262 98.63
R15305 gnd.n2782 gnd.t286 98.63
R15306 gnd.n1948 gnd.t236 98.63
R15307 gnd.n1977 gnd.t223 98.63
R15308 gnd.n180 gnd.t292 98.63
R15309 gnd.n7706 gnd.t211 98.63
R15310 gnd.n1031 gnd.t196 98.63
R15311 gnd.n1053 gnd.t284 98.63
R15312 gnd.n2634 gnd.t289 98.63
R15313 gnd.n2545 gnd.t203 98.63
R15314 gnd.n3041 gnd.t229 98.63
R15315 gnd.n1789 gnd.t199 98.63
R15316 gnd.n2450 gnd.t268 96.6984
R15317 gnd.n2032 gnd.t249 96.6984
R15318 gnd.n2447 gnd.t216 96.6906
R15319 gnd.n4231 gnd.t273 96.6906
R15320 gnd.n7388 gnd.n106 94.5225
R15321 gnd.n2434 gnd.n2433 81.8399
R15322 gnd.n5708 gnd.t280 74.8376
R15323 gnd.n5162 gnd.t208 74.8376
R15324 gnd.n2451 gnd.t267 72.8438
R15325 gnd.n2033 gnd.t250 72.8438
R15326 gnd.n2435 gnd.n2428 72.8411
R15327 gnd.n2441 gnd.n2426 72.8411
R15328 gnd.n4227 gnd.n4226 72.8411
R15329 gnd.n2657 gnd.t242 72.836
R15330 gnd.n2448 gnd.t215 72.836
R15331 gnd.n4232 gnd.t274 72.836
R15332 gnd.n7614 gnd.t271 72.836
R15333 gnd.n1646 gnd.t261 72.836
R15334 gnd.n2783 gnd.t287 72.836
R15335 gnd.n1949 gnd.t235 72.836
R15336 gnd.n1978 gnd.t222 72.836
R15337 gnd.n181 gnd.t293 72.836
R15338 gnd.n7707 gnd.t212 72.836
R15339 gnd.n1032 gnd.t195 72.836
R15340 gnd.n1054 gnd.t283 72.836
R15341 gnd.n2635 gnd.t290 72.836
R15342 gnd.n2546 gnd.t204 72.836
R15343 gnd.n3042 gnd.t228 72.836
R15344 gnd.n1790 gnd.t200 72.836
R15345 gnd.n4295 gnd.n1853 71.676
R15346 gnd.n4291 gnd.n1854 71.676
R15347 gnd.n4287 gnd.n1855 71.676
R15348 gnd.n4283 gnd.n1856 71.676
R15349 gnd.n4279 gnd.n1857 71.676
R15350 gnd.n4275 gnd.n1858 71.676
R15351 gnd.n4271 gnd.n1859 71.676
R15352 gnd.n4267 gnd.n1860 71.676
R15353 gnd.n4263 gnd.n1861 71.676
R15354 gnd.n4259 gnd.n1862 71.676
R15355 gnd.n4255 gnd.n1863 71.676
R15356 gnd.n4251 gnd.n1864 71.676
R15357 gnd.n4247 gnd.n1865 71.676
R15358 gnd.n4243 gnd.n1866 71.676
R15359 gnd.n4238 gnd.n1867 71.676
R15360 gnd.n4234 gnd.n1868 71.676
R15361 gnd.n4368 gnd.n1888 71.676
R15362 gnd.n4364 gnd.n1887 71.676
R15363 gnd.n4359 gnd.n1886 71.676
R15364 gnd.n4355 gnd.n1885 71.676
R15365 gnd.n4351 gnd.n1884 71.676
R15366 gnd.n4347 gnd.n1883 71.676
R15367 gnd.n4343 gnd.n1882 71.676
R15368 gnd.n4339 gnd.n1881 71.676
R15369 gnd.n4335 gnd.n1880 71.676
R15370 gnd.n4331 gnd.n1879 71.676
R15371 gnd.n4327 gnd.n1878 71.676
R15372 gnd.n4323 gnd.n1877 71.676
R15373 gnd.n4319 gnd.n1876 71.676
R15374 gnd.n4315 gnd.n1875 71.676
R15375 gnd.n4311 gnd.n1874 71.676
R15376 gnd.n4307 gnd.n1873 71.676
R15377 gnd.n4303 gnd.n1872 71.676
R15378 gnd.n3562 gnd.n3561 71.676
R15379 gnd.n3556 gnd.n2388 71.676
R15380 gnd.n3553 gnd.n2389 71.676
R15381 gnd.n3549 gnd.n2390 71.676
R15382 gnd.n3545 gnd.n2391 71.676
R15383 gnd.n3541 gnd.n2392 71.676
R15384 gnd.n3537 gnd.n2393 71.676
R15385 gnd.n3533 gnd.n2394 71.676
R15386 gnd.n3529 gnd.n2395 71.676
R15387 gnd.n3525 gnd.n2396 71.676
R15388 gnd.n3521 gnd.n2397 71.676
R15389 gnd.n3517 gnd.n2398 71.676
R15390 gnd.n3513 gnd.n2399 71.676
R15391 gnd.n3509 gnd.n2400 71.676
R15392 gnd.n3505 gnd.n2401 71.676
R15393 gnd.n3501 gnd.n2402 71.676
R15394 gnd.n3497 gnd.n2404 71.676
R15395 gnd.n2539 gnd.n2405 71.676
R15396 gnd.n2534 gnd.n2406 71.676
R15397 gnd.n2530 gnd.n2407 71.676
R15398 gnd.n2526 gnd.n2408 71.676
R15399 gnd.n2522 gnd.n2409 71.676
R15400 gnd.n2518 gnd.n2410 71.676
R15401 gnd.n2514 gnd.n2411 71.676
R15402 gnd.n2510 gnd.n2412 71.676
R15403 gnd.n2506 gnd.n2413 71.676
R15404 gnd.n2502 gnd.n2414 71.676
R15405 gnd.n2498 gnd.n2415 71.676
R15406 gnd.n2494 gnd.n2416 71.676
R15407 gnd.n2490 gnd.n2417 71.676
R15408 gnd.n2486 gnd.n2418 71.676
R15409 gnd.n2482 gnd.n2419 71.676
R15410 gnd.n3562 gnd.n2423 71.676
R15411 gnd.n3554 gnd.n2388 71.676
R15412 gnd.n3550 gnd.n2389 71.676
R15413 gnd.n3546 gnd.n2390 71.676
R15414 gnd.n3542 gnd.n2391 71.676
R15415 gnd.n3538 gnd.n2392 71.676
R15416 gnd.n3534 gnd.n2393 71.676
R15417 gnd.n3530 gnd.n2394 71.676
R15418 gnd.n3526 gnd.n2395 71.676
R15419 gnd.n3522 gnd.n2396 71.676
R15420 gnd.n3518 gnd.n2397 71.676
R15421 gnd.n3514 gnd.n2398 71.676
R15422 gnd.n3510 gnd.n2399 71.676
R15423 gnd.n3506 gnd.n2400 71.676
R15424 gnd.n3502 gnd.n2401 71.676
R15425 gnd.n3498 gnd.n2403 71.676
R15426 gnd.n2540 gnd.n2404 71.676
R15427 gnd.n2535 gnd.n2405 71.676
R15428 gnd.n2531 gnd.n2406 71.676
R15429 gnd.n2527 gnd.n2407 71.676
R15430 gnd.n2523 gnd.n2408 71.676
R15431 gnd.n2519 gnd.n2409 71.676
R15432 gnd.n2515 gnd.n2410 71.676
R15433 gnd.n2511 gnd.n2411 71.676
R15434 gnd.n2507 gnd.n2412 71.676
R15435 gnd.n2503 gnd.n2413 71.676
R15436 gnd.n2499 gnd.n2414 71.676
R15437 gnd.n2495 gnd.n2415 71.676
R15438 gnd.n2491 gnd.n2416 71.676
R15439 gnd.n2487 gnd.n2417 71.676
R15440 gnd.n2483 gnd.n2418 71.676
R15441 gnd.n2479 gnd.n2419 71.676
R15442 gnd.n4306 gnd.n1872 71.676
R15443 gnd.n4310 gnd.n1873 71.676
R15444 gnd.n4314 gnd.n1874 71.676
R15445 gnd.n4318 gnd.n1875 71.676
R15446 gnd.n4322 gnd.n1876 71.676
R15447 gnd.n4326 gnd.n1877 71.676
R15448 gnd.n4330 gnd.n1878 71.676
R15449 gnd.n4334 gnd.n1879 71.676
R15450 gnd.n4338 gnd.n1880 71.676
R15451 gnd.n4342 gnd.n1881 71.676
R15452 gnd.n4346 gnd.n1882 71.676
R15453 gnd.n4350 gnd.n1883 71.676
R15454 gnd.n4354 gnd.n1884 71.676
R15455 gnd.n4358 gnd.n1885 71.676
R15456 gnd.n4363 gnd.n1886 71.676
R15457 gnd.n4367 gnd.n1887 71.676
R15458 gnd.n4233 gnd.n1869 71.676
R15459 gnd.n4237 gnd.n1868 71.676
R15460 gnd.n4242 gnd.n1867 71.676
R15461 gnd.n4246 gnd.n1866 71.676
R15462 gnd.n4250 gnd.n1865 71.676
R15463 gnd.n4254 gnd.n1864 71.676
R15464 gnd.n4258 gnd.n1863 71.676
R15465 gnd.n4262 gnd.n1862 71.676
R15466 gnd.n4266 gnd.n1861 71.676
R15467 gnd.n4270 gnd.n1860 71.676
R15468 gnd.n4274 gnd.n1859 71.676
R15469 gnd.n4278 gnd.n1858 71.676
R15470 gnd.n4282 gnd.n1857 71.676
R15471 gnd.n4286 gnd.n1856 71.676
R15472 gnd.n4290 gnd.n1855 71.676
R15473 gnd.n4294 gnd.n1854 71.676
R15474 gnd.n2039 gnd.n1853 71.676
R15475 gnd.n10 gnd.t324 69.1507
R15476 gnd.n18 gnd.t13 68.4792
R15477 gnd.n17 gnd.t162 68.4792
R15478 gnd.n16 gnd.t62 68.4792
R15479 gnd.n15 gnd.t34 68.4792
R15480 gnd.n14 gnd.t94 68.4792
R15481 gnd.n13 gnd.t11 68.4792
R15482 gnd.n12 gnd.t166 68.4792
R15483 gnd.n11 gnd.t92 68.4792
R15484 gnd.n10 gnd.t96 68.4792
R15485 gnd.n5620 gnd.n5521 64.369
R15486 gnd.n2537 gnd.n2451 59.5399
R15487 gnd.n4361 gnd.n2033 59.5399
R15488 gnd.n2449 gnd.n2448 59.5399
R15489 gnd.n4240 gnd.n4232 59.5399
R15490 gnd.n2446 gnd.n2444 59.1804
R15491 gnd.n6490 gnd.n966 57.3586
R15492 gnd.n5138 gnd.n1009 57.3586
R15493 gnd.n5327 gnd.t325 56.607
R15494 gnd.n52 gnd.t24 56.607
R15495 gnd.n5296 gnd.t9 56.407
R15496 gnd.n5311 gnd.t102 56.407
R15497 gnd.n21 gnd.t65 56.407
R15498 gnd.n36 gnd.t23 56.407
R15499 gnd.n5340 gnd.t111 55.8337
R15500 gnd.n5309 gnd.t42 55.8337
R15501 gnd.n5324 gnd.t319 55.8337
R15502 gnd.n65 gnd.t86 55.8337
R15503 gnd.n34 gnd.t105 55.8337
R15504 gnd.n49 gnd.t140 55.8337
R15505 gnd.n2432 gnd.n2431 54.358
R15506 gnd.n4224 gnd.n4223 54.358
R15507 gnd.n5327 gnd.n5326 53.0052
R15508 gnd.n5329 gnd.n5328 53.0052
R15509 gnd.n5331 gnd.n5330 53.0052
R15510 gnd.n5333 gnd.n5332 53.0052
R15511 gnd.n5335 gnd.n5334 53.0052
R15512 gnd.n5337 gnd.n5336 53.0052
R15513 gnd.n5339 gnd.n5338 53.0052
R15514 gnd.n5296 gnd.n5295 53.0052
R15515 gnd.n5298 gnd.n5297 53.0052
R15516 gnd.n5300 gnd.n5299 53.0052
R15517 gnd.n5302 gnd.n5301 53.0052
R15518 gnd.n5304 gnd.n5303 53.0052
R15519 gnd.n5306 gnd.n5305 53.0052
R15520 gnd.n5308 gnd.n5307 53.0052
R15521 gnd.n5311 gnd.n5310 53.0052
R15522 gnd.n5313 gnd.n5312 53.0052
R15523 gnd.n5315 gnd.n5314 53.0052
R15524 gnd.n5317 gnd.n5316 53.0052
R15525 gnd.n5319 gnd.n5318 53.0052
R15526 gnd.n5321 gnd.n5320 53.0052
R15527 gnd.n5323 gnd.n5322 53.0052
R15528 gnd.n64 gnd.n63 53.0052
R15529 gnd.n62 gnd.n61 53.0052
R15530 gnd.n60 gnd.n59 53.0052
R15531 gnd.n58 gnd.n57 53.0052
R15532 gnd.n56 gnd.n55 53.0052
R15533 gnd.n54 gnd.n53 53.0052
R15534 gnd.n52 gnd.n51 53.0052
R15535 gnd.n33 gnd.n32 53.0052
R15536 gnd.n31 gnd.n30 53.0052
R15537 gnd.n29 gnd.n28 53.0052
R15538 gnd.n27 gnd.n26 53.0052
R15539 gnd.n25 gnd.n24 53.0052
R15540 gnd.n23 gnd.n22 53.0052
R15541 gnd.n21 gnd.n20 53.0052
R15542 gnd.n48 gnd.n47 53.0052
R15543 gnd.n46 gnd.n45 53.0052
R15544 gnd.n44 gnd.n43 53.0052
R15545 gnd.n42 gnd.n41 53.0052
R15546 gnd.n40 gnd.n39 53.0052
R15547 gnd.n38 gnd.n37 53.0052
R15548 gnd.n36 gnd.n35 53.0052
R15549 gnd.n4215 gnd.n4214 52.4801
R15550 gnd.n6359 gnd.t168 52.3082
R15551 gnd.n6327 gnd.t164 52.3082
R15552 gnd.n6295 gnd.t119 52.3082
R15553 gnd.n6264 gnd.t1 52.3082
R15554 gnd.n6232 gnd.t327 52.3082
R15555 gnd.n6200 gnd.t3 52.3082
R15556 gnd.n6168 gnd.t317 52.3082
R15557 gnd.n6137 gnd.t15 52.3082
R15558 gnd.n6189 gnd.n6157 51.4173
R15559 gnd.n6253 gnd.n6252 50.455
R15560 gnd.n6221 gnd.n6220 50.455
R15561 gnd.n6189 gnd.n6188 50.455
R15562 gnd.n5558 gnd.n5557 45.1884
R15563 gnd.n5188 gnd.n5187 45.1884
R15564 gnd.n4298 gnd.n4230 44.3322
R15565 gnd.n2435 gnd.n2434 44.3189
R15566 gnd.n7743 gnd.n106 43.6564
R15567 gnd.n2658 gnd.n2657 42.4732
R15568 gnd.n1791 gnd.n1790 42.4732
R15569 gnd.n5570 gnd.n5558 42.2793
R15570 gnd.n5189 gnd.n5188 42.2793
R15571 gnd.n5710 gnd.n5708 42.2793
R15572 gnd.n6462 gnd.n5162 42.2793
R15573 gnd.n7619 gnd.n7614 42.2793
R15574 gnd.n1647 gnd.n1646 42.2793
R15575 gnd.n2784 gnd.n2783 42.2793
R15576 gnd.n1979 gnd.n1978 42.2793
R15577 gnd.n7671 gnd.n181 42.2793
R15578 gnd.n7708 gnd.n7707 42.2793
R15579 gnd.n5102 gnd.n1032 42.2793
R15580 gnd.n1055 gnd.n1054 42.2793
R15581 gnd.n2636 gnd.n2635 42.2793
R15582 gnd.n3043 gnd.n3042 42.2793
R15583 gnd.n2433 gnd.n2432 41.6274
R15584 gnd.n4225 gnd.n4224 41.6274
R15585 gnd.n2442 gnd.n2441 40.8975
R15586 gnd.n4228 gnd.n4227 40.8975
R15587 gnd.n6695 gnd.n740 38.7329
R15588 gnd.n6689 gnd.n740 38.7329
R15589 gnd.n6689 gnd.n6688 38.7329
R15590 gnd.n6688 gnd.n6687 38.7329
R15591 gnd.n6687 gnd.n747 38.7329
R15592 gnd.n6681 gnd.n747 38.7329
R15593 gnd.n6681 gnd.n6680 38.7329
R15594 gnd.n6680 gnd.n6679 38.7329
R15595 gnd.n6679 gnd.n755 38.7329
R15596 gnd.n6673 gnd.n755 38.7329
R15597 gnd.n6673 gnd.n6672 38.7329
R15598 gnd.n6672 gnd.n6671 38.7329
R15599 gnd.n6671 gnd.n763 38.7329
R15600 gnd.n6665 gnd.n763 38.7329
R15601 gnd.n6665 gnd.n6664 38.7329
R15602 gnd.n6664 gnd.n6663 38.7329
R15603 gnd.n6663 gnd.n771 38.7329
R15604 gnd.n6657 gnd.n771 38.7329
R15605 gnd.n6657 gnd.n6656 38.7329
R15606 gnd.n6656 gnd.n6655 38.7329
R15607 gnd.n6655 gnd.n779 38.7329
R15608 gnd.n6649 gnd.n779 38.7329
R15609 gnd.n6649 gnd.n6648 38.7329
R15610 gnd.n6648 gnd.n6647 38.7329
R15611 gnd.n6647 gnd.n787 38.7329
R15612 gnd.n6641 gnd.n787 38.7329
R15613 gnd.n6641 gnd.n6640 38.7329
R15614 gnd.n6640 gnd.n6639 38.7329
R15615 gnd.n6639 gnd.n795 38.7329
R15616 gnd.n6633 gnd.n795 38.7329
R15617 gnd.n6633 gnd.n6632 38.7329
R15618 gnd.n6632 gnd.n6631 38.7329
R15619 gnd.n6631 gnd.n803 38.7329
R15620 gnd.n6625 gnd.n803 38.7329
R15621 gnd.n6625 gnd.n6624 38.7329
R15622 gnd.n6624 gnd.n6623 38.7329
R15623 gnd.n6623 gnd.n811 38.7329
R15624 gnd.n6617 gnd.n811 38.7329
R15625 gnd.n6617 gnd.n6616 38.7329
R15626 gnd.n6616 gnd.n6615 38.7329
R15627 gnd.n6615 gnd.n819 38.7329
R15628 gnd.n6609 gnd.n819 38.7329
R15629 gnd.n6609 gnd.n6608 38.7329
R15630 gnd.n6608 gnd.n6607 38.7329
R15631 gnd.n6607 gnd.n827 38.7329
R15632 gnd.n6601 gnd.n827 38.7329
R15633 gnd.n6601 gnd.n6600 38.7329
R15634 gnd.n6600 gnd.n6599 38.7329
R15635 gnd.n6599 gnd.n835 38.7329
R15636 gnd.n6593 gnd.n835 38.7329
R15637 gnd.n6593 gnd.n6592 38.7329
R15638 gnd.n6592 gnd.n6591 38.7329
R15639 gnd.n6591 gnd.n843 38.7329
R15640 gnd.n6585 gnd.n843 38.7329
R15641 gnd.n6585 gnd.n6584 38.7329
R15642 gnd.n6584 gnd.n6583 38.7329
R15643 gnd.n6583 gnd.n851 38.7329
R15644 gnd.n6577 gnd.n851 38.7329
R15645 gnd.n6577 gnd.n6576 38.7329
R15646 gnd.n6576 gnd.n6575 38.7329
R15647 gnd.n6575 gnd.n859 38.7329
R15648 gnd.n6569 gnd.n859 38.7329
R15649 gnd.n6569 gnd.n6568 38.7329
R15650 gnd.n6568 gnd.n6567 38.7329
R15651 gnd.n6567 gnd.n867 38.7329
R15652 gnd.n6561 gnd.n867 38.7329
R15653 gnd.n6561 gnd.n6560 38.7329
R15654 gnd.n6560 gnd.n6559 38.7329
R15655 gnd.n6559 gnd.n875 38.7329
R15656 gnd.n6553 gnd.n875 38.7329
R15657 gnd.n6553 gnd.n6552 38.7329
R15658 gnd.n6552 gnd.n6551 38.7329
R15659 gnd.n6551 gnd.n883 38.7329
R15660 gnd.n6545 gnd.n883 38.7329
R15661 gnd.n6545 gnd.n6544 38.7329
R15662 gnd.n6544 gnd.n6543 38.7329
R15663 gnd.n6543 gnd.n891 38.7329
R15664 gnd.n6537 gnd.n891 38.7329
R15665 gnd.n6537 gnd.n6536 38.7329
R15666 gnd.n6536 gnd.n6535 38.7329
R15667 gnd.n6535 gnd.n899 38.7329
R15668 gnd.n6529 gnd.n899 38.7329
R15669 gnd.n6529 gnd.n6528 38.7329
R15670 gnd.n2030 gnd.n1949 36.9518
R15671 gnd.n3495 gnd.n2546 36.9518
R15672 gnd.n2441 gnd.n2440 35.055
R15673 gnd.n2436 gnd.n2435 35.055
R15674 gnd.n4217 gnd.n4216 35.055
R15675 gnd.n4227 gnd.n4213 35.055
R15676 gnd.n5620 gnd.n5516 31.8661
R15677 gnd.n5628 gnd.n5516 31.8661
R15678 gnd.n5636 gnd.n5510 31.8661
R15679 gnd.n5636 gnd.n5504 31.8661
R15680 gnd.n5644 gnd.n5504 31.8661
R15681 gnd.n5644 gnd.n5497 31.8661
R15682 gnd.n5652 gnd.n5497 31.8661
R15683 gnd.n5652 gnd.n5498 31.8661
R15684 gnd.n5751 gnd.n5483 31.8661
R15685 gnd.n3100 gnd.n1009 31.8661
R15686 gnd.n5051 gnd.n1063 31.8661
R15687 gnd.n5051 gnd.n1065 31.8661
R15688 gnd.n5045 gnd.n1065 31.8661
R15689 gnd.n5045 gnd.n1077 31.8661
R15690 gnd.n5039 gnd.n1088 31.8661
R15691 gnd.n5033 gnd.n1088 31.8661
R15692 gnd.n5027 gnd.n1105 31.8661
R15693 gnd.n3327 gnd.n3325 31.8661
R15694 gnd.n3327 gnd.n3326 31.8661
R15695 gnd.n3336 gnd.n3335 31.8661
R15696 gnd.n4739 gnd.n1458 31.8661
R15697 gnd.n4733 gnd.n4732 31.8661
R15698 gnd.n4732 gnd.n4731 31.8661
R15699 gnd.n7556 gnd.n218 31.8661
R15700 gnd.n7564 gnd.n208 31.8661
R15701 gnd.n7564 gnd.n211 31.8661
R15702 gnd.n7572 gnd.n193 31.8661
R15703 gnd.n7655 gnd.n193 31.8661
R15704 gnd.n7655 gnd.n186 31.8661
R15705 gnd.n7663 gnd.n186 31.8661
R15706 gnd.n7743 gnd.n104 31.8661
R15707 gnd.n4304 gnd.n2034 30.4395
R15708 gnd.n2480 gnd.n2452 30.4395
R15709 gnd.n3141 gnd.n1116 29.3168
R15710 gnd.n5021 gnd.n1119 29.3168
R15711 gnd.n5015 gnd.n1130 29.3168
R15712 gnd.n3157 gnd.n1138 29.3168
R15713 gnd.n3165 gnd.n1148 29.3168
R15714 gnd.n3173 gnd.n1158 29.3168
R15715 gnd.n4997 gnd.n1161 29.3168
R15716 gnd.n4991 gnd.n1172 29.3168
R15717 gnd.n3189 gnd.n1178 29.3168
R15718 gnd.n3198 gnd.n1188 29.3168
R15719 gnd.n3207 gnd.n1195 29.3168
R15720 gnd.n4972 gnd.n1198 29.3168
R15721 gnd.n4966 gnd.n1209 29.3168
R15722 gnd.n3223 gnd.n1216 29.3168
R15723 gnd.n3231 gnd.n1226 29.3168
R15724 gnd.n3239 gnd.n1236 29.3168
R15725 gnd.n4948 gnd.n1239 29.3168
R15726 gnd.n4942 gnd.n1250 29.3168
R15727 gnd.n3256 gnd.n1258 29.3168
R15728 gnd.n3264 gnd.n1268 29.3168
R15729 gnd.n3299 gnd.n1278 29.3168
R15730 gnd.n4924 gnd.n1281 29.3168
R15731 gnd.n4918 gnd.n1292 29.3168
R15732 gnd.n3276 gnd.n1300 29.3168
R15733 gnd.n4912 gnd.n1303 29.3168
R15734 gnd.n3285 gnd.n1311 29.3168
R15735 gnd.n3450 gnd.n1320 29.3168
R15736 gnd.n4900 gnd.n1323 29.3168
R15737 gnd.n1477 gnd.n1476 29.3168
R15738 gnd.n4725 gnd.n4724 29.3168
R15739 gnd.n4718 gnd.n1490 29.3168
R15740 gnd.n1635 gnd.n1493 29.3168
R15741 gnd.n4528 gnd.n1634 29.3168
R15742 gnd.n4520 gnd.n1616 29.3168
R15743 gnd.n4550 gnd.n1605 29.3168
R15744 gnd.n4548 gnd.n1608 29.3168
R15745 gnd.n1598 gnd.n1589 29.3168
R15746 gnd.n4589 gnd.n1578 29.3168
R15747 gnd.n4588 gnd.n1581 29.3168
R15748 gnd.n1572 gnd.n1569 29.3168
R15749 gnd.n4612 gnd.n1561 29.3168
R15750 gnd.n4678 gnd.n1528 29.3168
R15751 gnd.n4625 gnd.n1520 29.3168
R15752 gnd.n7501 gnd.n277 29.3168
R15753 gnd.n4636 gnd.n1541 29.3168
R15754 gnd.n4665 gnd.n4664 29.3168
R15755 gnd.n4659 gnd.n4648 29.3168
R15756 gnd.n7485 gnd.n294 29.3168
R15757 gnd.n7474 gnd.n296 29.3168
R15758 gnd.n7406 gnd.n264 29.3168
R15759 gnd.n7516 gnd.n255 29.3168
R15760 gnd.n7524 gnd.n247 29.3168
R15761 gnd.n7532 gnd.n239 29.3168
R15762 gnd.n7457 gnd.n241 29.3168
R15763 gnd.n7450 gnd.n233 29.3168
R15764 gnd.n7548 gnd.n225 29.3168
R15765 gnd.n2606 gnd.n1323 28.0422
R15766 gnd.n1476 gnd.n1468 28.0422
R15767 gnd.n5003 gnd.t76 27.0862
R15768 gnd.n7413 gnd.t35 27.0862
R15769 gnd.n4979 gnd.t52 26.4489
R15770 gnd.n4660 gnd.t70 26.4489
R15771 gnd.n4954 gnd.t20 25.8116
R15772 gnd.n4679 gnd.t4 25.8116
R15773 gnd.n2657 gnd.n2656 25.7944
R15774 gnd.n5708 gnd.n5707 25.7944
R15775 gnd.n5162 gnd.n5161 25.7944
R15776 gnd.n7614 gnd.n7613 25.7944
R15777 gnd.n1646 gnd.n1645 25.7944
R15778 gnd.n2783 gnd.n2782 25.7944
R15779 gnd.n1949 gnd.n1948 25.7944
R15780 gnd.n1978 gnd.n1977 25.7944
R15781 gnd.n181 gnd.n180 25.7944
R15782 gnd.n7707 gnd.n7706 25.7944
R15783 gnd.n1032 gnd.n1031 25.7944
R15784 gnd.n1054 gnd.n1053 25.7944
R15785 gnd.n2635 gnd.n2634 25.7944
R15786 gnd.n2546 gnd.n2545 25.7944
R15787 gnd.n3042 gnd.n3041 25.7944
R15788 gnd.n1790 gnd.n1789 25.7944
R15789 gnd.n1105 gnd.t106 25.1743
R15790 gnd.n2872 gnd.t48 25.1743
R15791 gnd.n4930 gnd.t39 25.1743
R15792 gnd.n4560 gnd.t88 25.1743
R15793 gnd.n4571 gnd.t31 25.1743
R15794 gnd.n7556 gnd.t6 25.1743
R15795 gnd.n5752 gnd.n5472 24.8557
R15796 gnd.n5475 gnd.n5466 24.8557
R15797 gnd.n5773 gnd.n5451 24.8557
R15798 gnd.n5792 gnd.n5791 24.8557
R15799 gnd.n5802 gnd.n5444 24.8557
R15800 gnd.n5815 gnd.n5432 24.8557
R15801 gnd.n5840 gnd.n5416 24.8557
R15802 gnd.n5839 gnd.n5418 24.8557
R15803 gnd.n5862 gnd.n5400 24.8557
R15804 gnd.n5851 gnd.n5392 24.8557
R15805 gnd.n5887 gnd.n5886 24.8557
R15806 gnd.n5897 gnd.n5385 24.8557
R15807 gnd.n5909 gnd.n5377 24.8557
R15808 gnd.n5908 gnd.n5365 24.8557
R15809 gnd.n5927 gnd.n5926 24.8557
R15810 gnd.n5948 gnd.n5346 24.8557
R15811 gnd.n5972 gnd.n5971 24.8557
R15812 gnd.n5983 gnd.n5281 24.8557
R15813 gnd.n5982 gnd.n5283 24.8557
R15814 gnd.n5994 gnd.n5274 24.8557
R15815 gnd.n6011 gnd.n6010 24.8557
R15816 gnd.n5265 gnd.n5254 24.8557
R15817 gnd.n6034 gnd.n5243 24.8557
R15818 gnd.n5245 gnd.n5244 24.8557
R15819 gnd.n6054 gnd.n5237 24.8557
R15820 gnd.n6066 gnd.n6065 24.8557
R15821 gnd.n6077 gnd.n5224 24.8557
R15822 gnd.n6090 gnd.n5214 24.8557
R15823 gnd.n6526 gnd.n909 24.8557
R15824 gnd.n6520 gnd.n6519 24.8557
R15825 gnd.n6119 gnd.n920 24.8557
R15826 gnd.n6512 gnd.n931 24.8557
R15827 gnd.n5198 gnd.n942 24.8557
R15828 gnd.n6506 gnd.n6505 24.8557
R15829 gnd.n6498 gnd.n956 24.8557
R15830 gnd.n2886 gnd.t133 24.537
R15831 gnd.n1530 gnd.t109 24.537
R15832 gnd.n2901 gnd.t50 23.8997
R15833 gnd.n3326 gnd.n2840 23.8997
R15834 gnd.n4733 gnd.n1467 23.8997
R15835 gnd.n4649 gnd.t130 23.8997
R15836 gnd.n2451 gnd.n2450 23.855
R15837 gnd.n2033 gnd.n2032 23.855
R15838 gnd.n2448 gnd.n2447 23.855
R15839 gnd.n4232 gnd.n4231 23.855
R15840 gnd.n5770 gnd.t14 23.2624
R15841 gnd.n3005 gnd.t303 23.2624
R15842 gnd.t27 gnd.n249 23.2624
R15843 gnd.n6528 gnd.n6527 23.2399
R15844 gnd.n5762 gnd.t279 22.6251
R15845 gnd.n3100 gnd.t194 22.6251
R15846 gnd.t210 gnd.n104 22.6251
R15847 gnd.t46 gnd.n1108 21.6691
R15848 gnd.n7396 gnd.t78 21.6691
R15849 gnd.n5742 gnd.t0 21.3504
R15850 gnd.t145 gnd.n907 20.7131
R15851 gnd.t147 gnd.n5255 20.0758
R15852 gnd.n2641 gnd.t202 20.0758
R15853 gnd.t221 gnd.n1480 20.0758
R15854 gnd.n2429 gnd.t277 19.8005
R15855 gnd.n2429 gnd.t226 19.8005
R15856 gnd.n2430 gnd.t259 19.8005
R15857 gnd.n2430 gnd.t246 19.8005
R15858 gnd.n4221 gnd.t192 19.8005
R15859 gnd.n4221 gnd.t265 19.8005
R15860 gnd.n4222 gnd.t239 19.8005
R15861 gnd.n4222 gnd.t256 19.8005
R15862 gnd.n2426 gnd.n2425 19.5087
R15863 gnd.n2439 gnd.n2426 19.5087
R15864 gnd.n2437 gnd.n2428 19.5087
R15865 gnd.n4226 gnd.n4220 19.5087
R15866 gnd.t151 gnd.n5290 19.4385
R15867 gnd.n3426 gnd.n3425 19.3944
R15868 gnd.n3425 gnd.n3424 19.3944
R15869 gnd.n3424 gnd.n2668 19.3944
R15870 gnd.n3420 gnd.n2668 19.3944
R15871 gnd.n3420 gnd.n3419 19.3944
R15872 gnd.n3419 gnd.n3418 19.3944
R15873 gnd.n3418 gnd.n2673 19.3944
R15874 gnd.n3414 gnd.n2673 19.3944
R15875 gnd.n3414 gnd.n3413 19.3944
R15876 gnd.n3413 gnd.n3412 19.3944
R15877 gnd.n3412 gnd.n2678 19.3944
R15878 gnd.n3408 gnd.n2678 19.3944
R15879 gnd.n3408 gnd.n3407 19.3944
R15880 gnd.n3407 gnd.n3406 19.3944
R15881 gnd.n3406 gnd.n2683 19.3944
R15882 gnd.n3402 gnd.n2683 19.3944
R15883 gnd.n3402 gnd.n2378 19.3944
R15884 gnd.n3575 gnd.n2378 19.3944
R15885 gnd.n3575 gnd.n2375 19.3944
R15886 gnd.n3580 gnd.n2375 19.3944
R15887 gnd.n3580 gnd.n2376 19.3944
R15888 gnd.n2376 gnd.n2349 19.3944
R15889 gnd.n3614 gnd.n2349 19.3944
R15890 gnd.n3614 gnd.n2346 19.3944
R15891 gnd.n3655 gnd.n2346 19.3944
R15892 gnd.n3655 gnd.n2347 19.3944
R15893 gnd.n3651 gnd.n2347 19.3944
R15894 gnd.n3651 gnd.n3650 19.3944
R15895 gnd.n3650 gnd.n3649 19.3944
R15896 gnd.n3649 gnd.n3621 19.3944
R15897 gnd.n3645 gnd.n3621 19.3944
R15898 gnd.n3645 gnd.n3644 19.3944
R15899 gnd.n3644 gnd.n3643 19.3944
R15900 gnd.n3643 gnd.n3627 19.3944
R15901 gnd.n3639 gnd.n3627 19.3944
R15902 gnd.n3639 gnd.n3638 19.3944
R15903 gnd.n3638 gnd.n3637 19.3944
R15904 gnd.n3637 gnd.n3634 19.3944
R15905 gnd.n3634 gnd.n2264 19.3944
R15906 gnd.n3792 gnd.n2264 19.3944
R15907 gnd.n3792 gnd.n2261 19.3944
R15908 gnd.n3831 gnd.n2261 19.3944
R15909 gnd.n3831 gnd.n2262 19.3944
R15910 gnd.n3827 gnd.n2262 19.3944
R15911 gnd.n3827 gnd.n3826 19.3944
R15912 gnd.n3826 gnd.n3825 19.3944
R15913 gnd.n3825 gnd.n3799 19.3944
R15914 gnd.n3821 gnd.n3799 19.3944
R15915 gnd.n3821 gnd.n3820 19.3944
R15916 gnd.n3820 gnd.n3819 19.3944
R15917 gnd.n3819 gnd.n3803 19.3944
R15918 gnd.n3815 gnd.n3803 19.3944
R15919 gnd.n3815 gnd.n3814 19.3944
R15920 gnd.n3814 gnd.n3813 19.3944
R15921 gnd.n3813 gnd.n3810 19.3944
R15922 gnd.n3810 gnd.n2177 19.3944
R15923 gnd.n3969 gnd.n2177 19.3944
R15924 gnd.n3969 gnd.n2174 19.3944
R15925 gnd.n3993 gnd.n2174 19.3944
R15926 gnd.n3993 gnd.n2175 19.3944
R15927 gnd.n3989 gnd.n2175 19.3944
R15928 gnd.n3989 gnd.n3988 19.3944
R15929 gnd.n3988 gnd.n3987 19.3944
R15930 gnd.n3987 gnd.n3976 19.3944
R15931 gnd.n3983 gnd.n3976 19.3944
R15932 gnd.n3983 gnd.n3982 19.3944
R15933 gnd.n3982 gnd.n3981 19.3944
R15934 gnd.n3981 gnd.n2112 19.3944
R15935 gnd.n4101 gnd.n2112 19.3944
R15936 gnd.n4101 gnd.n2109 19.3944
R15937 gnd.n4106 gnd.n2109 19.3944
R15938 gnd.n4106 gnd.n2110 19.3944
R15939 gnd.n2110 gnd.n2085 19.3944
R15940 gnd.n4140 gnd.n2085 19.3944
R15941 gnd.n4140 gnd.n2082 19.3944
R15942 gnd.n4158 gnd.n2082 19.3944
R15943 gnd.n4158 gnd.n2083 19.3944
R15944 gnd.n4154 gnd.n2083 19.3944
R15945 gnd.n4154 gnd.n4153 19.3944
R15946 gnd.n4153 gnd.n4152 19.3944
R15947 gnd.n4152 gnd.n4147 19.3944
R15948 gnd.n4148 gnd.n4147 19.3944
R15949 gnd.n4148 gnd.n1850 19.3944
R15950 gnd.n4372 gnd.n1850 19.3944
R15951 gnd.n4372 gnd.n1848 19.3944
R15952 gnd.n4376 gnd.n1848 19.3944
R15953 gnd.n4376 gnd.n1838 19.3944
R15954 gnd.n4392 gnd.n1838 19.3944
R15955 gnd.n4392 gnd.n1836 19.3944
R15956 gnd.n4396 gnd.n1836 19.3944
R15957 gnd.n4396 gnd.n1825 19.3944
R15958 gnd.n4412 gnd.n1825 19.3944
R15959 gnd.n4412 gnd.n1823 19.3944
R15960 gnd.n4416 gnd.n1823 19.3944
R15961 gnd.n4416 gnd.n1812 19.3944
R15962 gnd.n4432 gnd.n1812 19.3944
R15963 gnd.n4432 gnd.n1810 19.3944
R15964 gnd.n4437 gnd.n1810 19.3944
R15965 gnd.n4437 gnd.n1801 19.3944
R15966 gnd.n4455 gnd.n1801 19.3944
R15967 gnd.n4456 gnd.n4455 19.3944
R15968 gnd.n3432 gnd.n3431 19.3944
R15969 gnd.n3431 gnd.n3430 19.3944
R15970 gnd.n3430 gnd.n2663 19.3944
R15971 gnd.n2837 gnd.n2836 19.3944
R15972 gnd.n2836 gnd.n2726 19.3944
R15973 gnd.n2829 gnd.n2726 19.3944
R15974 gnd.n2829 gnd.n2828 19.3944
R15975 gnd.n2828 gnd.n2742 19.3944
R15976 gnd.n2821 gnd.n2742 19.3944
R15977 gnd.n2821 gnd.n2820 19.3944
R15978 gnd.n2820 gnd.n2752 19.3944
R15979 gnd.n2813 gnd.n2752 19.3944
R15980 gnd.n2813 gnd.n2812 19.3944
R15981 gnd.n2812 gnd.n2765 19.3944
R15982 gnd.n2805 gnd.n2765 19.3944
R15983 gnd.n2805 gnd.n2804 19.3944
R15984 gnd.n2804 gnd.n2775 19.3944
R15985 gnd.n2797 gnd.n2775 19.3944
R15986 gnd.n2797 gnd.n2796 19.3944
R15987 gnd.n2796 gnd.n2647 19.3944
R15988 gnd.n3443 gnd.n2647 19.3944
R15989 gnd.n3443 gnd.n3442 19.3944
R15990 gnd.n3442 gnd.n3441 19.3944
R15991 gnd.n3441 gnd.n2651 19.3944
R15992 gnd.n3437 gnd.n2651 19.3944
R15993 gnd.n3437 gnd.n3436 19.3944
R15994 gnd.n3436 gnd.n3435 19.3944
R15995 gnd.n5615 gnd.n5614 19.3944
R15996 gnd.n5614 gnd.n5524 19.3944
R15997 gnd.n5609 gnd.n5524 19.3944
R15998 gnd.n5609 gnd.n5608 19.3944
R15999 gnd.n5608 gnd.n5529 19.3944
R16000 gnd.n5603 gnd.n5529 19.3944
R16001 gnd.n5603 gnd.n5602 19.3944
R16002 gnd.n5602 gnd.n5601 19.3944
R16003 gnd.n5601 gnd.n5535 19.3944
R16004 gnd.n5595 gnd.n5535 19.3944
R16005 gnd.n5595 gnd.n5594 19.3944
R16006 gnd.n5594 gnd.n5593 19.3944
R16007 gnd.n5593 gnd.n5541 19.3944
R16008 gnd.n5587 gnd.n5541 19.3944
R16009 gnd.n5587 gnd.n5586 19.3944
R16010 gnd.n5586 gnd.n5585 19.3944
R16011 gnd.n5585 gnd.n5547 19.3944
R16012 gnd.n5579 gnd.n5547 19.3944
R16013 gnd.n5579 gnd.n5578 19.3944
R16014 gnd.n5578 gnd.n5577 19.3944
R16015 gnd.n5577 gnd.n5553 19.3944
R16016 gnd.n5571 gnd.n5553 19.3944
R16017 gnd.n5569 gnd.n5568 19.3944
R16018 gnd.n5568 gnd.n5563 19.3944
R16019 gnd.n5563 gnd.n5561 19.3944
R16020 gnd.n6412 gnd.n6411 19.3944
R16021 gnd.n6411 gnd.n6408 19.3944
R16022 gnd.n6408 gnd.n6407 19.3944
R16023 gnd.n6457 gnd.n6456 19.3944
R16024 gnd.n6456 gnd.n6455 19.3944
R16025 gnd.n6455 gnd.n6452 19.3944
R16026 gnd.n6452 gnd.n6451 19.3944
R16027 gnd.n6451 gnd.n6448 19.3944
R16028 gnd.n6448 gnd.n6447 19.3944
R16029 gnd.n6447 gnd.n6444 19.3944
R16030 gnd.n6444 gnd.n6443 19.3944
R16031 gnd.n6443 gnd.n6440 19.3944
R16032 gnd.n6440 gnd.n6439 19.3944
R16033 gnd.n6439 gnd.n6436 19.3944
R16034 gnd.n6436 gnd.n6435 19.3944
R16035 gnd.n6435 gnd.n6432 19.3944
R16036 gnd.n6432 gnd.n6431 19.3944
R16037 gnd.n6431 gnd.n6428 19.3944
R16038 gnd.n6428 gnd.n6427 19.3944
R16039 gnd.n6427 gnd.n6424 19.3944
R16040 gnd.n6424 gnd.n6423 19.3944
R16041 gnd.n6423 gnd.n6420 19.3944
R16042 gnd.n6420 gnd.n6419 19.3944
R16043 gnd.n6419 gnd.n6416 19.3944
R16044 gnd.n6416 gnd.n6415 19.3944
R16045 gnd.n5755 gnd.n5754 19.3944
R16046 gnd.n5756 gnd.n5755 19.3944
R16047 gnd.n5756 gnd.n5465 19.3944
R16048 gnd.n5465 gnd.n5459 19.3944
R16049 gnd.n5781 gnd.n5459 19.3944
R16050 gnd.n5782 gnd.n5781 19.3944
R16051 gnd.n5782 gnd.n5442 19.3944
R16052 gnd.n5442 gnd.n5440 19.3944
R16053 gnd.n5806 gnd.n5440 19.3944
R16054 gnd.n5809 gnd.n5806 19.3944
R16055 gnd.n5809 gnd.n5808 19.3944
R16056 gnd.n5808 gnd.n5412 19.3944
R16057 gnd.n5847 gnd.n5412 19.3944
R16058 gnd.n5847 gnd.n5410 19.3944
R16059 gnd.n5853 gnd.n5410 19.3944
R16060 gnd.n5854 gnd.n5853 19.3944
R16061 gnd.n5854 gnd.n5380 19.3944
R16062 gnd.n5904 gnd.n5380 19.3944
R16063 gnd.n5905 gnd.n5904 19.3944
R16064 gnd.n5905 gnd.n5373 19.3944
R16065 gnd.n5916 gnd.n5373 19.3944
R16066 gnd.n5917 gnd.n5916 19.3944
R16067 gnd.n5917 gnd.n5356 19.3944
R16068 gnd.n5356 gnd.n5354 19.3944
R16069 gnd.n5941 gnd.n5354 19.3944
R16070 gnd.n5942 gnd.n5941 19.3944
R16071 gnd.n5942 gnd.n5277 19.3944
R16072 gnd.n5989 gnd.n5277 19.3944
R16073 gnd.n5990 gnd.n5989 19.3944
R16074 gnd.n5990 gnd.n5270 19.3944
R16075 gnd.n6001 gnd.n5270 19.3944
R16076 gnd.n6002 gnd.n6001 19.3944
R16077 gnd.n6002 gnd.n5253 19.3944
R16078 gnd.n5253 gnd.n5250 19.3944
R16079 gnd.n6029 gnd.n5250 19.3944
R16080 gnd.n6029 gnd.n5251 19.3944
R16081 gnd.n5251 gnd.n5233 19.3944
R16082 gnd.n6062 gnd.n5233 19.3944
R16083 gnd.n6062 gnd.n6061 19.3944
R16084 gnd.n6061 gnd.n5217 19.3944
R16085 gnd.n6087 gnd.n5217 19.3944
R16086 gnd.n6087 gnd.n5209 19.3944
R16087 gnd.n6100 gnd.n5209 19.3944
R16088 gnd.n6100 gnd.n6099 19.3944
R16089 gnd.n6099 gnd.n5202 19.3944
R16090 gnd.n6122 gnd.n5202 19.3944
R16091 gnd.n6123 gnd.n6122 19.3944
R16092 gnd.n6123 gnd.n5200 19.3944
R16093 gnd.n6385 gnd.n5200 19.3944
R16094 gnd.n6387 gnd.n6385 19.3944
R16095 gnd.n6395 gnd.n6387 19.3944
R16096 gnd.n6395 gnd.n6394 19.3944
R16097 gnd.n6394 gnd.n6393 19.3944
R16098 gnd.n5738 gnd.n5737 19.3944
R16099 gnd.n5737 gnd.n5736 19.3944
R16100 gnd.n5736 gnd.n5735 19.3944
R16101 gnd.n5735 gnd.n5733 19.3944
R16102 gnd.n5733 gnd.n5730 19.3944
R16103 gnd.n5730 gnd.n5729 19.3944
R16104 gnd.n5729 gnd.n5726 19.3944
R16105 gnd.n5726 gnd.n5725 19.3944
R16106 gnd.n5725 gnd.n5722 19.3944
R16107 gnd.n5722 gnd.n5721 19.3944
R16108 gnd.n5721 gnd.n5718 19.3944
R16109 gnd.n5718 gnd.n5717 19.3944
R16110 gnd.n5717 gnd.n5714 19.3944
R16111 gnd.n5714 gnd.n5713 19.3944
R16112 gnd.n5764 gnd.n5470 19.3944
R16113 gnd.n5764 gnd.n5468 19.3944
R16114 gnd.n5768 gnd.n5468 19.3944
R16115 gnd.n5768 gnd.n5449 19.3944
R16116 gnd.n5794 gnd.n5449 19.3944
R16117 gnd.n5794 gnd.n5447 19.3944
R16118 gnd.n5800 gnd.n5447 19.3944
R16119 gnd.n5800 gnd.n5799 19.3944
R16120 gnd.n5799 gnd.n5423 19.3944
R16121 gnd.n5828 gnd.n5423 19.3944
R16122 gnd.n5828 gnd.n5421 19.3944
R16123 gnd.n5837 gnd.n5421 19.3944
R16124 gnd.n5837 gnd.n5836 19.3944
R16125 gnd.n5836 gnd.n5835 19.3944
R16126 gnd.n5835 gnd.n5390 19.3944
R16127 gnd.n5889 gnd.n5390 19.3944
R16128 gnd.n5889 gnd.n5388 19.3944
R16129 gnd.n5895 gnd.n5388 19.3944
R16130 gnd.n5895 gnd.n5894 19.3944
R16131 gnd.n5894 gnd.n5363 19.3944
R16132 gnd.n5929 gnd.n5363 19.3944
R16133 gnd.n5929 gnd.n5361 19.3944
R16134 gnd.n5935 gnd.n5361 19.3944
R16135 gnd.n5935 gnd.n5934 19.3944
R16136 gnd.n5934 gnd.n5288 19.3944
R16137 gnd.n5974 gnd.n5288 19.3944
R16138 gnd.n5974 gnd.n5286 19.3944
R16139 gnd.n5980 gnd.n5286 19.3944
R16140 gnd.n5980 gnd.n5979 19.3944
R16141 gnd.n5979 gnd.n5260 19.3944
R16142 gnd.n6013 gnd.n5260 19.3944
R16143 gnd.n6013 gnd.n5258 19.3944
R16144 gnd.n6022 gnd.n5258 19.3944
R16145 gnd.n6022 gnd.n6021 19.3944
R16146 gnd.n6021 gnd.n6020 19.3944
R16147 gnd.n6020 gnd.n5229 19.3944
R16148 gnd.n6068 gnd.n5229 19.3944
R16149 gnd.n6068 gnd.n5227 19.3944
R16150 gnd.n6075 gnd.n5227 19.3944
R16151 gnd.n6075 gnd.n6074 19.3944
R16152 gnd.n6074 gnd.n912 19.3944
R16153 gnd.n6524 gnd.n912 19.3944
R16154 gnd.n6524 gnd.n6523 19.3944
R16155 gnd.n6523 gnd.n6522 19.3944
R16156 gnd.n6522 gnd.n916 19.3944
R16157 gnd.n934 gnd.n916 19.3944
R16158 gnd.n6510 gnd.n934 19.3944
R16159 gnd.n6510 gnd.n6509 19.3944
R16160 gnd.n6509 gnd.n6508 19.3944
R16161 gnd.n6508 gnd.n940 19.3944
R16162 gnd.n959 gnd.n940 19.3944
R16163 gnd.n6496 gnd.n959 19.3944
R16164 gnd.n6496 gnd.n6495 19.3944
R16165 gnd.n6492 gnd.n964 19.3944
R16166 gnd.n6487 gnd.n964 19.3944
R16167 gnd.n6487 gnd.n6486 19.3944
R16168 gnd.n6486 gnd.n6485 19.3944
R16169 gnd.n6485 gnd.n6482 19.3944
R16170 gnd.n6482 gnd.n6481 19.3944
R16171 gnd.n6481 gnd.n6478 19.3944
R16172 gnd.n6478 gnd.n6477 19.3944
R16173 gnd.n6477 gnd.n6474 19.3944
R16174 gnd.n6474 gnd.n6473 19.3944
R16175 gnd.n6473 gnd.n6470 19.3944
R16176 gnd.n6470 gnd.n6469 19.3944
R16177 gnd.n6469 gnd.n6466 19.3944
R16178 gnd.n6466 gnd.n6465 19.3944
R16179 gnd.n5622 gnd.n5518 19.3944
R16180 gnd.n5626 gnd.n5518 19.3944
R16181 gnd.n5626 gnd.n5508 19.3944
R16182 gnd.n5638 gnd.n5508 19.3944
R16183 gnd.n5638 gnd.n5506 19.3944
R16184 gnd.n5642 gnd.n5506 19.3944
R16185 gnd.n5642 gnd.n5495 19.3944
R16186 gnd.n5654 gnd.n5495 19.3944
R16187 gnd.n5654 gnd.n5493 19.3944
R16188 gnd.n5680 gnd.n5493 19.3944
R16189 gnd.n5680 gnd.n5679 19.3944
R16190 gnd.n5679 gnd.n5678 19.3944
R16191 gnd.n5678 gnd.n5677 19.3944
R16192 gnd.n5677 gnd.n5675 19.3944
R16193 gnd.n5675 gnd.n5674 19.3944
R16194 gnd.n5674 gnd.n5672 19.3944
R16195 gnd.n5672 gnd.n5671 19.3944
R16196 gnd.n5671 gnd.n5669 19.3944
R16197 gnd.n5669 gnd.n5668 19.3944
R16198 gnd.n5668 gnd.n5430 19.3944
R16199 gnd.n5817 gnd.n5430 19.3944
R16200 gnd.n5817 gnd.n5428 19.3944
R16201 gnd.n5823 gnd.n5428 19.3944
R16202 gnd.n5823 gnd.n5822 19.3944
R16203 gnd.n5822 gnd.n5397 19.3944
R16204 gnd.n5864 gnd.n5397 19.3944
R16205 gnd.n5864 gnd.n5395 19.3944
R16206 gnd.n5868 gnd.n5395 19.3944
R16207 gnd.n5882 gnd.n5868 19.3944
R16208 gnd.n5880 gnd.n5879 19.3944
R16209 gnd.n5876 gnd.n5875 19.3944
R16210 gnd.n5872 gnd.n5871 19.3944
R16211 gnd.n5950 gnd.n5344 19.3944
R16212 gnd.n5950 gnd.n5294 19.3944
R16213 gnd.n5969 gnd.n5294 19.3944
R16214 gnd.n5969 gnd.n5968 19.3944
R16215 gnd.n5968 gnd.n5967 19.3944
R16216 gnd.n5967 gnd.n5965 19.3944
R16217 gnd.n5965 gnd.n5964 19.3944
R16218 gnd.n5964 gnd.n5962 19.3944
R16219 gnd.n5962 gnd.n5961 19.3944
R16220 gnd.n5961 gnd.n5241 19.3944
R16221 gnd.n6036 gnd.n5241 19.3944
R16222 gnd.n6036 gnd.n5239 19.3944
R16223 gnd.n6052 gnd.n5239 19.3944
R16224 gnd.n6052 gnd.n6051 19.3944
R16225 gnd.n6051 gnd.n6050 19.3944
R16226 gnd.n6050 gnd.n6049 19.3944
R16227 gnd.n6049 gnd.n6047 19.3944
R16228 gnd.n6047 gnd.n6046 19.3944
R16229 gnd.n6046 gnd.n5207 19.3944
R16230 gnd.n6105 gnd.n5207 19.3944
R16231 gnd.n6105 gnd.n5205 19.3944
R16232 gnd.n6117 gnd.n5205 19.3944
R16233 gnd.n6117 gnd.n6116 19.3944
R16234 gnd.n6116 gnd.n6115 19.3944
R16235 gnd.n6115 gnd.n6112 19.3944
R16236 gnd.n6112 gnd.n5196 19.3944
R16237 gnd.n6400 gnd.n5196 19.3944
R16238 gnd.n6400 gnd.n5194 19.3944
R16239 gnd.n6404 gnd.n5194 19.3944
R16240 gnd.n5618 gnd.n5514 19.3944
R16241 gnd.n5630 gnd.n5514 19.3944
R16242 gnd.n5630 gnd.n5512 19.3944
R16243 gnd.n5634 gnd.n5512 19.3944
R16244 gnd.n5634 gnd.n5502 19.3944
R16245 gnd.n5646 gnd.n5502 19.3944
R16246 gnd.n5646 gnd.n5500 19.3944
R16247 gnd.n5650 gnd.n5500 19.3944
R16248 gnd.n5650 gnd.n5489 19.3944
R16249 gnd.n5744 gnd.n5489 19.3944
R16250 gnd.n5744 gnd.n5486 19.3944
R16251 gnd.n5749 gnd.n5486 19.3944
R16252 gnd.n5749 gnd.n5477 19.3944
R16253 gnd.n5759 gnd.n5477 19.3944
R16254 gnd.n5759 gnd.n5461 19.3944
R16255 gnd.n5776 gnd.n5461 19.3944
R16256 gnd.n5776 gnd.n5457 19.3944
R16257 gnd.n5789 gnd.n5457 19.3944
R16258 gnd.n5789 gnd.n5788 19.3944
R16259 gnd.n5788 gnd.n5436 19.3944
R16260 gnd.n5813 gnd.n5436 19.3944
R16261 gnd.n5813 gnd.n5812 19.3944
R16262 gnd.n5812 gnd.n5414 19.3944
R16263 gnd.n5842 gnd.n5414 19.3944
R16264 gnd.n5842 gnd.n5404 19.3944
R16265 gnd.n5860 gnd.n5404 19.3944
R16266 gnd.n5860 gnd.n5859 19.3944
R16267 gnd.n5859 gnd.n5858 19.3944
R16268 gnd.n5858 gnd.n5382 19.3944
R16269 gnd.n5900 gnd.n5382 19.3944
R16270 gnd.n5900 gnd.n5375 19.3944
R16271 gnd.n5911 gnd.n5375 19.3944
R16272 gnd.n5911 gnd.n5371 19.3944
R16273 gnd.n5924 gnd.n5371 19.3944
R16274 gnd.n5924 gnd.n5923 19.3944
R16275 gnd.n5923 gnd.n5350 19.3944
R16276 gnd.n5946 gnd.n5350 19.3944
R16277 gnd.n5946 gnd.n5945 19.3944
R16278 gnd.n5945 gnd.n5279 19.3944
R16279 gnd.n5985 gnd.n5279 19.3944
R16280 gnd.n5985 gnd.n5272 19.3944
R16281 gnd.n5996 gnd.n5272 19.3944
R16282 gnd.n5996 gnd.n5268 19.3944
R16283 gnd.n6008 gnd.n5268 19.3944
R16284 gnd.n6008 gnd.n6007 19.3944
R16285 gnd.n6007 gnd.n5247 19.3944
R16286 gnd.n6032 gnd.n5247 19.3944
R16287 gnd.n6032 gnd.n5235 19.3944
R16288 gnd.n6056 gnd.n5235 19.3944
R16289 gnd.n6056 gnd.n5219 19.3944
R16290 gnd.n6080 gnd.n5219 19.3944
R16291 gnd.n6081 gnd.n6080 19.3944
R16292 gnd.n6081 gnd.n5213 19.3944
R16293 gnd.n5213 gnd.n5211 19.3944
R16294 gnd.n6094 gnd.n5211 19.3944
R16295 gnd.n6094 gnd.n923 19.3944
R16296 gnd.n6517 gnd.n923 19.3944
R16297 gnd.n6517 gnd.n6516 19.3944
R16298 gnd.n6516 gnd.n6515 19.3944
R16299 gnd.n6515 gnd.n927 19.3944
R16300 gnd.n948 gnd.n927 19.3944
R16301 gnd.n6503 gnd.n948 19.3944
R16302 gnd.n6503 gnd.n6502 19.3944
R16303 gnd.n6502 gnd.n6501 19.3944
R16304 gnd.n6501 gnd.n952 19.3944
R16305 gnd.n4480 gnd.n1641 19.3944
R16306 gnd.n4485 gnd.n1641 19.3944
R16307 gnd.n4485 gnd.n1642 19.3944
R16308 gnd.n1642 gnd.n1622 19.3944
R16309 gnd.n4530 gnd.n1622 19.3944
R16310 gnd.n4530 gnd.n1619 19.3944
R16311 gnd.n4535 gnd.n1619 19.3944
R16312 gnd.n4535 gnd.n1620 19.3944
R16313 gnd.n1620 gnd.n1595 19.3944
R16314 gnd.n4562 gnd.n1595 19.3944
R16315 gnd.n4562 gnd.n1592 19.3944
R16316 gnd.n4567 gnd.n1592 19.3944
R16317 gnd.n4567 gnd.n1593 19.3944
R16318 gnd.n1593 gnd.n1566 19.3944
R16319 gnd.n4601 gnd.n1566 19.3944
R16320 gnd.n4601 gnd.n1563 19.3944
R16321 gnd.n4609 gnd.n1563 19.3944
R16322 gnd.n4609 gnd.n1564 19.3944
R16323 gnd.n4605 gnd.n1564 19.3944
R16324 gnd.n4605 gnd.n1555 19.3944
R16325 gnd.n4627 gnd.n1555 19.3944
R16326 gnd.n4627 gnd.n1552 19.3944
R16327 gnd.n4634 gnd.n1552 19.3944
R16328 gnd.n4634 gnd.n1553 19.3944
R16329 gnd.n4630 gnd.n1553 19.3944
R16330 gnd.n4630 gnd.n69 19.3944
R16331 gnd.n7783 gnd.n69 19.3944
R16332 gnd.n7783 gnd.n7782 19.3944
R16333 gnd.n7782 gnd.n7781 19.3944
R16334 gnd.n7781 gnd.n73 19.3944
R16335 gnd.n7777 gnd.n73 19.3944
R16336 gnd.n7777 gnd.n7776 19.3944
R16337 gnd.n7776 gnd.n7775 19.3944
R16338 gnd.n7775 gnd.n78 19.3944
R16339 gnd.n7771 gnd.n78 19.3944
R16340 gnd.n7771 gnd.n7770 19.3944
R16341 gnd.n7770 gnd.n7769 19.3944
R16342 gnd.n7769 gnd.n83 19.3944
R16343 gnd.n7765 gnd.n83 19.3944
R16344 gnd.n7765 gnd.n7764 19.3944
R16345 gnd.n7764 gnd.n7763 19.3944
R16346 gnd.n7763 gnd.n88 19.3944
R16347 gnd.n7759 gnd.n88 19.3944
R16348 gnd.n7759 gnd.n7758 19.3944
R16349 gnd.n7758 gnd.n7757 19.3944
R16350 gnd.n7757 gnd.n93 19.3944
R16351 gnd.n7753 gnd.n93 19.3944
R16352 gnd.n7753 gnd.n7752 19.3944
R16353 gnd.n7752 gnd.n7751 19.3944
R16354 gnd.n7751 gnd.n98 19.3944
R16355 gnd.n7747 gnd.n98 19.3944
R16356 gnd.n7747 gnd.n7746 19.3944
R16357 gnd.n7746 gnd.n7745 19.3944
R16358 gnd.n7644 gnd.n7643 19.3944
R16359 gnd.n7643 gnd.n7642 19.3944
R16360 gnd.n7642 gnd.n7584 19.3944
R16361 gnd.n7638 gnd.n7584 19.3944
R16362 gnd.n7638 gnd.n7637 19.3944
R16363 gnd.n7637 gnd.n7636 19.3944
R16364 gnd.n7636 gnd.n7592 19.3944
R16365 gnd.n7632 gnd.n7592 19.3944
R16366 gnd.n7632 gnd.n7631 19.3944
R16367 gnd.n7631 gnd.n7630 19.3944
R16368 gnd.n7630 gnd.n7600 19.3944
R16369 gnd.n7626 gnd.n7600 19.3944
R16370 gnd.n7626 gnd.n7625 19.3944
R16371 gnd.n7625 gnd.n7624 19.3944
R16372 gnd.n7624 gnd.n7608 19.3944
R16373 gnd.n7620 gnd.n7608 19.3944
R16374 gnd.n1684 gnd.n1683 19.3944
R16375 gnd.n1704 gnd.n1683 19.3944
R16376 gnd.n1704 gnd.n1681 19.3944
R16377 gnd.n1710 gnd.n1681 19.3944
R16378 gnd.n1710 gnd.n1674 19.3944
R16379 gnd.n1723 gnd.n1674 19.3944
R16380 gnd.n1723 gnd.n1672 19.3944
R16381 gnd.n1729 gnd.n1672 19.3944
R16382 gnd.n1729 gnd.n1665 19.3944
R16383 gnd.n1742 gnd.n1665 19.3944
R16384 gnd.n1742 gnd.n1663 19.3944
R16385 gnd.n1748 gnd.n1663 19.3944
R16386 gnd.n1748 gnd.n1656 19.3944
R16387 gnd.n1761 gnd.n1656 19.3944
R16388 gnd.n1761 gnd.n1654 19.3944
R16389 gnd.n1767 gnd.n1654 19.3944
R16390 gnd.n1690 gnd.n1689 19.3944
R16391 gnd.n1689 gnd.n1496 19.3944
R16392 gnd.n4716 gnd.n1496 19.3944
R16393 gnd.n4716 gnd.n1497 19.3944
R16394 gnd.n4712 gnd.n1497 19.3944
R16395 gnd.n4712 gnd.n4711 19.3944
R16396 gnd.n4711 gnd.n4710 19.3944
R16397 gnd.n4710 gnd.n1503 19.3944
R16398 gnd.n4706 gnd.n1503 19.3944
R16399 gnd.n4706 gnd.n4705 19.3944
R16400 gnd.n4705 gnd.n4704 19.3944
R16401 gnd.n4704 gnd.n1508 19.3944
R16402 gnd.n4700 gnd.n1508 19.3944
R16403 gnd.n4700 gnd.n4699 19.3944
R16404 gnd.n4699 gnd.n4698 19.3944
R16405 gnd.n4698 gnd.n1513 19.3944
R16406 gnd.n4694 gnd.n1513 19.3944
R16407 gnd.n4694 gnd.n4693 19.3944
R16408 gnd.n4693 gnd.n4692 19.3944
R16409 gnd.n4692 gnd.n4689 19.3944
R16410 gnd.n4689 gnd.n283 19.3944
R16411 gnd.n7499 gnd.n283 19.3944
R16412 gnd.n7499 gnd.n284 19.3944
R16413 gnd.n7495 gnd.n284 19.3944
R16414 gnd.n7495 gnd.n7494 19.3944
R16415 gnd.n7494 gnd.n7493 19.3944
R16416 gnd.n7493 gnd.n290 19.3944
R16417 gnd.n7488 gnd.n290 19.3944
R16418 gnd.n7488 gnd.n7487 19.3944
R16419 gnd.n7487 gnd.n261 19.3944
R16420 gnd.n7510 gnd.n261 19.3944
R16421 gnd.n7510 gnd.n259 19.3944
R16422 gnd.n7514 gnd.n259 19.3944
R16423 gnd.n7514 gnd.n245 19.3944
R16424 gnd.n7526 gnd.n245 19.3944
R16425 gnd.n7526 gnd.n243 19.3944
R16426 gnd.n7530 gnd.n243 19.3944
R16427 gnd.n7530 gnd.n230 19.3944
R16428 gnd.n7542 gnd.n230 19.3944
R16429 gnd.n7542 gnd.n228 19.3944
R16430 gnd.n7546 gnd.n228 19.3944
R16431 gnd.n7546 gnd.n215 19.3944
R16432 gnd.n7558 gnd.n215 19.3944
R16433 gnd.n7558 gnd.n213 19.3944
R16434 gnd.n7562 gnd.n213 19.3944
R16435 gnd.n7562 gnd.n200 19.3944
R16436 gnd.n7574 gnd.n200 19.3944
R16437 gnd.n7574 gnd.n197 19.3944
R16438 gnd.n7653 gnd.n197 19.3944
R16439 gnd.n7653 gnd.n198 19.3944
R16440 gnd.n7649 gnd.n198 19.3944
R16441 gnd.n7649 gnd.n7648 19.3944
R16442 gnd.n7648 gnd.n7647 19.3944
R16443 gnd.n2730 gnd.n1326 19.3944
R16444 gnd.n2730 gnd.n2729 19.3944
R16445 gnd.n2833 gnd.n2729 19.3944
R16446 gnd.n2833 gnd.n2832 19.3944
R16447 gnd.n2832 gnd.n2737 19.3944
R16448 gnd.n2825 gnd.n2737 19.3944
R16449 gnd.n2825 gnd.n2824 19.3944
R16450 gnd.n2824 gnd.n2748 19.3944
R16451 gnd.n2817 gnd.n2748 19.3944
R16452 gnd.n2817 gnd.n2816 19.3944
R16453 gnd.n2816 gnd.n2759 19.3944
R16454 gnd.n2809 gnd.n2759 19.3944
R16455 gnd.n2809 gnd.n2808 19.3944
R16456 gnd.n2808 gnd.n2771 19.3944
R16457 gnd.n2801 gnd.n2771 19.3944
R16458 gnd.n2801 gnd.n2800 19.3944
R16459 gnd.n7184 gnd.n445 19.3944
R16460 gnd.n7190 gnd.n445 19.3944
R16461 gnd.n7190 gnd.n443 19.3944
R16462 gnd.n7194 gnd.n443 19.3944
R16463 gnd.n7194 gnd.n439 19.3944
R16464 gnd.n7200 gnd.n439 19.3944
R16465 gnd.n7200 gnd.n437 19.3944
R16466 gnd.n7204 gnd.n437 19.3944
R16467 gnd.n7204 gnd.n433 19.3944
R16468 gnd.n7210 gnd.n433 19.3944
R16469 gnd.n7210 gnd.n431 19.3944
R16470 gnd.n7214 gnd.n431 19.3944
R16471 gnd.n7214 gnd.n427 19.3944
R16472 gnd.n7220 gnd.n427 19.3944
R16473 gnd.n7220 gnd.n425 19.3944
R16474 gnd.n7224 gnd.n425 19.3944
R16475 gnd.n7224 gnd.n421 19.3944
R16476 gnd.n7230 gnd.n421 19.3944
R16477 gnd.n7230 gnd.n419 19.3944
R16478 gnd.n7234 gnd.n419 19.3944
R16479 gnd.n7234 gnd.n415 19.3944
R16480 gnd.n7240 gnd.n415 19.3944
R16481 gnd.n7240 gnd.n413 19.3944
R16482 gnd.n7244 gnd.n413 19.3944
R16483 gnd.n7244 gnd.n409 19.3944
R16484 gnd.n7250 gnd.n409 19.3944
R16485 gnd.n7250 gnd.n407 19.3944
R16486 gnd.n7254 gnd.n407 19.3944
R16487 gnd.n7254 gnd.n403 19.3944
R16488 gnd.n7260 gnd.n403 19.3944
R16489 gnd.n7260 gnd.n401 19.3944
R16490 gnd.n7264 gnd.n401 19.3944
R16491 gnd.n7264 gnd.n397 19.3944
R16492 gnd.n7270 gnd.n397 19.3944
R16493 gnd.n7270 gnd.n395 19.3944
R16494 gnd.n7274 gnd.n395 19.3944
R16495 gnd.n7274 gnd.n391 19.3944
R16496 gnd.n7280 gnd.n391 19.3944
R16497 gnd.n7280 gnd.n389 19.3944
R16498 gnd.n7284 gnd.n389 19.3944
R16499 gnd.n7284 gnd.n385 19.3944
R16500 gnd.n7290 gnd.n385 19.3944
R16501 gnd.n7290 gnd.n383 19.3944
R16502 gnd.n7294 gnd.n383 19.3944
R16503 gnd.n7294 gnd.n379 19.3944
R16504 gnd.n7300 gnd.n379 19.3944
R16505 gnd.n7300 gnd.n377 19.3944
R16506 gnd.n7304 gnd.n377 19.3944
R16507 gnd.n7304 gnd.n373 19.3944
R16508 gnd.n7310 gnd.n373 19.3944
R16509 gnd.n7310 gnd.n371 19.3944
R16510 gnd.n7314 gnd.n371 19.3944
R16511 gnd.n7314 gnd.n367 19.3944
R16512 gnd.n7320 gnd.n367 19.3944
R16513 gnd.n7320 gnd.n365 19.3944
R16514 gnd.n7324 gnd.n365 19.3944
R16515 gnd.n7324 gnd.n361 19.3944
R16516 gnd.n7330 gnd.n361 19.3944
R16517 gnd.n7330 gnd.n359 19.3944
R16518 gnd.n7334 gnd.n359 19.3944
R16519 gnd.n7334 gnd.n355 19.3944
R16520 gnd.n7340 gnd.n355 19.3944
R16521 gnd.n7340 gnd.n353 19.3944
R16522 gnd.n7344 gnd.n353 19.3944
R16523 gnd.n7344 gnd.n349 19.3944
R16524 gnd.n7350 gnd.n349 19.3944
R16525 gnd.n7350 gnd.n347 19.3944
R16526 gnd.n7354 gnd.n347 19.3944
R16527 gnd.n7354 gnd.n343 19.3944
R16528 gnd.n7360 gnd.n343 19.3944
R16529 gnd.n7360 gnd.n341 19.3944
R16530 gnd.n7364 gnd.n341 19.3944
R16531 gnd.n7364 gnd.n337 19.3944
R16532 gnd.n7370 gnd.n337 19.3944
R16533 gnd.n7370 gnd.n335 19.3944
R16534 gnd.n7374 gnd.n335 19.3944
R16535 gnd.n7374 gnd.n331 19.3944
R16536 gnd.n7380 gnd.n331 19.3944
R16537 gnd.n7380 gnd.n329 19.3944
R16538 gnd.n7384 gnd.n329 19.3944
R16539 gnd.n7384 gnd.n325 19.3944
R16540 gnd.n7391 gnd.n325 19.3944
R16541 gnd.n7391 gnd.n323 19.3944
R16542 gnd.n7395 gnd.n323 19.3944
R16543 gnd.n6699 gnd.n738 19.3944
R16544 gnd.n6699 gnd.n736 19.3944
R16545 gnd.n6703 gnd.n736 19.3944
R16546 gnd.n6703 gnd.n732 19.3944
R16547 gnd.n6709 gnd.n732 19.3944
R16548 gnd.n6709 gnd.n730 19.3944
R16549 gnd.n6713 gnd.n730 19.3944
R16550 gnd.n6713 gnd.n726 19.3944
R16551 gnd.n6719 gnd.n726 19.3944
R16552 gnd.n6719 gnd.n724 19.3944
R16553 gnd.n6723 gnd.n724 19.3944
R16554 gnd.n6723 gnd.n720 19.3944
R16555 gnd.n6729 gnd.n720 19.3944
R16556 gnd.n6729 gnd.n718 19.3944
R16557 gnd.n6733 gnd.n718 19.3944
R16558 gnd.n6733 gnd.n714 19.3944
R16559 gnd.n6739 gnd.n714 19.3944
R16560 gnd.n6739 gnd.n712 19.3944
R16561 gnd.n6743 gnd.n712 19.3944
R16562 gnd.n6743 gnd.n708 19.3944
R16563 gnd.n6749 gnd.n708 19.3944
R16564 gnd.n6749 gnd.n706 19.3944
R16565 gnd.n6753 gnd.n706 19.3944
R16566 gnd.n6753 gnd.n702 19.3944
R16567 gnd.n6759 gnd.n702 19.3944
R16568 gnd.n6759 gnd.n700 19.3944
R16569 gnd.n6763 gnd.n700 19.3944
R16570 gnd.n6763 gnd.n696 19.3944
R16571 gnd.n6769 gnd.n696 19.3944
R16572 gnd.n6769 gnd.n694 19.3944
R16573 gnd.n6773 gnd.n694 19.3944
R16574 gnd.n6773 gnd.n690 19.3944
R16575 gnd.n6779 gnd.n690 19.3944
R16576 gnd.n6779 gnd.n688 19.3944
R16577 gnd.n6783 gnd.n688 19.3944
R16578 gnd.n6783 gnd.n684 19.3944
R16579 gnd.n6789 gnd.n684 19.3944
R16580 gnd.n6789 gnd.n682 19.3944
R16581 gnd.n6793 gnd.n682 19.3944
R16582 gnd.n6793 gnd.n678 19.3944
R16583 gnd.n6799 gnd.n678 19.3944
R16584 gnd.n6799 gnd.n676 19.3944
R16585 gnd.n6803 gnd.n676 19.3944
R16586 gnd.n6803 gnd.n672 19.3944
R16587 gnd.n6809 gnd.n672 19.3944
R16588 gnd.n6809 gnd.n670 19.3944
R16589 gnd.n6813 gnd.n670 19.3944
R16590 gnd.n6813 gnd.n666 19.3944
R16591 gnd.n6819 gnd.n666 19.3944
R16592 gnd.n6819 gnd.n664 19.3944
R16593 gnd.n6823 gnd.n664 19.3944
R16594 gnd.n6823 gnd.n660 19.3944
R16595 gnd.n6829 gnd.n660 19.3944
R16596 gnd.n6829 gnd.n658 19.3944
R16597 gnd.n6833 gnd.n658 19.3944
R16598 gnd.n6833 gnd.n654 19.3944
R16599 gnd.n6839 gnd.n654 19.3944
R16600 gnd.n6839 gnd.n652 19.3944
R16601 gnd.n6843 gnd.n652 19.3944
R16602 gnd.n6843 gnd.n648 19.3944
R16603 gnd.n6849 gnd.n648 19.3944
R16604 gnd.n6849 gnd.n646 19.3944
R16605 gnd.n6853 gnd.n646 19.3944
R16606 gnd.n6853 gnd.n642 19.3944
R16607 gnd.n6859 gnd.n642 19.3944
R16608 gnd.n6859 gnd.n640 19.3944
R16609 gnd.n6863 gnd.n640 19.3944
R16610 gnd.n6863 gnd.n636 19.3944
R16611 gnd.n6869 gnd.n636 19.3944
R16612 gnd.n6869 gnd.n634 19.3944
R16613 gnd.n6873 gnd.n634 19.3944
R16614 gnd.n6873 gnd.n630 19.3944
R16615 gnd.n6879 gnd.n630 19.3944
R16616 gnd.n6879 gnd.n628 19.3944
R16617 gnd.n6883 gnd.n628 19.3944
R16618 gnd.n6883 gnd.n624 19.3944
R16619 gnd.n6889 gnd.n624 19.3944
R16620 gnd.n6889 gnd.n622 19.3944
R16621 gnd.n6893 gnd.n622 19.3944
R16622 gnd.n6893 gnd.n618 19.3944
R16623 gnd.n6899 gnd.n618 19.3944
R16624 gnd.n6899 gnd.n616 19.3944
R16625 gnd.n6903 gnd.n616 19.3944
R16626 gnd.n6903 gnd.n612 19.3944
R16627 gnd.n6909 gnd.n612 19.3944
R16628 gnd.n6909 gnd.n610 19.3944
R16629 gnd.n6913 gnd.n610 19.3944
R16630 gnd.n6913 gnd.n606 19.3944
R16631 gnd.n6919 gnd.n606 19.3944
R16632 gnd.n6919 gnd.n604 19.3944
R16633 gnd.n6923 gnd.n604 19.3944
R16634 gnd.n6923 gnd.n600 19.3944
R16635 gnd.n6929 gnd.n600 19.3944
R16636 gnd.n6929 gnd.n598 19.3944
R16637 gnd.n6933 gnd.n598 19.3944
R16638 gnd.n6933 gnd.n594 19.3944
R16639 gnd.n6939 gnd.n594 19.3944
R16640 gnd.n6939 gnd.n592 19.3944
R16641 gnd.n6943 gnd.n592 19.3944
R16642 gnd.n6943 gnd.n588 19.3944
R16643 gnd.n6949 gnd.n588 19.3944
R16644 gnd.n6949 gnd.n586 19.3944
R16645 gnd.n6953 gnd.n586 19.3944
R16646 gnd.n6953 gnd.n582 19.3944
R16647 gnd.n6959 gnd.n582 19.3944
R16648 gnd.n6959 gnd.n580 19.3944
R16649 gnd.n6963 gnd.n580 19.3944
R16650 gnd.n6963 gnd.n576 19.3944
R16651 gnd.n6969 gnd.n576 19.3944
R16652 gnd.n6969 gnd.n574 19.3944
R16653 gnd.n6973 gnd.n574 19.3944
R16654 gnd.n6973 gnd.n570 19.3944
R16655 gnd.n6979 gnd.n570 19.3944
R16656 gnd.n6979 gnd.n568 19.3944
R16657 gnd.n6983 gnd.n568 19.3944
R16658 gnd.n6983 gnd.n564 19.3944
R16659 gnd.n6989 gnd.n564 19.3944
R16660 gnd.n6989 gnd.n562 19.3944
R16661 gnd.n6993 gnd.n562 19.3944
R16662 gnd.n6993 gnd.n558 19.3944
R16663 gnd.n6999 gnd.n558 19.3944
R16664 gnd.n6999 gnd.n556 19.3944
R16665 gnd.n7003 gnd.n556 19.3944
R16666 gnd.n7003 gnd.n552 19.3944
R16667 gnd.n7009 gnd.n552 19.3944
R16668 gnd.n7009 gnd.n550 19.3944
R16669 gnd.n7013 gnd.n550 19.3944
R16670 gnd.n7013 gnd.n546 19.3944
R16671 gnd.n7019 gnd.n546 19.3944
R16672 gnd.n7019 gnd.n544 19.3944
R16673 gnd.n7023 gnd.n544 19.3944
R16674 gnd.n7023 gnd.n540 19.3944
R16675 gnd.n7029 gnd.n540 19.3944
R16676 gnd.n7029 gnd.n538 19.3944
R16677 gnd.n7033 gnd.n538 19.3944
R16678 gnd.n7033 gnd.n534 19.3944
R16679 gnd.n7039 gnd.n534 19.3944
R16680 gnd.n7039 gnd.n532 19.3944
R16681 gnd.n7043 gnd.n532 19.3944
R16682 gnd.n7043 gnd.n528 19.3944
R16683 gnd.n7049 gnd.n528 19.3944
R16684 gnd.n7049 gnd.n526 19.3944
R16685 gnd.n7053 gnd.n526 19.3944
R16686 gnd.n7053 gnd.n522 19.3944
R16687 gnd.n7059 gnd.n522 19.3944
R16688 gnd.n7059 gnd.n520 19.3944
R16689 gnd.n7063 gnd.n520 19.3944
R16690 gnd.n7063 gnd.n516 19.3944
R16691 gnd.n7069 gnd.n516 19.3944
R16692 gnd.n7069 gnd.n514 19.3944
R16693 gnd.n7073 gnd.n514 19.3944
R16694 gnd.n7073 gnd.n510 19.3944
R16695 gnd.n7079 gnd.n510 19.3944
R16696 gnd.n7079 gnd.n508 19.3944
R16697 gnd.n7083 gnd.n508 19.3944
R16698 gnd.n7083 gnd.n504 19.3944
R16699 gnd.n7089 gnd.n504 19.3944
R16700 gnd.n7089 gnd.n502 19.3944
R16701 gnd.n7093 gnd.n502 19.3944
R16702 gnd.n7093 gnd.n498 19.3944
R16703 gnd.n7099 gnd.n498 19.3944
R16704 gnd.n7099 gnd.n496 19.3944
R16705 gnd.n7103 gnd.n496 19.3944
R16706 gnd.n7103 gnd.n492 19.3944
R16707 gnd.n7109 gnd.n492 19.3944
R16708 gnd.n7109 gnd.n490 19.3944
R16709 gnd.n7113 gnd.n490 19.3944
R16710 gnd.n7113 gnd.n486 19.3944
R16711 gnd.n7119 gnd.n486 19.3944
R16712 gnd.n7119 gnd.n484 19.3944
R16713 gnd.n7123 gnd.n484 19.3944
R16714 gnd.n7123 gnd.n480 19.3944
R16715 gnd.n7129 gnd.n480 19.3944
R16716 gnd.n7129 gnd.n478 19.3944
R16717 gnd.n7133 gnd.n478 19.3944
R16718 gnd.n7133 gnd.n474 19.3944
R16719 gnd.n7139 gnd.n474 19.3944
R16720 gnd.n7139 gnd.n472 19.3944
R16721 gnd.n7143 gnd.n472 19.3944
R16722 gnd.n7143 gnd.n468 19.3944
R16723 gnd.n7149 gnd.n468 19.3944
R16724 gnd.n7149 gnd.n466 19.3944
R16725 gnd.n7153 gnd.n466 19.3944
R16726 gnd.n7153 gnd.n462 19.3944
R16727 gnd.n7159 gnd.n462 19.3944
R16728 gnd.n7159 gnd.n460 19.3944
R16729 gnd.n7163 gnd.n460 19.3944
R16730 gnd.n7163 gnd.n456 19.3944
R16731 gnd.n7169 gnd.n456 19.3944
R16732 gnd.n7169 gnd.n454 19.3944
R16733 gnd.n7174 gnd.n454 19.3944
R16734 gnd.n7174 gnd.n450 19.3944
R16735 gnd.n7180 gnd.n450 19.3944
R16736 gnd.n7181 gnd.n7180 19.3944
R16737 gnd.n1912 gnd.n1908 19.3944
R16738 gnd.n1912 gnd.n1905 19.3944
R16739 gnd.n1916 gnd.n1905 19.3944
R16740 gnd.n1916 gnd.n1903 19.3944
R16741 gnd.n1922 gnd.n1903 19.3944
R16742 gnd.n1922 gnd.n1901 19.3944
R16743 gnd.n1926 gnd.n1901 19.3944
R16744 gnd.n1926 gnd.n1899 19.3944
R16745 gnd.n1932 gnd.n1899 19.3944
R16746 gnd.n1932 gnd.n1897 19.3944
R16747 gnd.n1937 gnd.n1897 19.3944
R16748 gnd.n1937 gnd.n1895 19.3944
R16749 gnd.n1895 gnd.n1892 19.3944
R16750 gnd.n1944 gnd.n1892 19.3944
R16751 gnd.n1944 gnd.n1889 19.3944
R16752 gnd.n2029 gnd.n1951 19.3944
R16753 gnd.n2023 gnd.n1951 19.3944
R16754 gnd.n2023 gnd.n2022 19.3944
R16755 gnd.n2022 gnd.n2021 19.3944
R16756 gnd.n2021 gnd.n1957 19.3944
R16757 gnd.n2015 gnd.n1957 19.3944
R16758 gnd.n2015 gnd.n2014 19.3944
R16759 gnd.n2014 gnd.n2013 19.3944
R16760 gnd.n2013 gnd.n1963 19.3944
R16761 gnd.n2007 gnd.n1963 19.3944
R16762 gnd.n2007 gnd.n2006 19.3944
R16763 gnd.n2006 gnd.n2005 19.3944
R16764 gnd.n2005 gnd.n1969 19.3944
R16765 gnd.n1999 gnd.n1969 19.3944
R16766 gnd.n1999 gnd.n1998 19.3944
R16767 gnd.n1998 gnd.n1997 19.3944
R16768 gnd.n1997 gnd.n1975 19.3944
R16769 gnd.n1991 gnd.n1975 19.3944
R16770 gnd.n1983 gnd.n1640 19.3944
R16771 gnd.n4489 gnd.n1640 19.3944
R16772 gnd.n4490 gnd.n4489 19.3944
R16773 gnd.n4490 gnd.n1638 19.3944
R16774 gnd.n4518 gnd.n1638 19.3944
R16775 gnd.n4518 gnd.n4517 19.3944
R16776 gnd.n4517 gnd.n4516 19.3944
R16777 gnd.n4516 gnd.n4515 19.3944
R16778 gnd.n4515 gnd.n4514 19.3944
R16779 gnd.n4514 gnd.n4512 19.3944
R16780 gnd.n4512 gnd.n4511 19.3944
R16781 gnd.n4511 gnd.n4509 19.3944
R16782 gnd.n4509 gnd.n4508 19.3944
R16783 gnd.n4508 gnd.n4507 19.3944
R16784 gnd.n4507 gnd.n4505 19.3944
R16785 gnd.n4505 gnd.n1558 19.3944
R16786 gnd.n4614 gnd.n1558 19.3944
R16787 gnd.n4615 gnd.n4614 19.3944
R16788 gnd.n4617 gnd.n4615 19.3944
R16789 gnd.n4617 gnd.n1556 19.3944
R16790 gnd.n4623 gnd.n1556 19.3944
R16791 gnd.n4623 gnd.n4622 19.3944
R16792 gnd.n4622 gnd.n1550 19.3944
R16793 gnd.n4640 gnd.n1550 19.3944
R16794 gnd.n4640 gnd.n1548 19.3944
R16795 gnd.n4644 gnd.n1548 19.3944
R16796 gnd.n4644 gnd.n299 19.3944
R16797 gnd.n7478 gnd.n299 19.3944
R16798 gnd.n7478 gnd.n7477 19.3944
R16799 gnd.n7477 gnd.n7476 19.3944
R16800 gnd.n7476 gnd.n304 19.3944
R16801 gnd.n7408 gnd.n304 19.3944
R16802 gnd.n7408 gnd.n7404 19.3944
R16803 gnd.n7415 gnd.n7404 19.3944
R16804 gnd.n7416 gnd.n7415 19.3944
R16805 gnd.n7419 gnd.n7416 19.3944
R16806 gnd.n7419 gnd.n7402 19.3944
R16807 gnd.n7454 gnd.n7402 19.3944
R16808 gnd.n7454 gnd.n7453 19.3944
R16809 gnd.n7453 gnd.n7452 19.3944
R16810 gnd.n7452 gnd.n7449 19.3944
R16811 gnd.n7449 gnd.n7448 19.3944
R16812 gnd.n7448 gnd.n7446 19.3944
R16813 gnd.n7446 gnd.n7445 19.3944
R16814 gnd.n7445 gnd.n7443 19.3944
R16815 gnd.n7443 gnd.n7442 19.3944
R16816 gnd.n7442 gnd.n7440 19.3944
R16817 gnd.n7440 gnd.n7439 19.3944
R16818 gnd.n7439 gnd.n7437 19.3944
R16819 gnd.n7437 gnd.n7436 19.3944
R16820 gnd.n7436 gnd.n183 19.3944
R16821 gnd.n7666 gnd.n183 19.3944
R16822 gnd.n7667 gnd.n7666 19.3944
R16823 gnd.n7705 gnd.n144 19.3944
R16824 gnd.n7700 gnd.n144 19.3944
R16825 gnd.n7700 gnd.n7699 19.3944
R16826 gnd.n7699 gnd.n7698 19.3944
R16827 gnd.n7698 gnd.n151 19.3944
R16828 gnd.n7693 gnd.n151 19.3944
R16829 gnd.n7693 gnd.n7692 19.3944
R16830 gnd.n7692 gnd.n7691 19.3944
R16831 gnd.n7691 gnd.n158 19.3944
R16832 gnd.n7686 gnd.n158 19.3944
R16833 gnd.n7686 gnd.n7685 19.3944
R16834 gnd.n7685 gnd.n7684 19.3944
R16835 gnd.n7684 gnd.n165 19.3944
R16836 gnd.n7679 gnd.n165 19.3944
R16837 gnd.n7679 gnd.n7678 19.3944
R16838 gnd.n7678 gnd.n7677 19.3944
R16839 gnd.n7677 gnd.n172 19.3944
R16840 gnd.n7672 gnd.n172 19.3944
R16841 gnd.n7738 gnd.n7737 19.3944
R16842 gnd.n7737 gnd.n7736 19.3944
R16843 gnd.n7736 gnd.n115 19.3944
R16844 gnd.n7731 gnd.n115 19.3944
R16845 gnd.n7731 gnd.n7730 19.3944
R16846 gnd.n7730 gnd.n7729 19.3944
R16847 gnd.n7729 gnd.n123 19.3944
R16848 gnd.n7724 gnd.n123 19.3944
R16849 gnd.n7724 gnd.n7723 19.3944
R16850 gnd.n7723 gnd.n7722 19.3944
R16851 gnd.n7722 gnd.n130 19.3944
R16852 gnd.n7717 gnd.n130 19.3944
R16853 gnd.n7717 gnd.n7716 19.3944
R16854 gnd.n7716 gnd.n7715 19.3944
R16855 gnd.n7715 gnd.n137 19.3944
R16856 gnd.n7710 gnd.n137 19.3944
R16857 gnd.n7710 gnd.n7709 19.3944
R16858 gnd.n4722 gnd.n1484 19.3944
R16859 gnd.n4722 gnd.n4721 19.3944
R16860 gnd.n4721 gnd.n4720 19.3944
R16861 gnd.n4720 gnd.n1488 19.3944
R16862 gnd.n4526 gnd.n1488 19.3944
R16863 gnd.n4526 gnd.n4525 19.3944
R16864 gnd.n4525 gnd.n1603 19.3944
R16865 gnd.n4552 gnd.n1603 19.3944
R16866 gnd.n4552 gnd.n1601 19.3944
R16867 gnd.n4558 gnd.n1601 19.3944
R16868 gnd.n4558 gnd.n4557 19.3944
R16869 gnd.n4557 gnd.n1576 19.3944
R16870 gnd.n4591 gnd.n1576 19.3944
R16871 gnd.n4591 gnd.n1574 19.3944
R16872 gnd.n4597 gnd.n1574 19.3944
R16873 gnd.n4597 gnd.n4596 19.3944
R16874 gnd.n4596 gnd.n1524 19.3944
R16875 gnd.n4681 gnd.n1524 19.3944
R16876 gnd.n4681 gnd.n1522 19.3944
R16877 gnd.n4685 gnd.n1522 19.3944
R16878 gnd.n4685 gnd.n274 19.3944
R16879 gnd.n7503 gnd.n274 19.3944
R16880 gnd.n273 gnd.n272 19.3944
R16881 gnd.n4662 gnd.n272 19.3944
R16882 gnd.n1547 gnd.n1546 19.3944
R16883 gnd.n7483 gnd.n7482 19.3944
R16884 gnd.n7506 gnd.n266 19.3944
R16885 gnd.n7506 gnd.n253 19.3944
R16886 gnd.n7518 gnd.n253 19.3944
R16887 gnd.n7518 gnd.n251 19.3944
R16888 gnd.n7522 gnd.n251 19.3944
R16889 gnd.n7522 gnd.n237 19.3944
R16890 gnd.n7534 gnd.n237 19.3944
R16891 gnd.n7534 gnd.n235 19.3944
R16892 gnd.n7538 gnd.n235 19.3944
R16893 gnd.n7538 gnd.n223 19.3944
R16894 gnd.n7550 gnd.n223 19.3944
R16895 gnd.n7550 gnd.n221 19.3944
R16896 gnd.n7554 gnd.n221 19.3944
R16897 gnd.n7554 gnd.n206 19.3944
R16898 gnd.n7566 gnd.n206 19.3944
R16899 gnd.n7566 gnd.n204 19.3944
R16900 gnd.n7570 gnd.n204 19.3944
R16901 gnd.n7570 gnd.n191 19.3944
R16902 gnd.n7657 gnd.n191 19.3944
R16903 gnd.n7657 gnd.n189 19.3944
R16904 gnd.n7661 gnd.n189 19.3944
R16905 gnd.n7661 gnd.n110 19.3944
R16906 gnd.n7741 gnd.n110 19.3944
R16907 gnd.n2928 gnd.n2921 19.3944
R16908 gnd.n2928 gnd.n2919 19.3944
R16909 gnd.n2932 gnd.n2919 19.3944
R16910 gnd.n2932 gnd.n2917 19.3944
R16911 gnd.n3003 gnd.n2917 19.3944
R16912 gnd.n3003 gnd.n3002 19.3944
R16913 gnd.n3002 gnd.n3001 19.3944
R16914 gnd.n3001 gnd.n2938 19.3944
R16915 gnd.n2997 gnd.n2938 19.3944
R16916 gnd.n2992 gnd.n2940 19.3944
R16917 gnd.n2988 gnd.n2945 19.3944
R16918 gnd.n2986 gnd.n2985 19.3944
R16919 gnd.n2982 gnd.n2981 19.3944
R16920 gnd.n2978 gnd.n2977 19.3944
R16921 gnd.n2977 gnd.n2976 19.3944
R16922 gnd.n2976 gnd.n2948 19.3944
R16923 gnd.n2972 gnd.n2948 19.3944
R16924 gnd.n2972 gnd.n2971 19.3944
R16925 gnd.n2971 gnd.n2970 19.3944
R16926 gnd.n2970 gnd.n2954 19.3944
R16927 gnd.n2966 gnd.n2954 19.3944
R16928 gnd.n2966 gnd.n2965 19.3944
R16929 gnd.n2965 gnd.n2964 19.3944
R16930 gnd.n2964 gnd.n2961 19.3944
R16931 gnd.n2961 gnd.n2856 19.3944
R16932 gnd.n3302 gnd.n2856 19.3944
R16933 gnd.n3302 gnd.n2854 19.3944
R16934 gnd.n3306 gnd.n2854 19.3944
R16935 gnd.n3306 gnd.n2852 19.3944
R16936 gnd.n3310 gnd.n2852 19.3944
R16937 gnd.n3310 gnd.n2850 19.3944
R16938 gnd.n3314 gnd.n2850 19.3944
R16939 gnd.n3314 gnd.n2848 19.3944
R16940 gnd.n3318 gnd.n2848 19.3944
R16941 gnd.n3318 gnd.n2846 19.3944
R16942 gnd.n3322 gnd.n2846 19.3944
R16943 gnd.n3322 gnd.n2844 19.3944
R16944 gnd.n3329 gnd.n2844 19.3944
R16945 gnd.n3329 gnd.n2842 19.3944
R16946 gnd.n3333 gnd.n2842 19.3944
R16947 gnd.n3333 gnd.n2706 19.3944
R16948 gnd.n3342 gnd.n2706 19.3944
R16949 gnd.n3342 gnd.n2704 19.3944
R16950 gnd.n3346 gnd.n2704 19.3944
R16951 gnd.n3346 gnd.n2700 19.3944
R16952 gnd.n3358 gnd.n2700 19.3944
R16953 gnd.n3358 gnd.n2698 19.3944
R16954 gnd.n3362 gnd.n2698 19.3944
R16955 gnd.n3362 gnd.n2694 19.3944
R16956 gnd.n3374 gnd.n2694 19.3944
R16957 gnd.n3374 gnd.n2692 19.3944
R16958 gnd.n3378 gnd.n2692 19.3944
R16959 gnd.n3378 gnd.n2688 19.3944
R16960 gnd.n3390 gnd.n2688 19.3944
R16961 gnd.n3390 gnd.n2686 19.3944
R16962 gnd.n3394 gnd.n2686 19.3944
R16963 gnd.n3394 gnd.n2385 19.3944
R16964 gnd.n3566 gnd.n2385 19.3944
R16965 gnd.n3566 gnd.n2383 19.3944
R16966 gnd.n3570 gnd.n2383 19.3944
R16967 gnd.n3570 gnd.n2363 19.3944
R16968 gnd.n3594 gnd.n2363 19.3944
R16969 gnd.n3594 gnd.n2361 19.3944
R16970 gnd.n3600 gnd.n2361 19.3944
R16971 gnd.n3600 gnd.n3599 19.3944
R16972 gnd.n3599 gnd.n2335 19.3944
R16973 gnd.n3668 gnd.n2335 19.3944
R16974 gnd.n3668 gnd.n2333 19.3944
R16975 gnd.n3672 gnd.n2333 19.3944
R16976 gnd.n3672 gnd.n2315 19.3944
R16977 gnd.n3693 gnd.n2315 19.3944
R16978 gnd.n3693 gnd.n2313 19.3944
R16979 gnd.n3697 gnd.n2313 19.3944
R16980 gnd.n3697 gnd.n2295 19.3944
R16981 gnd.n3727 gnd.n2295 19.3944
R16982 gnd.n3727 gnd.n2293 19.3944
R16983 gnd.n3731 gnd.n2293 19.3944
R16984 gnd.n3731 gnd.n2278 19.3944
R16985 gnd.n3772 gnd.n2278 19.3944
R16986 gnd.n3772 gnd.n2276 19.3944
R16987 gnd.n3778 gnd.n2276 19.3944
R16988 gnd.n3778 gnd.n3777 19.3944
R16989 gnd.n3777 gnd.n2250 19.3944
R16990 gnd.n3845 gnd.n2250 19.3944
R16991 gnd.n3845 gnd.n2248 19.3944
R16992 gnd.n3849 gnd.n2248 19.3944
R16993 gnd.n3849 gnd.n2230 19.3944
R16994 gnd.n3871 gnd.n2230 19.3944
R16995 gnd.n3871 gnd.n2228 19.3944
R16996 gnd.n3875 gnd.n2228 19.3944
R16997 gnd.n3875 gnd.n2207 19.3944
R16998 gnd.n3904 gnd.n2207 19.3944
R16999 gnd.n3904 gnd.n2205 19.3944
R17000 gnd.n3908 gnd.n2205 19.3944
R17001 gnd.n3908 gnd.n2190 19.3944
R17002 gnd.n3950 gnd.n2190 19.3944
R17003 gnd.n3950 gnd.n2188 19.3944
R17004 gnd.n3956 gnd.n2188 19.3944
R17005 gnd.n3956 gnd.n3955 19.3944
R17006 gnd.n3955 gnd.n2163 19.3944
R17007 gnd.n4007 gnd.n2163 19.3944
R17008 gnd.n4007 gnd.n2161 19.3944
R17009 gnd.n4011 gnd.n2161 19.3944
R17010 gnd.n4011 gnd.n2142 19.3944
R17011 gnd.n4032 gnd.n2142 19.3944
R17012 gnd.n4032 gnd.n2140 19.3944
R17013 gnd.n4036 gnd.n2140 19.3944
R17014 gnd.n4036 gnd.n2120 19.3944
R17015 gnd.n4092 gnd.n2120 19.3944
R17016 gnd.n4092 gnd.n2118 19.3944
R17017 gnd.n4096 gnd.n2118 19.3944
R17018 gnd.n4096 gnd.n2098 19.3944
R17019 gnd.n4121 gnd.n2098 19.3944
R17020 gnd.n4121 gnd.n2096 19.3944
R17021 gnd.n4127 gnd.n2096 19.3944
R17022 gnd.n4127 gnd.n4126 19.3944
R17023 gnd.n4126 gnd.n2070 19.3944
R17024 gnd.n4171 gnd.n2070 19.3944
R17025 gnd.n4171 gnd.n2068 19.3944
R17026 gnd.n4175 gnd.n2068 19.3944
R17027 gnd.n4175 gnd.n2049 19.3944
R17028 gnd.n4197 gnd.n2049 19.3944
R17029 gnd.n4197 gnd.n2047 19.3944
R17030 gnd.n4203 gnd.n2047 19.3944
R17031 gnd.n4203 gnd.n4202 19.3944
R17032 gnd.n4202 gnd.n1845 19.3944
R17033 gnd.n4382 gnd.n1845 19.3944
R17034 gnd.n4382 gnd.n1843 19.3944
R17035 gnd.n4386 gnd.n1843 19.3944
R17036 gnd.n4386 gnd.n1832 19.3944
R17037 gnd.n4402 gnd.n1832 19.3944
R17038 gnd.n4402 gnd.n1830 19.3944
R17039 gnd.n4406 gnd.n1830 19.3944
R17040 gnd.n4406 gnd.n1819 19.3944
R17041 gnd.n4422 gnd.n1819 19.3944
R17042 gnd.n4422 gnd.n1817 19.3944
R17043 gnd.n4426 gnd.n1817 19.3944
R17044 gnd.n4426 gnd.n1806 19.3944
R17045 gnd.n4445 gnd.n1806 19.3944
R17046 gnd.n4445 gnd.n1804 19.3944
R17047 gnd.n4450 gnd.n1804 19.3944
R17048 gnd.n4450 gnd.n1461 19.3944
R17049 gnd.n4737 gnd.n1461 19.3944
R17050 gnd.n4737 gnd.n4736 19.3944
R17051 gnd.n4736 gnd.n4735 19.3944
R17052 gnd.n4735 gnd.n1465 19.3944
R17053 gnd.n4729 gnd.n1465 19.3944
R17054 gnd.n4729 gnd.n4728 19.3944
R17055 gnd.n4728 gnd.n4727 19.3944
R17056 gnd.n4727 gnd.n1474 19.3944
R17057 gnd.n1628 gnd.n1474 19.3944
R17058 gnd.n1628 gnd.n1625 19.3944
R17059 gnd.n1632 gnd.n1625 19.3944
R17060 gnd.n1632 gnd.n1614 19.3944
R17061 gnd.n4540 gnd.n1614 19.3944
R17062 gnd.n4540 gnd.n1612 19.3944
R17063 gnd.n4546 gnd.n1612 19.3944
R17064 gnd.n4546 gnd.n4545 19.3944
R17065 gnd.n4545 gnd.n1587 19.3944
R17066 gnd.n4573 gnd.n1587 19.3944
R17067 gnd.n4573 gnd.n1585 19.3944
R17068 gnd.n4586 gnd.n1585 19.3944
R17069 gnd.n4586 gnd.n4585 19.3944
R17070 gnd.n4585 gnd.n4584 19.3944
R17071 gnd.n4584 gnd.n4581 19.3944
R17072 gnd.n4581 gnd.n1532 19.3944
R17073 gnd.n4676 gnd.n1532 19.3944
R17074 gnd.n4676 gnd.n4675 19.3944
R17075 gnd.n4675 gnd.n4674 19.3944
R17076 gnd.n4674 gnd.n1537 19.3944
R17077 gnd.n4670 gnd.n1537 19.3944
R17078 gnd.n4668 gnd.n4667 19.3944
R17079 gnd.n4657 gnd.n4651 19.3944
R17080 gnd.n4655 gnd.n4654 19.3944
R17081 gnd.n7471 gnd.n308 19.3944
R17082 gnd.n7469 gnd.n7468 19.3944
R17083 gnd.n7468 gnd.n310 19.3944
R17084 gnd.n7464 gnd.n310 19.3944
R17085 gnd.n7464 gnd.n7463 19.3944
R17086 gnd.n7463 gnd.n7462 19.3944
R17087 gnd.n7462 gnd.n316 19.3944
R17088 gnd.n7401 gnd.n316 19.3944
R17089 gnd.n7401 gnd.n7400 19.3944
R17090 gnd.n7400 gnd.n7399 19.3944
R17091 gnd.n5135 gnd.n5134 19.3944
R17092 gnd.n5134 gnd.n5133 19.3944
R17093 gnd.n5133 gnd.n5132 19.3944
R17094 gnd.n5132 gnd.n5130 19.3944
R17095 gnd.n5130 gnd.n5127 19.3944
R17096 gnd.n5127 gnd.n5126 19.3944
R17097 gnd.n5126 gnd.n5123 19.3944
R17098 gnd.n5123 gnd.n5122 19.3944
R17099 gnd.n5122 gnd.n5119 19.3944
R17100 gnd.n5119 gnd.n5118 19.3944
R17101 gnd.n5118 gnd.n5115 19.3944
R17102 gnd.n5115 gnd.n5114 19.3944
R17103 gnd.n5114 gnd.n5111 19.3944
R17104 gnd.n5111 gnd.n5110 19.3944
R17105 gnd.n5110 gnd.n5107 19.3944
R17106 gnd.n5107 gnd.n5106 19.3944
R17107 gnd.n5106 gnd.n5103 19.3944
R17108 gnd.n5101 gnd.n5098 19.3944
R17109 gnd.n5098 gnd.n5097 19.3944
R17110 gnd.n5097 gnd.n5094 19.3944
R17111 gnd.n5094 gnd.n5093 19.3944
R17112 gnd.n5093 gnd.n5090 19.3944
R17113 gnd.n5090 gnd.n5089 19.3944
R17114 gnd.n5089 gnd.n5086 19.3944
R17115 gnd.n5086 gnd.n5085 19.3944
R17116 gnd.n5085 gnd.n5082 19.3944
R17117 gnd.n5082 gnd.n5081 19.3944
R17118 gnd.n5081 gnd.n5078 19.3944
R17119 gnd.n5078 gnd.n5077 19.3944
R17120 gnd.n5077 gnd.n5074 19.3944
R17121 gnd.n5074 gnd.n5073 19.3944
R17122 gnd.n5073 gnd.n5070 19.3944
R17123 gnd.n5070 gnd.n5069 19.3944
R17124 gnd.n5069 gnd.n5066 19.3944
R17125 gnd.n5066 gnd.n5065 19.3944
R17126 gnd.n5058 gnd.n5057 19.3944
R17127 gnd.n5057 gnd.n1058 19.3944
R17128 gnd.n5053 gnd.n1058 19.3944
R17129 gnd.n5053 gnd.n1060 19.3944
R17130 gnd.n3125 gnd.n1060 19.3944
R17131 gnd.n3127 gnd.n3125 19.3944
R17132 gnd.n3127 gnd.n3123 19.3944
R17133 gnd.n3132 gnd.n3123 19.3944
R17134 gnd.n3133 gnd.n3132 19.3944
R17135 gnd.n3135 gnd.n3133 19.3944
R17136 gnd.n3135 gnd.n3121 19.3944
R17137 gnd.n3139 gnd.n3121 19.3944
R17138 gnd.n3139 gnd.n3011 19.3944
R17139 gnd.n3151 gnd.n3011 19.3944
R17140 gnd.n3151 gnd.n3009 19.3944
R17141 gnd.n3155 gnd.n3009 19.3944
R17142 gnd.n3155 gnd.n2914 19.3944
R17143 gnd.n3167 gnd.n2914 19.3944
R17144 gnd.n3167 gnd.n2912 19.3944
R17145 gnd.n3171 gnd.n2912 19.3944
R17146 gnd.n3171 gnd.n2907 19.3944
R17147 gnd.n3183 gnd.n2907 19.3944
R17148 gnd.n3183 gnd.n2905 19.3944
R17149 gnd.n3187 gnd.n2905 19.3944
R17150 gnd.n3187 gnd.n2900 19.3944
R17151 gnd.n3200 gnd.n2900 19.3944
R17152 gnd.n3200 gnd.n2897 19.3944
R17153 gnd.n3205 gnd.n2897 19.3944
R17154 gnd.n3205 gnd.n2892 19.3944
R17155 gnd.n3217 gnd.n2892 19.3944
R17156 gnd.n3217 gnd.n2890 19.3944
R17157 gnd.n3221 gnd.n2890 19.3944
R17158 gnd.n3221 gnd.n2885 19.3944
R17159 gnd.n3233 gnd.n2885 19.3944
R17160 gnd.n3233 gnd.n2883 19.3944
R17161 gnd.n3237 gnd.n2883 19.3944
R17162 gnd.n3237 gnd.n2878 19.3944
R17163 gnd.n3249 gnd.n2878 19.3944
R17164 gnd.n3249 gnd.n2876 19.3944
R17165 gnd.n3254 gnd.n2876 19.3944
R17166 gnd.n3254 gnd.n2870 19.3944
R17167 gnd.n3266 gnd.n2870 19.3944
R17168 gnd.n3267 gnd.n3266 19.3944
R17169 gnd.n3268 gnd.n3267 19.3944
R17170 gnd.n3268 gnd.n2868 19.3944
R17171 gnd.n3274 gnd.n2868 19.3944
R17172 gnd.n3275 gnd.n3274 19.3944
R17173 gnd.n3278 gnd.n3275 19.3944
R17174 gnd.n3278 gnd.n2866 19.3944
R17175 gnd.n3283 gnd.n2866 19.3944
R17176 gnd.n3283 gnd.n2640 19.3944
R17177 gnd.n3452 gnd.n2640 19.3944
R17178 gnd.n3453 gnd.n3452 19.3944
R17179 gnd.n3491 gnd.n2543 19.3944
R17180 gnd.n3491 gnd.n2550 19.3944
R17181 gnd.n2607 gnd.n2550 19.3944
R17182 gnd.n3484 gnd.n2607 19.3944
R17183 gnd.n3484 gnd.n3483 19.3944
R17184 gnd.n3483 gnd.n3482 19.3944
R17185 gnd.n3482 gnd.n2613 19.3944
R17186 gnd.n3477 gnd.n2613 19.3944
R17187 gnd.n3477 gnd.n3476 19.3944
R17188 gnd.n3476 gnd.n3475 19.3944
R17189 gnd.n3475 gnd.n2620 19.3944
R17190 gnd.n3470 gnd.n2620 19.3944
R17191 gnd.n3470 gnd.n3469 19.3944
R17192 gnd.n3469 gnd.n3468 19.3944
R17193 gnd.n3468 gnd.n2627 19.3944
R17194 gnd.n3463 gnd.n2627 19.3944
R17195 gnd.n3463 gnd.n3462 19.3944
R17196 gnd.n3462 gnd.n3461 19.3944
R17197 gnd.n2563 gnd.n2562 19.3944
R17198 gnd.n2603 gnd.n2562 19.3944
R17199 gnd.n2603 gnd.n2602 19.3944
R17200 gnd.n2602 gnd.n2601 19.3944
R17201 gnd.n2601 gnd.n2598 19.3944
R17202 gnd.n2598 gnd.n2597 19.3944
R17203 gnd.n2597 gnd.n2594 19.3944
R17204 gnd.n2594 gnd.n2593 19.3944
R17205 gnd.n2593 gnd.n2590 19.3944
R17206 gnd.n2590 gnd.n2589 19.3944
R17207 gnd.n2589 gnd.n2586 19.3944
R17208 gnd.n2586 gnd.n2585 19.3944
R17209 gnd.n2585 gnd.n2582 19.3944
R17210 gnd.n2582 gnd.n2581 19.3944
R17211 gnd.n2581 gnd.n2544 19.3944
R17212 gnd.n3092 gnd.n3023 19.3944
R17213 gnd.n3092 gnd.n3024 19.3944
R17214 gnd.n3088 gnd.n3024 19.3944
R17215 gnd.n3088 gnd.n1080 19.3944
R17216 gnd.n5043 gnd.n1080 19.3944
R17217 gnd.n5043 gnd.n5042 19.3944
R17218 gnd.n5042 gnd.n5041 19.3944
R17219 gnd.n5041 gnd.n1084 19.3944
R17220 gnd.n5031 gnd.n1084 19.3944
R17221 gnd.n5031 gnd.n5030 19.3944
R17222 gnd.n5030 gnd.n5029 19.3944
R17223 gnd.n5029 gnd.n1103 19.3944
R17224 gnd.n5019 gnd.n1103 19.3944
R17225 gnd.n5019 gnd.n5018 19.3944
R17226 gnd.n5018 gnd.n5017 19.3944
R17227 gnd.n5017 gnd.n1125 19.3944
R17228 gnd.n5007 gnd.n1125 19.3944
R17229 gnd.n5007 gnd.n5006 19.3944
R17230 gnd.n5006 gnd.n5005 19.3944
R17231 gnd.n5005 gnd.n1146 19.3944
R17232 gnd.n4995 gnd.n1146 19.3944
R17233 gnd.n4995 gnd.n4994 19.3944
R17234 gnd.n4994 gnd.n4993 19.3944
R17235 gnd.n4993 gnd.n1167 19.3944
R17236 gnd.n4983 gnd.n1167 19.3944
R17237 gnd.n4983 gnd.n4982 19.3944
R17238 gnd.n4982 gnd.n4981 19.3944
R17239 gnd.n4981 gnd.n1186 19.3944
R17240 gnd.n4970 gnd.n1186 19.3944
R17241 gnd.n4970 gnd.n4969 19.3944
R17242 gnd.n4969 gnd.n4968 19.3944
R17243 gnd.n4968 gnd.n1204 19.3944
R17244 gnd.n4958 gnd.n1204 19.3944
R17245 gnd.n4958 gnd.n4957 19.3944
R17246 gnd.n4957 gnd.n4956 19.3944
R17247 gnd.n4956 gnd.n1224 19.3944
R17248 gnd.n4946 gnd.n1224 19.3944
R17249 gnd.n4946 gnd.n4945 19.3944
R17250 gnd.n4945 gnd.n4944 19.3944
R17251 gnd.n4944 gnd.n1245 19.3944
R17252 gnd.n4934 gnd.n1245 19.3944
R17253 gnd.n4934 gnd.n4933 19.3944
R17254 gnd.n4933 gnd.n4932 19.3944
R17255 gnd.n4932 gnd.n1266 19.3944
R17256 gnd.n4922 gnd.n1266 19.3944
R17257 gnd.n4922 gnd.n4921 19.3944
R17258 gnd.n4921 gnd.n4920 19.3944
R17259 gnd.n4920 gnd.n1287 19.3944
R17260 gnd.n4910 gnd.n1287 19.3944
R17261 gnd.n4910 gnd.n4909 19.3944
R17262 gnd.n4909 gnd.n4908 19.3944
R17263 gnd.n4908 gnd.n1309 19.3944
R17264 gnd.n4898 gnd.n1309 19.3944
R17265 gnd.n3084 gnd.n3082 19.3944
R17266 gnd.n3082 gnd.n3079 19.3944
R17267 gnd.n3079 gnd.n3078 19.3944
R17268 gnd.n3078 gnd.n3075 19.3944
R17269 gnd.n3075 gnd.n3074 19.3944
R17270 gnd.n3074 gnd.n3071 19.3944
R17271 gnd.n3071 gnd.n3070 19.3944
R17272 gnd.n3070 gnd.n3067 19.3944
R17273 gnd.n3067 gnd.n3066 19.3944
R17274 gnd.n3066 gnd.n3063 19.3944
R17275 gnd.n3063 gnd.n3062 19.3944
R17276 gnd.n3062 gnd.n3059 19.3944
R17277 gnd.n3059 gnd.n3058 19.3944
R17278 gnd.n3058 gnd.n3055 19.3944
R17279 gnd.n3055 gnd.n3054 19.3944
R17280 gnd.n3054 gnd.n3051 19.3944
R17281 gnd.n3045 gnd.n3018 19.3944
R17282 gnd.n3103 gnd.n3018 19.3944
R17283 gnd.n3104 gnd.n3103 19.3944
R17284 gnd.n3106 gnd.n3104 19.3944
R17285 gnd.n3106 gnd.n3016 19.3944
R17286 gnd.n3111 gnd.n3016 19.3944
R17287 gnd.n3112 gnd.n3111 19.3944
R17288 gnd.n3114 gnd.n3112 19.3944
R17289 gnd.n3114 gnd.n3014 19.3944
R17290 gnd.n3119 gnd.n3014 19.3944
R17291 gnd.n3120 gnd.n3119 19.3944
R17292 gnd.n3143 gnd.n3120 19.3944
R17293 gnd.n3143 gnd.n3012 19.3944
R17294 gnd.n3147 gnd.n3012 19.3944
R17295 gnd.n3147 gnd.n3008 19.3944
R17296 gnd.n3159 gnd.n3008 19.3944
R17297 gnd.n3159 gnd.n3006 19.3944
R17298 gnd.n3163 gnd.n3006 19.3944
R17299 gnd.n3163 gnd.n2910 19.3944
R17300 gnd.n3175 gnd.n2910 19.3944
R17301 gnd.n3175 gnd.n2908 19.3944
R17302 gnd.n3179 gnd.n2908 19.3944
R17303 gnd.n3179 gnd.n2904 19.3944
R17304 gnd.n3191 gnd.n2904 19.3944
R17305 gnd.n3191 gnd.n2902 19.3944
R17306 gnd.n3196 gnd.n2902 19.3944
R17307 gnd.n3196 gnd.n2895 19.3944
R17308 gnd.n3209 gnd.n2895 19.3944
R17309 gnd.n3209 gnd.n2893 19.3944
R17310 gnd.n3213 gnd.n2893 19.3944
R17311 gnd.n3213 gnd.n2889 19.3944
R17312 gnd.n3225 gnd.n2889 19.3944
R17313 gnd.n3225 gnd.n2887 19.3944
R17314 gnd.n3229 gnd.n2887 19.3944
R17315 gnd.n3229 gnd.n2881 19.3944
R17316 gnd.n3241 gnd.n2881 19.3944
R17317 gnd.n3241 gnd.n2879 19.3944
R17318 gnd.n3245 gnd.n2879 19.3944
R17319 gnd.n3245 gnd.n2875 19.3944
R17320 gnd.n3258 gnd.n2875 19.3944
R17321 gnd.n3258 gnd.n2873 19.3944
R17322 gnd.n3262 gnd.n2873 19.3944
R17323 gnd.n3262 gnd.n2859 19.3944
R17324 gnd.n3297 gnd.n2859 19.3944
R17325 gnd.n3297 gnd.n2860 19.3944
R17326 gnd.n3293 gnd.n2860 19.3944
R17327 gnd.n3293 gnd.n3292 19.3944
R17328 gnd.n3292 gnd.n3291 19.3944
R17329 gnd.n3291 gnd.n2865 19.3944
R17330 gnd.n3287 gnd.n2865 19.3944
R17331 gnd.n3287 gnd.n2642 19.3944
R17332 gnd.n3448 gnd.n2642 19.3944
R17333 gnd.n3448 gnd.n2643 19.3944
R17334 gnd.n3098 gnd.n3094 19.3944
R17335 gnd.n3098 gnd.n1069 19.3944
R17336 gnd.n5049 gnd.n1069 19.3944
R17337 gnd.n5049 gnd.n5048 19.3944
R17338 gnd.n5048 gnd.n5047 19.3944
R17339 gnd.n5047 gnd.n1073 19.3944
R17340 gnd.n5037 gnd.n1073 19.3944
R17341 gnd.n5037 gnd.n5036 19.3944
R17342 gnd.n5036 gnd.n5035 19.3944
R17343 gnd.n5035 gnd.n1094 19.3944
R17344 gnd.n5025 gnd.n1094 19.3944
R17345 gnd.n5025 gnd.n5024 19.3944
R17346 gnd.n5024 gnd.n5023 19.3944
R17347 gnd.n5023 gnd.n1114 19.3944
R17348 gnd.n5013 gnd.n1114 19.3944
R17349 gnd.n5013 gnd.n5012 19.3944
R17350 gnd.n5012 gnd.n5011 19.3944
R17351 gnd.n5011 gnd.n1136 19.3944
R17352 gnd.n5001 gnd.n1136 19.3944
R17353 gnd.n5001 gnd.n5000 19.3944
R17354 gnd.n5000 gnd.n4999 19.3944
R17355 gnd.n4999 gnd.n1156 19.3944
R17356 gnd.n4989 gnd.n4988 19.3944
R17357 gnd.n4988 gnd.n4987 19.3944
R17358 gnd.n4977 gnd.n1192 19.3944
R17359 gnd.n4975 gnd.n4974 19.3944
R17360 gnd.n4964 gnd.n1211 19.3944
R17361 gnd.n4964 gnd.n4963 19.3944
R17362 gnd.n4963 gnd.n4962 19.3944
R17363 gnd.n4962 gnd.n1214 19.3944
R17364 gnd.n4952 gnd.n1214 19.3944
R17365 gnd.n4952 gnd.n4951 19.3944
R17366 gnd.n4951 gnd.n4950 19.3944
R17367 gnd.n4950 gnd.n1234 19.3944
R17368 gnd.n4940 gnd.n1234 19.3944
R17369 gnd.n4940 gnd.n4939 19.3944
R17370 gnd.n4939 gnd.n4938 19.3944
R17371 gnd.n4938 gnd.n1256 19.3944
R17372 gnd.n4928 gnd.n1256 19.3944
R17373 gnd.n4928 gnd.n4927 19.3944
R17374 gnd.n4927 gnd.n4926 19.3944
R17375 gnd.n4926 gnd.n1276 19.3944
R17376 gnd.n4916 gnd.n1276 19.3944
R17377 gnd.n4916 gnd.n4915 19.3944
R17378 gnd.n4915 gnd.n4914 19.3944
R17379 gnd.n4914 gnd.n1298 19.3944
R17380 gnd.n4904 gnd.n1298 19.3944
R17381 gnd.n4904 gnd.n4903 19.3944
R17382 gnd.n4903 gnd.n4902 19.3944
R17383 gnd.n6693 gnd.n6692 19.3944
R17384 gnd.n6692 gnd.n6691 19.3944
R17385 gnd.n6691 gnd.n745 19.3944
R17386 gnd.n6685 gnd.n745 19.3944
R17387 gnd.n6685 gnd.n6684 19.3944
R17388 gnd.n6684 gnd.n6683 19.3944
R17389 gnd.n6683 gnd.n753 19.3944
R17390 gnd.n6677 gnd.n753 19.3944
R17391 gnd.n6677 gnd.n6676 19.3944
R17392 gnd.n6676 gnd.n6675 19.3944
R17393 gnd.n6675 gnd.n761 19.3944
R17394 gnd.n6669 gnd.n761 19.3944
R17395 gnd.n6669 gnd.n6668 19.3944
R17396 gnd.n6668 gnd.n6667 19.3944
R17397 gnd.n6667 gnd.n769 19.3944
R17398 gnd.n6661 gnd.n769 19.3944
R17399 gnd.n6661 gnd.n6660 19.3944
R17400 gnd.n6660 gnd.n6659 19.3944
R17401 gnd.n6659 gnd.n777 19.3944
R17402 gnd.n6653 gnd.n777 19.3944
R17403 gnd.n6653 gnd.n6652 19.3944
R17404 gnd.n6652 gnd.n6651 19.3944
R17405 gnd.n6651 gnd.n785 19.3944
R17406 gnd.n6645 gnd.n785 19.3944
R17407 gnd.n6645 gnd.n6644 19.3944
R17408 gnd.n6644 gnd.n6643 19.3944
R17409 gnd.n6643 gnd.n793 19.3944
R17410 gnd.n6637 gnd.n793 19.3944
R17411 gnd.n6637 gnd.n6636 19.3944
R17412 gnd.n6636 gnd.n6635 19.3944
R17413 gnd.n6635 gnd.n801 19.3944
R17414 gnd.n6629 gnd.n801 19.3944
R17415 gnd.n6629 gnd.n6628 19.3944
R17416 gnd.n6628 gnd.n6627 19.3944
R17417 gnd.n6627 gnd.n809 19.3944
R17418 gnd.n6621 gnd.n809 19.3944
R17419 gnd.n6621 gnd.n6620 19.3944
R17420 gnd.n6620 gnd.n6619 19.3944
R17421 gnd.n6619 gnd.n817 19.3944
R17422 gnd.n6613 gnd.n817 19.3944
R17423 gnd.n6613 gnd.n6612 19.3944
R17424 gnd.n6612 gnd.n6611 19.3944
R17425 gnd.n6611 gnd.n825 19.3944
R17426 gnd.n6605 gnd.n825 19.3944
R17427 gnd.n6605 gnd.n6604 19.3944
R17428 gnd.n6604 gnd.n6603 19.3944
R17429 gnd.n6603 gnd.n833 19.3944
R17430 gnd.n6597 gnd.n833 19.3944
R17431 gnd.n6597 gnd.n6596 19.3944
R17432 gnd.n6596 gnd.n6595 19.3944
R17433 gnd.n6595 gnd.n841 19.3944
R17434 gnd.n6589 gnd.n841 19.3944
R17435 gnd.n6589 gnd.n6588 19.3944
R17436 gnd.n6588 gnd.n6587 19.3944
R17437 gnd.n6587 gnd.n849 19.3944
R17438 gnd.n6581 gnd.n849 19.3944
R17439 gnd.n6581 gnd.n6580 19.3944
R17440 gnd.n6580 gnd.n6579 19.3944
R17441 gnd.n6579 gnd.n857 19.3944
R17442 gnd.n6573 gnd.n857 19.3944
R17443 gnd.n6573 gnd.n6572 19.3944
R17444 gnd.n6572 gnd.n6571 19.3944
R17445 gnd.n6571 gnd.n865 19.3944
R17446 gnd.n6565 gnd.n865 19.3944
R17447 gnd.n6565 gnd.n6564 19.3944
R17448 gnd.n6564 gnd.n6563 19.3944
R17449 gnd.n6563 gnd.n873 19.3944
R17450 gnd.n6557 gnd.n873 19.3944
R17451 gnd.n6557 gnd.n6556 19.3944
R17452 gnd.n6556 gnd.n6555 19.3944
R17453 gnd.n6555 gnd.n881 19.3944
R17454 gnd.n6549 gnd.n881 19.3944
R17455 gnd.n6549 gnd.n6548 19.3944
R17456 gnd.n6548 gnd.n6547 19.3944
R17457 gnd.n6547 gnd.n889 19.3944
R17458 gnd.n6541 gnd.n889 19.3944
R17459 gnd.n6541 gnd.n6540 19.3944
R17460 gnd.n6540 gnd.n6539 19.3944
R17461 gnd.n6539 gnd.n897 19.3944
R17462 gnd.n6533 gnd.n897 19.3944
R17463 gnd.n6533 gnd.n6532 19.3944
R17464 gnd.n6532 gnd.n6531 19.3944
R17465 gnd.n6531 gnd.n905 19.3944
R17466 gnd.n2924 gnd.n905 19.3944
R17467 gnd.n4893 gnd.n4892 19.3944
R17468 gnd.n4892 gnd.n4891 19.3944
R17469 gnd.n4891 gnd.n1332 19.3944
R17470 gnd.n4887 gnd.n1332 19.3944
R17471 gnd.n4887 gnd.n4886 19.3944
R17472 gnd.n4886 gnd.n4885 19.3944
R17473 gnd.n4885 gnd.n1337 19.3944
R17474 gnd.n4881 gnd.n1337 19.3944
R17475 gnd.n4881 gnd.n4880 19.3944
R17476 gnd.n4880 gnd.n4879 19.3944
R17477 gnd.n4879 gnd.n1342 19.3944
R17478 gnd.n4875 gnd.n1342 19.3944
R17479 gnd.n4875 gnd.n4874 19.3944
R17480 gnd.n4874 gnd.n4873 19.3944
R17481 gnd.n4873 gnd.n1347 19.3944
R17482 gnd.n4869 gnd.n1347 19.3944
R17483 gnd.n4869 gnd.n4868 19.3944
R17484 gnd.n4868 gnd.n4867 19.3944
R17485 gnd.n4867 gnd.n1352 19.3944
R17486 gnd.n4863 gnd.n1352 19.3944
R17487 gnd.n4863 gnd.n4862 19.3944
R17488 gnd.n4862 gnd.n4861 19.3944
R17489 gnd.n4861 gnd.n1357 19.3944
R17490 gnd.n4857 gnd.n1357 19.3944
R17491 gnd.n4857 gnd.n4856 19.3944
R17492 gnd.n4856 gnd.n4855 19.3944
R17493 gnd.n4855 gnd.n1362 19.3944
R17494 gnd.n4851 gnd.n1362 19.3944
R17495 gnd.n4851 gnd.n4850 19.3944
R17496 gnd.n4850 gnd.n4849 19.3944
R17497 gnd.n4849 gnd.n1367 19.3944
R17498 gnd.n4845 gnd.n1367 19.3944
R17499 gnd.n4845 gnd.n4844 19.3944
R17500 gnd.n4844 gnd.n4843 19.3944
R17501 gnd.n4843 gnd.n1372 19.3944
R17502 gnd.n4839 gnd.n1372 19.3944
R17503 gnd.n4839 gnd.n4838 19.3944
R17504 gnd.n4838 gnd.n4837 19.3944
R17505 gnd.n4837 gnd.n1377 19.3944
R17506 gnd.n4833 gnd.n1377 19.3944
R17507 gnd.n4833 gnd.n4832 19.3944
R17508 gnd.n4832 gnd.n4831 19.3944
R17509 gnd.n4831 gnd.n1382 19.3944
R17510 gnd.n4827 gnd.n1382 19.3944
R17511 gnd.n4827 gnd.n4826 19.3944
R17512 gnd.n4826 gnd.n4825 19.3944
R17513 gnd.n4825 gnd.n1387 19.3944
R17514 gnd.n4821 gnd.n1387 19.3944
R17515 gnd.n4821 gnd.n4820 19.3944
R17516 gnd.n4820 gnd.n4819 19.3944
R17517 gnd.n4819 gnd.n1392 19.3944
R17518 gnd.n4815 gnd.n1392 19.3944
R17519 gnd.n4815 gnd.n4814 19.3944
R17520 gnd.n4814 gnd.n4813 19.3944
R17521 gnd.n4813 gnd.n1397 19.3944
R17522 gnd.n4809 gnd.n1397 19.3944
R17523 gnd.n4809 gnd.n4808 19.3944
R17524 gnd.n4808 gnd.n4807 19.3944
R17525 gnd.n4807 gnd.n1402 19.3944
R17526 gnd.n4803 gnd.n1402 19.3944
R17527 gnd.n4803 gnd.n4802 19.3944
R17528 gnd.n4802 gnd.n4801 19.3944
R17529 gnd.n4801 gnd.n1407 19.3944
R17530 gnd.n4797 gnd.n1407 19.3944
R17531 gnd.n4797 gnd.n4796 19.3944
R17532 gnd.n4796 gnd.n4795 19.3944
R17533 gnd.n4795 gnd.n1412 19.3944
R17534 gnd.n4791 gnd.n1412 19.3944
R17535 gnd.n4791 gnd.n4790 19.3944
R17536 gnd.n4790 gnd.n4789 19.3944
R17537 gnd.n4789 gnd.n1417 19.3944
R17538 gnd.n4785 gnd.n1417 19.3944
R17539 gnd.n4785 gnd.n4784 19.3944
R17540 gnd.n4784 gnd.n4783 19.3944
R17541 gnd.n4783 gnd.n1422 19.3944
R17542 gnd.n4779 gnd.n1422 19.3944
R17543 gnd.n4779 gnd.n4778 19.3944
R17544 gnd.n4778 gnd.n4777 19.3944
R17545 gnd.n4777 gnd.n1427 19.3944
R17546 gnd.n4773 gnd.n1427 19.3944
R17547 gnd.n4773 gnd.n4772 19.3944
R17548 gnd.n4772 gnd.n4771 19.3944
R17549 gnd.n4771 gnd.n1432 19.3944
R17550 gnd.n4767 gnd.n1432 19.3944
R17551 gnd.n4767 gnd.n4766 19.3944
R17552 gnd.n4766 gnd.n4765 19.3944
R17553 gnd.n4765 gnd.n1437 19.3944
R17554 gnd.n4761 gnd.n1437 19.3944
R17555 gnd.n4761 gnd.n4760 19.3944
R17556 gnd.n4760 gnd.n4759 19.3944
R17557 gnd.n4759 gnd.n1442 19.3944
R17558 gnd.n4755 gnd.n1442 19.3944
R17559 gnd.n4755 gnd.n4754 19.3944
R17560 gnd.n4754 gnd.n4753 19.3944
R17561 gnd.n4753 gnd.n1447 19.3944
R17562 gnd.n4749 gnd.n1447 19.3944
R17563 gnd.n4749 gnd.n4748 19.3944
R17564 gnd.n4748 gnd.n4747 19.3944
R17565 gnd.n4747 gnd.n1452 19.3944
R17566 gnd.n4743 gnd.n1452 19.3944
R17567 gnd.n4743 gnd.n4742 19.3944
R17568 gnd.n4462 gnd.n4461 19.3944
R17569 gnd.n4461 gnd.n4460 19.3944
R17570 gnd.n4460 gnd.n1799 19.3944
R17571 gnd.n1701 gnd.n1697 19.3944
R17572 gnd.n1701 gnd.n1679 19.3944
R17573 gnd.n1714 gnd.n1679 19.3944
R17574 gnd.n1714 gnd.n1677 19.3944
R17575 gnd.n1720 gnd.n1677 19.3944
R17576 gnd.n1720 gnd.n1670 19.3944
R17577 gnd.n1733 gnd.n1670 19.3944
R17578 gnd.n1733 gnd.n1668 19.3944
R17579 gnd.n1739 gnd.n1668 19.3944
R17580 gnd.n1739 gnd.n1661 19.3944
R17581 gnd.n1752 gnd.n1661 19.3944
R17582 gnd.n1752 gnd.n1659 19.3944
R17583 gnd.n1758 gnd.n1659 19.3944
R17584 gnd.n1758 gnd.n1652 19.3944
R17585 gnd.n1771 gnd.n1652 19.3944
R17586 gnd.n1771 gnd.n1650 19.3944
R17587 gnd.n4474 gnd.n1650 19.3944
R17588 gnd.n4474 gnd.n4473 19.3944
R17589 gnd.n4473 gnd.n4472 19.3944
R17590 gnd.n4472 gnd.n1779 19.3944
R17591 gnd.n4468 gnd.n1779 19.3944
R17592 gnd.n4468 gnd.n4467 19.3944
R17593 gnd.n4467 gnd.n4466 19.3944
R17594 gnd.n4466 gnd.n1787 19.3944
R17595 gnd.n5898 gnd.t153 18.8012
R17596 gnd.n5937 gnd.t163 18.8012
R17597 gnd.n5741 gnd.n5483 18.4825
R17598 gnd.n2030 gnd.n1889 18.4247
R17599 gnd.n3495 gnd.n2544 18.4247
R17600 gnd.n2446 gnd.n2445 18.2639
R17601 gnd.n4299 gnd.n4298 18.2639
R17602 gnd.n7620 gnd.n7619 18.2308
R17603 gnd.n1767 gnd.n1647 18.2308
R17604 gnd.n2800 gnd.n2784 18.2308
R17605 gnd.n3051 gnd.n3043 18.2308
R17606 gnd.t154 gnd.n5425 18.1639
R17607 gnd.n5454 gnd.t156 17.5266
R17608 gnd.t41 gnd.n1077 17.5266
R17609 gnd.n7572 gnd.t85 17.5266
R17610 gnd.t150 gnd.n5401 16.8893
R17611 gnd.n3149 gnd.t80 16.8893
R17612 gnd.n7540 gnd.t82 16.8893
R17613 gnd.t231 gnd.n5510 16.2519
R17614 gnd.n5368 gnd.t144 16.2519
R17615 gnd.n3181 gnd.t37 16.2519
R17616 gnd.n7508 gnd.t25 16.2519
R17617 gnd.n3337 gnd.n3336 15.9333
R17618 gnd.n3340 gnd.n3337 15.9333
R17619 gnd.n3340 gnd.n3339 15.9333
R17620 gnd.n3339 gnd.n3338 15.9333
R17621 gnd.n3348 gnd.n2702 15.9333
R17622 gnd.n3351 gnd.n3348 15.9333
R17623 gnd.n3352 gnd.n3351 15.9333
R17624 gnd.n3353 gnd.n3352 15.9333
R17625 gnd.n3356 gnd.n3353 15.9333
R17626 gnd.n3356 gnd.n3355 15.9333
R17627 gnd.n3355 gnd.n3354 15.9333
R17628 gnd.n3354 gnd.n2696 15.9333
R17629 gnd.n3364 gnd.n2696 15.9333
R17630 gnd.n3368 gnd.n3367 15.9333
R17631 gnd.n3369 gnd.n3368 15.9333
R17632 gnd.n3372 gnd.n3369 15.9333
R17633 gnd.n3372 gnd.n3371 15.9333
R17634 gnd.n3371 gnd.n3370 15.9333
R17635 gnd.n3370 gnd.n2690 15.9333
R17636 gnd.n3380 gnd.n2690 15.9333
R17637 gnd.n3383 gnd.n3380 15.9333
R17638 gnd.n3385 gnd.n3384 15.9333
R17639 gnd.n3388 gnd.n3385 15.9333
R17640 gnd.n3388 gnd.n3387 15.9333
R17641 gnd.n3387 gnd.n3386 15.9333
R17642 gnd.n3386 gnd.n2684 15.9333
R17643 gnd.n3396 gnd.n2684 15.9333
R17644 gnd.n3399 gnd.n3396 15.9333
R17645 gnd.n3399 gnd.n3397 15.9333
R17646 gnd.n3564 gnd.n2387 15.9333
R17647 gnd.n2421 gnd.n2420 15.9333
R17648 gnd.n3573 gnd.n3572 15.9333
R17649 gnd.n3603 gnd.n3602 15.9333
R17650 gnd.n3666 gnd.n3665 15.9333
R17651 gnd.n3674 gnd.n2331 15.9333
R17652 gnd.n3699 gnd.n2303 15.9333
R17653 gnd.n3725 gnd.n2298 15.9333
R17654 gnd.n3733 gnd.n2291 15.9333
R17655 gnd.n3770 gnd.n2280 15.9333
R17656 gnd.n3782 gnd.n3780 15.9333
R17657 gnd.n3747 gnd.n2258 15.9333
R17658 gnd.n3843 gnd.n3842 15.9333
R17659 gnd.n3851 gnd.n2246 15.9333
R17660 gnd.n3869 gnd.n3868 15.9333
R17661 gnd.n3877 gnd.n2217 15.9333
R17662 gnd.n3902 gnd.n2209 15.9333
R17663 gnd.n3902 gnd.n2212 15.9333
R17664 gnd.n3910 gnd.n2203 15.9333
R17665 gnd.n3948 gnd.n2192 15.9333
R17666 gnd.n3959 gnd.n3958 15.9333
R17667 gnd.n3925 gnd.n2171 15.9333
R17668 gnd.n4005 gnd.n4004 15.9333
R17669 gnd.n4013 gnd.n2159 15.9333
R17670 gnd.n4030 gnd.n4029 15.9333
R17671 gnd.n4038 gnd.n2129 15.9333
R17672 gnd.n4090 gnd.n2123 15.9333
R17673 gnd.n4099 gnd.n4098 15.9333
R17674 gnd.n4130 gnd.n4129 15.9333
R17675 gnd.n4069 gnd.n2079 15.9333
R17676 gnd.n4169 gnd.n4168 15.9333
R17677 gnd.n4177 gnd.n2066 15.9333
R17678 gnd.n4370 gnd.n1852 15.9333
R17679 gnd.n1871 gnd.n1870 15.9333
R17680 gnd.n4380 gnd.n4379 15.9333
R17681 gnd.n4379 gnd.n4378 15.9333
R17682 gnd.n4378 gnd.n1841 15.9333
R17683 gnd.n4388 gnd.n1841 15.9333
R17684 gnd.n4390 gnd.n4388 15.9333
R17685 gnd.n4390 gnd.n4389 15.9333
R17686 gnd.n4389 gnd.n1834 15.9333
R17687 gnd.n4400 gnd.n1834 15.9333
R17688 gnd.n4399 gnd.n4398 15.9333
R17689 gnd.n4398 gnd.n1828 15.9333
R17690 gnd.n4408 gnd.n1828 15.9333
R17691 gnd.n4410 gnd.n4408 15.9333
R17692 gnd.n4410 gnd.n4409 15.9333
R17693 gnd.n4409 gnd.n1821 15.9333
R17694 gnd.n4420 gnd.n1821 15.9333
R17695 gnd.n4420 gnd.n4419 15.9333
R17696 gnd.n4418 gnd.n1815 15.9333
R17697 gnd.n4428 gnd.n1815 15.9333
R17698 gnd.n4430 gnd.n4428 15.9333
R17699 gnd.n4430 gnd.n4429 15.9333
R17700 gnd.n4429 gnd.n1808 15.9333
R17701 gnd.n4443 gnd.n1808 15.9333
R17702 gnd.n4443 gnd.n4442 15.9333
R17703 gnd.n4442 gnd.n4441 15.9333
R17704 gnd.n4441 gnd.n4440 15.9333
R17705 gnd.n4453 gnd.n4452 15.9333
R17706 gnd.n4453 gnd.n1456 15.9333
R17707 gnd.n4740 gnd.n1456 15.9333
R17708 gnd.n4740 gnd.n4739 15.9333
R17709 gnd.n6360 gnd.n6358 15.6674
R17710 gnd.n6328 gnd.n6326 15.6674
R17711 gnd.n6296 gnd.n6294 15.6674
R17712 gnd.n6265 gnd.n6263 15.6674
R17713 gnd.n6233 gnd.n6231 15.6674
R17714 gnd.n6201 gnd.n6199 15.6674
R17715 gnd.n6169 gnd.n6167 15.6674
R17716 gnd.n6138 gnd.n6136 15.6674
R17717 gnd.n5628 gnd.t231 15.6146
R17718 gnd.n6398 gnd.t187 15.6146
R17719 gnd.n6499 gnd.t206 15.6146
R17720 gnd.n3215 gnd.t123 15.6146
R17721 gnd.n4637 gnd.t73 15.6146
R17722 gnd.n2463 gnd.n2352 15.296
R17723 gnd.n4167 gnd.n2075 15.296
R17724 gnd.n4216 gnd.n4215 15.0827
R17725 gnd.n2433 gnd.n2428 15.0481
R17726 gnd.n4226 gnd.n4225 15.0481
R17727 gnd.n6064 gnd.t157 14.9773
R17728 gnd.n3247 gnd.t29 14.9773
R17729 gnd.t8 gnd.n1289 14.9773
R17730 gnd.n3582 gnd.t95 14.9773
R17731 gnd.t97 gnd.n4194 14.9773
R17732 gnd.n4538 gnd.t22 14.9773
R17733 gnd.n4599 gnd.t63 14.9773
R17734 gnd.n2381 gnd.n2370 14.6587
R17735 gnd.n2454 gnd.t300 14.6587
R17736 gnd.n3702 gnd.n3700 14.6587
R17737 gnd.n2116 gnd.n2115 14.6587
R17738 gnd.t294 gnd.n2089 14.6587
R17739 gnd.n4207 gnd.n4206 14.6587
R17740 gnd.t326 gnd.n6102 14.34
R17741 gnd.n6120 gnd.t155 14.34
R17742 gnd.n5039 gnd.t41 14.34
R17743 gnd.t29 gnd.n1247 14.34
R17744 gnd.n3272 gnd.t8 14.34
R17745 gnd.t22 gnd.n4537 14.34
R17746 gnd.n1583 gnd.t63 14.34
R17747 gnd.n211 gnd.t85 14.34
R17748 gnd.n3604 gnd.n2356 14.0214
R17749 gnd.n2330 gnd.t298 14.0214
R17750 gnd.n3783 gnd.n2272 14.0214
R17751 gnd.n2245 gnd.n2244 14.0214
R17752 gnd.n3960 gnd.n2184 14.0214
R17753 gnd.n2158 gnd.n2157 14.0214
R17754 gnd.n4131 gnd.t180 14.0214
R17755 gnd.t118 gnd.n5825 13.7027
R17756 gnd.t123 gnd.n1206 13.7027
R17757 gnd.t73 gnd.n280 13.7027
R17758 gnd.n117 gnd.n106 13.7027
R17759 gnd.n5710 gnd.n5706 13.5763
R17760 gnd.n6462 gnd.n5160 13.5763
R17761 gnd.n1991 gnd.n1979 13.5763
R17762 gnd.n7672 gnd.n7671 13.5763
R17763 gnd.n5065 gnd.n1055 13.5763
R17764 gnd.n3461 gnd.n2636 13.5763
R17765 gnd.n5742 gnd.n5741 13.384
R17766 gnd.n3591 gnd.t245 13.384
R17767 gnd.n2322 gnd.n2317 13.384
R17768 gnd.n3625 gnd.t17 13.384
R17769 gnd.n3769 gnd.n2282 13.384
R17770 gnd.n2237 gnd.n2232 13.384
R17771 gnd.n3947 gnd.n2195 13.384
R17772 gnd.n2150 gnd.n2144 13.384
R17773 gnd.n4047 gnd.t297 13.384
R17774 gnd.n4118 gnd.n2101 13.384
R17775 gnd.n2064 gnd.t238 13.384
R17776 gnd.n2056 gnd.n2051 13.384
R17777 gnd.n2444 gnd.n2425 13.1884
R17778 gnd.n2439 gnd.n2438 13.1884
R17779 gnd.n2438 gnd.n2437 13.1884
R17780 gnd.n4219 gnd.n4214 13.1884
R17781 gnd.n4220 gnd.n4219 13.1884
R17782 gnd.n2440 gnd.n2427 13.146
R17783 gnd.n2436 gnd.n2427 13.146
R17784 gnd.n4218 gnd.n4217 13.146
R17785 gnd.n4218 gnd.n4213 13.146
R17786 gnd.t37 gnd.n1169 13.0654
R17787 gnd.n7473 gnd.t25 13.0654
R17788 gnd.n6361 gnd.n6357 12.8005
R17789 gnd.n6329 gnd.n6325 12.8005
R17790 gnd.n6297 gnd.n6293 12.8005
R17791 gnd.n6266 gnd.n6262 12.8005
R17792 gnd.n6234 gnd.n6230 12.8005
R17793 gnd.n6202 gnd.n6198 12.8005
R17794 gnd.n6170 gnd.n6166 12.8005
R17795 gnd.n6139 gnd.n6135 12.8005
R17796 gnd.n3584 gnd.n3583 12.7467
R17797 gnd.n3689 gnd.n2309 12.7467
R17798 gnd.n3762 gnd.n3761 12.7467
R17799 gnd.n3866 gnd.n2224 12.7467
R17800 gnd.n3940 gnd.n3939 12.7467
R17801 gnd.n4028 gnd.n2136 12.7467
R17802 gnd.n4111 gnd.n4110 12.7467
R17803 gnd.t80 gnd.n1127 12.4281
R17804 gnd.n3367 gnd.t159 12.4281
R17805 gnd.n4419 gnd.t12 12.4281
R17806 gnd.n7458 gnd.t82 12.4281
R17807 gnd.n5713 gnd.n5710 12.4126
R17808 gnd.n6465 gnd.n6462 12.4126
R17809 gnd.n1987 gnd.n1979 12.4126
R17810 gnd.n7671 gnd.n179 12.4126
R17811 gnd.n5061 gnd.n1055 12.4126
R17812 gnd.n3456 gnd.n2636 12.4126
R17813 gnd.n3560 gnd.n2446 12.1761
R17814 gnd.n4298 gnd.n4297 12.1761
R17815 gnd.n3675 gnd.n2328 12.1094
R17816 gnd.n3790 gnd.n2266 12.1094
R17817 gnd.n3852 gnd.n2242 12.1094
R17818 gnd.n3967 gnd.n2179 12.1094
R17819 gnd.n4014 gnd.n2155 12.1094
R17820 gnd.n4138 gnd.n2087 12.1094
R17821 gnd.n4178 gnd.n2061 12.1094
R17822 gnd.n6365 gnd.n6364 12.0247
R17823 gnd.n6333 gnd.n6332 12.0247
R17824 gnd.n6301 gnd.n6300 12.0247
R17825 gnd.n6270 gnd.n6269 12.0247
R17826 gnd.n6238 gnd.n6237 12.0247
R17827 gnd.n6206 gnd.n6205 12.0247
R17828 gnd.n6174 gnd.n6173 12.0247
R17829 gnd.n6143 gnd.n6142 12.0247
R17830 gnd.n3718 gnd.n2304 11.4721
R17831 gnd.n3710 gnd.n3709 11.4721
R17832 gnd.n3895 gnd.n2218 11.4721
R17833 gnd.n3887 gnd.n3886 11.4721
R17834 gnd.n4056 gnd.n2130 11.4721
R17835 gnd.n4048 gnd.n2114 11.4721
R17836 gnd.t255 gnd.n2042 11.4721
R17837 gnd.n4301 gnd.n1852 11.4721
R17838 gnd.n6368 gnd.n6355 11.249
R17839 gnd.n6336 gnd.n6323 11.249
R17840 gnd.n6304 gnd.n6291 11.249
R17841 gnd.n6273 gnd.n6260 11.249
R17842 gnd.n6241 gnd.n6228 11.249
R17843 gnd.n6209 gnd.n6196 11.249
R17844 gnd.n6177 gnd.n6164 11.249
R17845 gnd.n6146 gnd.n6133 11.249
R17846 gnd.n5826 gnd.t118 11.1535
R17847 gnd.n3397 gnd.t55 11.1535
R17848 gnd.n4380 gnd.t161 11.1535
R17849 gnd.n3612 gnd.t276 10.8348
R17850 gnd.n3658 gnd.n3657 10.8348
R17851 gnd.n3734 gnd.t44 10.8348
R17852 gnd.n3834 gnd.n3833 10.8348
R17853 gnd.n3833 gnd.n2252 10.8348
R17854 gnd.n3997 gnd.n3996 10.8348
R17855 gnd.n3996 gnd.n2165 10.8348
R17856 gnd.t19 gnd.n4039 10.8348
R17857 gnd.n4160 gnd.n2072 10.8348
R17858 gnd.n4366 gnd.n4365 10.6151
R17859 gnd.n4365 gnd.n4362 10.6151
R17860 gnd.n4360 gnd.n4357 10.6151
R17861 gnd.n4357 gnd.n4356 10.6151
R17862 gnd.n4356 gnd.n4353 10.6151
R17863 gnd.n4353 gnd.n4352 10.6151
R17864 gnd.n4352 gnd.n4349 10.6151
R17865 gnd.n4349 gnd.n4348 10.6151
R17866 gnd.n4348 gnd.n4345 10.6151
R17867 gnd.n4345 gnd.n4344 10.6151
R17868 gnd.n4344 gnd.n4341 10.6151
R17869 gnd.n4341 gnd.n4340 10.6151
R17870 gnd.n4340 gnd.n4337 10.6151
R17871 gnd.n4337 gnd.n4336 10.6151
R17872 gnd.n4336 gnd.n4333 10.6151
R17873 gnd.n4333 gnd.n4332 10.6151
R17874 gnd.n4332 gnd.n4329 10.6151
R17875 gnd.n4329 gnd.n4328 10.6151
R17876 gnd.n4328 gnd.n4325 10.6151
R17877 gnd.n4325 gnd.n4324 10.6151
R17878 gnd.n4324 gnd.n4321 10.6151
R17879 gnd.n4321 gnd.n4320 10.6151
R17880 gnd.n4320 gnd.n4317 10.6151
R17881 gnd.n4317 gnd.n4316 10.6151
R17882 gnd.n4316 gnd.n4313 10.6151
R17883 gnd.n4313 gnd.n4312 10.6151
R17884 gnd.n4312 gnd.n4309 10.6151
R17885 gnd.n4309 gnd.n4308 10.6151
R17886 gnd.n4308 gnd.n4305 10.6151
R17887 gnd.n4305 gnd.n4304 10.6151
R17888 gnd.n2476 gnd.n2452 10.6151
R17889 gnd.n2476 gnd.n2475 10.6151
R17890 gnd.n2475 gnd.n2474 10.6151
R17891 gnd.n2474 gnd.n2473 10.6151
R17892 gnd.n2473 gnd.n2472 10.6151
R17893 gnd.n2472 gnd.n2469 10.6151
R17894 gnd.n2469 gnd.n2468 10.6151
R17895 gnd.n2468 gnd.n2466 10.6151
R17896 gnd.n2466 gnd.n2465 10.6151
R17897 gnd.n2465 gnd.n2461 10.6151
R17898 gnd.n2461 gnd.n2460 10.6151
R17899 gnd.n2460 gnd.n2458 10.6151
R17900 gnd.n2458 gnd.n2457 10.6151
R17901 gnd.n2457 gnd.n2453 10.6151
R17902 gnd.n2453 gnd.n2320 10.6151
R17903 gnd.n3684 gnd.n2320 10.6151
R17904 gnd.n3685 gnd.n3684 10.6151
R17905 gnd.n3687 gnd.n3685 10.6151
R17906 gnd.n3687 gnd.n3686 10.6151
R17907 gnd.n3686 gnd.n2301 10.6151
R17908 gnd.n3720 gnd.n2301 10.6151
R17909 gnd.n3721 gnd.n3720 10.6151
R17910 gnd.n3723 gnd.n3721 10.6151
R17911 gnd.n3723 gnd.n3722 10.6151
R17912 gnd.n3722 gnd.n2288 10.6151
R17913 gnd.n3736 gnd.n2288 10.6151
R17914 gnd.n3737 gnd.n3736 10.6151
R17915 gnd.n3759 gnd.n3737 10.6151
R17916 gnd.n3759 gnd.n3758 10.6151
R17917 gnd.n3758 gnd.n3757 10.6151
R17918 gnd.n3757 gnd.n3754 10.6151
R17919 gnd.n3754 gnd.n3753 10.6151
R17920 gnd.n3753 gnd.n3751 10.6151
R17921 gnd.n3751 gnd.n3750 10.6151
R17922 gnd.n3750 gnd.n3746 10.6151
R17923 gnd.n3746 gnd.n3745 10.6151
R17924 gnd.n3745 gnd.n3743 10.6151
R17925 gnd.n3743 gnd.n3742 10.6151
R17926 gnd.n3742 gnd.n3738 10.6151
R17927 gnd.n3738 gnd.n2235 10.6151
R17928 gnd.n3861 gnd.n2235 10.6151
R17929 gnd.n3862 gnd.n3861 10.6151
R17930 gnd.n3864 gnd.n3862 10.6151
R17931 gnd.n3864 gnd.n3863 10.6151
R17932 gnd.n3863 gnd.n2215 10.6151
R17933 gnd.n3897 gnd.n2215 10.6151
R17934 gnd.n3898 gnd.n3897 10.6151
R17935 gnd.n3900 gnd.n3898 10.6151
R17936 gnd.n3900 gnd.n3899 10.6151
R17937 gnd.n3899 gnd.n2201 10.6151
R17938 gnd.n3913 gnd.n2201 10.6151
R17939 gnd.n3914 gnd.n3913 10.6151
R17940 gnd.n3937 gnd.n3914 10.6151
R17941 gnd.n3937 gnd.n3936 10.6151
R17942 gnd.n3936 gnd.n3935 10.6151
R17943 gnd.n3935 gnd.n3932 10.6151
R17944 gnd.n3932 gnd.n3931 10.6151
R17945 gnd.n3931 gnd.n3929 10.6151
R17946 gnd.n3929 gnd.n3928 10.6151
R17947 gnd.n3928 gnd.n3923 10.6151
R17948 gnd.n3923 gnd.n3922 10.6151
R17949 gnd.n3922 gnd.n3920 10.6151
R17950 gnd.n3920 gnd.n3919 10.6151
R17951 gnd.n3919 gnd.n3915 10.6151
R17952 gnd.n3915 gnd.n2147 10.6151
R17953 gnd.n4023 gnd.n2147 10.6151
R17954 gnd.n4024 gnd.n4023 10.6151
R17955 gnd.n4026 gnd.n4024 10.6151
R17956 gnd.n4026 gnd.n4025 10.6151
R17957 gnd.n4025 gnd.n2127 10.6151
R17958 gnd.n4058 gnd.n2127 10.6151
R17959 gnd.n4059 gnd.n4058 10.6151
R17960 gnd.n4088 gnd.n4059 10.6151
R17961 gnd.n4088 gnd.n4087 10.6151
R17962 gnd.n4087 gnd.n4086 10.6151
R17963 gnd.n4086 gnd.n4083 10.6151
R17964 gnd.n4083 gnd.n4082 10.6151
R17965 gnd.n4082 gnd.n4081 10.6151
R17966 gnd.n4081 gnd.n4080 10.6151
R17967 gnd.n4080 gnd.n4079 10.6151
R17968 gnd.n4079 gnd.n4076 10.6151
R17969 gnd.n4076 gnd.n4075 10.6151
R17970 gnd.n4075 gnd.n4073 10.6151
R17971 gnd.n4073 gnd.n4072 10.6151
R17972 gnd.n4072 gnd.n4067 10.6151
R17973 gnd.n4067 gnd.n4066 10.6151
R17974 gnd.n4066 gnd.n4064 10.6151
R17975 gnd.n4064 gnd.n4063 10.6151
R17976 gnd.n4063 gnd.n4060 10.6151
R17977 gnd.n4060 gnd.n2054 10.6151
R17978 gnd.n4187 gnd.n2054 10.6151
R17979 gnd.n4188 gnd.n4187 10.6151
R17980 gnd.n4191 gnd.n4188 10.6151
R17981 gnd.n4191 gnd.n4190 10.6151
R17982 gnd.n4190 gnd.n4189 10.6151
R17983 gnd.n4189 gnd.n2034 10.6151
R17984 gnd.n2542 gnd.n2541 10.6151
R17985 gnd.n2541 gnd.n2538 10.6151
R17986 gnd.n2536 gnd.n2533 10.6151
R17987 gnd.n2533 gnd.n2532 10.6151
R17988 gnd.n2532 gnd.n2529 10.6151
R17989 gnd.n2529 gnd.n2528 10.6151
R17990 gnd.n2528 gnd.n2525 10.6151
R17991 gnd.n2525 gnd.n2524 10.6151
R17992 gnd.n2524 gnd.n2521 10.6151
R17993 gnd.n2521 gnd.n2520 10.6151
R17994 gnd.n2520 gnd.n2517 10.6151
R17995 gnd.n2517 gnd.n2516 10.6151
R17996 gnd.n2516 gnd.n2513 10.6151
R17997 gnd.n2513 gnd.n2512 10.6151
R17998 gnd.n2512 gnd.n2509 10.6151
R17999 gnd.n2509 gnd.n2508 10.6151
R18000 gnd.n2508 gnd.n2505 10.6151
R18001 gnd.n2505 gnd.n2504 10.6151
R18002 gnd.n2504 gnd.n2501 10.6151
R18003 gnd.n2501 gnd.n2500 10.6151
R18004 gnd.n2500 gnd.n2497 10.6151
R18005 gnd.n2497 gnd.n2496 10.6151
R18006 gnd.n2496 gnd.n2493 10.6151
R18007 gnd.n2493 gnd.n2492 10.6151
R18008 gnd.n2492 gnd.n2489 10.6151
R18009 gnd.n2489 gnd.n2488 10.6151
R18010 gnd.n2488 gnd.n2485 10.6151
R18011 gnd.n2485 gnd.n2484 10.6151
R18012 gnd.n2484 gnd.n2481 10.6151
R18013 gnd.n2481 gnd.n2480 10.6151
R18014 gnd.n3560 gnd.n3559 10.6151
R18015 gnd.n3559 gnd.n3558 10.6151
R18016 gnd.n3558 gnd.n3557 10.6151
R18017 gnd.n3557 gnd.n3555 10.6151
R18018 gnd.n3555 gnd.n3552 10.6151
R18019 gnd.n3552 gnd.n3551 10.6151
R18020 gnd.n3551 gnd.n3548 10.6151
R18021 gnd.n3548 gnd.n3547 10.6151
R18022 gnd.n3547 gnd.n3544 10.6151
R18023 gnd.n3544 gnd.n3543 10.6151
R18024 gnd.n3543 gnd.n3540 10.6151
R18025 gnd.n3540 gnd.n3539 10.6151
R18026 gnd.n3539 gnd.n3536 10.6151
R18027 gnd.n3536 gnd.n3535 10.6151
R18028 gnd.n3535 gnd.n3532 10.6151
R18029 gnd.n3532 gnd.n3531 10.6151
R18030 gnd.n3531 gnd.n3528 10.6151
R18031 gnd.n3528 gnd.n3527 10.6151
R18032 gnd.n3527 gnd.n3524 10.6151
R18033 gnd.n3524 gnd.n3523 10.6151
R18034 gnd.n3523 gnd.n3520 10.6151
R18035 gnd.n3520 gnd.n3519 10.6151
R18036 gnd.n3519 gnd.n3516 10.6151
R18037 gnd.n3516 gnd.n3515 10.6151
R18038 gnd.n3515 gnd.n3512 10.6151
R18039 gnd.n3512 gnd.n3511 10.6151
R18040 gnd.n3511 gnd.n3508 10.6151
R18041 gnd.n3508 gnd.n3507 10.6151
R18042 gnd.n3504 gnd.n3503 10.6151
R18043 gnd.n3503 gnd.n3500 10.6151
R18044 gnd.n4297 gnd.n4296 10.6151
R18045 gnd.n4296 gnd.n4293 10.6151
R18046 gnd.n4293 gnd.n4292 10.6151
R18047 gnd.n4292 gnd.n4289 10.6151
R18048 gnd.n4289 gnd.n4288 10.6151
R18049 gnd.n4288 gnd.n4285 10.6151
R18050 gnd.n4285 gnd.n4284 10.6151
R18051 gnd.n4284 gnd.n4281 10.6151
R18052 gnd.n4281 gnd.n4280 10.6151
R18053 gnd.n4280 gnd.n4277 10.6151
R18054 gnd.n4277 gnd.n4276 10.6151
R18055 gnd.n4276 gnd.n4273 10.6151
R18056 gnd.n4273 gnd.n4272 10.6151
R18057 gnd.n4272 gnd.n4269 10.6151
R18058 gnd.n4269 gnd.n4268 10.6151
R18059 gnd.n4268 gnd.n4265 10.6151
R18060 gnd.n4265 gnd.n4264 10.6151
R18061 gnd.n4264 gnd.n4261 10.6151
R18062 gnd.n4261 gnd.n4260 10.6151
R18063 gnd.n4260 gnd.n4257 10.6151
R18064 gnd.n4257 gnd.n4256 10.6151
R18065 gnd.n4256 gnd.n4253 10.6151
R18066 gnd.n4253 gnd.n4252 10.6151
R18067 gnd.n4252 gnd.n4249 10.6151
R18068 gnd.n4249 gnd.n4248 10.6151
R18069 gnd.n4248 gnd.n4245 10.6151
R18070 gnd.n4245 gnd.n4244 10.6151
R18071 gnd.n4244 gnd.n4241 10.6151
R18072 gnd.n4239 gnd.n4236 10.6151
R18073 gnd.n4236 gnd.n4235 10.6151
R18074 gnd.n2445 gnd.n2367 10.6151
R18075 gnd.n3587 gnd.n2367 10.6151
R18076 gnd.n3588 gnd.n3587 10.6151
R18077 gnd.n3589 gnd.n3588 10.6151
R18078 gnd.n3589 gnd.n2354 10.6151
R18079 gnd.n3606 gnd.n2354 10.6151
R18080 gnd.n3607 gnd.n3606 10.6151
R18081 gnd.n3608 gnd.n3607 10.6151
R18082 gnd.n3608 gnd.n2341 10.6151
R18083 gnd.n3660 gnd.n2341 10.6151
R18084 gnd.n3661 gnd.n3660 10.6151
R18085 gnd.n3662 gnd.n3661 10.6151
R18086 gnd.n3662 gnd.n2325 10.6151
R18087 gnd.n3677 gnd.n2325 10.6151
R18088 gnd.n3678 gnd.n3677 10.6151
R18089 gnd.n3680 gnd.n3678 10.6151
R18090 gnd.n3680 gnd.n3679 10.6151
R18091 gnd.n3679 gnd.n2307 10.6151
R18092 gnd.n3705 gnd.n2307 10.6151
R18093 gnd.n3706 gnd.n3705 10.6151
R18094 gnd.n3716 gnd.n3706 10.6151
R18095 gnd.n3716 gnd.n3715 10.6151
R18096 gnd.n3715 gnd.n3714 10.6151
R18097 gnd.n3714 gnd.n3713 10.6151
R18098 gnd.n3713 gnd.n3707 10.6151
R18099 gnd.n3707 gnd.n2284 10.6151
R18100 gnd.n3765 gnd.n2284 10.6151
R18101 gnd.n3766 gnd.n3765 10.6151
R18102 gnd.n3767 gnd.n3766 10.6151
R18103 gnd.n3767 gnd.n2270 10.6151
R18104 gnd.n3785 gnd.n2270 10.6151
R18105 gnd.n3786 gnd.n3785 10.6151
R18106 gnd.n3787 gnd.n3786 10.6151
R18107 gnd.n3787 gnd.n2256 10.6151
R18108 gnd.n3836 gnd.n2256 10.6151
R18109 gnd.n3837 gnd.n3836 10.6151
R18110 gnd.n3838 gnd.n3837 10.6151
R18111 gnd.n3838 gnd.n2240 10.6151
R18112 gnd.n3854 gnd.n2240 10.6151
R18113 gnd.n3855 gnd.n3854 10.6151
R18114 gnd.n3857 gnd.n3855 10.6151
R18115 gnd.n3857 gnd.n3856 10.6151
R18116 gnd.n3856 gnd.n2222 10.6151
R18117 gnd.n3882 gnd.n2222 10.6151
R18118 gnd.n3883 gnd.n3882 10.6151
R18119 gnd.n3893 gnd.n3883 10.6151
R18120 gnd.n3893 gnd.n3892 10.6151
R18121 gnd.n3892 gnd.n3891 10.6151
R18122 gnd.n3891 gnd.n3890 10.6151
R18123 gnd.n3890 gnd.n3884 10.6151
R18124 gnd.n3884 gnd.n2197 10.6151
R18125 gnd.n3943 gnd.n2197 10.6151
R18126 gnd.n3944 gnd.n3943 10.6151
R18127 gnd.n3945 gnd.n3944 10.6151
R18128 gnd.n3945 gnd.n2182 10.6151
R18129 gnd.n3962 gnd.n2182 10.6151
R18130 gnd.n3963 gnd.n3962 10.6151
R18131 gnd.n3964 gnd.n3963 10.6151
R18132 gnd.n3964 gnd.n2169 10.6151
R18133 gnd.n3999 gnd.n2169 10.6151
R18134 gnd.n4000 gnd.n3999 10.6151
R18135 gnd.n4001 gnd.n4000 10.6151
R18136 gnd.n4001 gnd.n2153 10.6151
R18137 gnd.n4016 gnd.n2153 10.6151
R18138 gnd.n4017 gnd.n4016 10.6151
R18139 gnd.n4019 gnd.n4017 10.6151
R18140 gnd.n4019 gnd.n4018 10.6151
R18141 gnd.n4018 gnd.n2134 10.6151
R18142 gnd.n4043 gnd.n2134 10.6151
R18143 gnd.n4044 gnd.n4043 10.6151
R18144 gnd.n4054 gnd.n4044 10.6151
R18145 gnd.n4054 gnd.n4053 10.6151
R18146 gnd.n4053 gnd.n4052 10.6151
R18147 gnd.n4052 gnd.n4051 10.6151
R18148 gnd.n4051 gnd.n4045 10.6151
R18149 gnd.n4045 gnd.n2103 10.6151
R18150 gnd.n4114 gnd.n2103 10.6151
R18151 gnd.n4115 gnd.n4114 10.6151
R18152 gnd.n4116 gnd.n4115 10.6151
R18153 gnd.n4116 gnd.n2091 10.6151
R18154 gnd.n4133 gnd.n2091 10.6151
R18155 gnd.n4134 gnd.n4133 10.6151
R18156 gnd.n4135 gnd.n4134 10.6151
R18157 gnd.n4135 gnd.n2077 10.6151
R18158 gnd.n4163 gnd.n2077 10.6151
R18159 gnd.n4164 gnd.n4163 10.6151
R18160 gnd.n4165 gnd.n4164 10.6151
R18161 gnd.n4165 gnd.n2059 10.6151
R18162 gnd.n4180 gnd.n2059 10.6151
R18163 gnd.n4181 gnd.n4180 10.6151
R18164 gnd.n4183 gnd.n4181 10.6151
R18165 gnd.n4183 gnd.n4182 10.6151
R18166 gnd.n4182 gnd.n2040 10.6151
R18167 gnd.n4210 gnd.n2040 10.6151
R18168 gnd.n4211 gnd.n4210 10.6151
R18169 gnd.n4299 gnd.n4211 10.6151
R18170 gnd.n5498 gnd.t0 10.5161
R18171 gnd.n6103 gnd.t326 10.5161
R18172 gnd.n6513 gnd.t155 10.5161
R18173 gnd.n6369 gnd.n6353 10.4732
R18174 gnd.n6337 gnd.n6321 10.4732
R18175 gnd.n6305 gnd.n6289 10.4732
R18176 gnd.n6274 gnd.n6258 10.4732
R18177 gnd.n6242 gnd.n6226 10.4732
R18178 gnd.n6210 gnd.n6194 10.4732
R18179 gnd.n6178 gnd.n6162 10.4732
R18180 gnd.n6147 gnd.n6131 10.4732
R18181 gnd.n2462 gnd.t225 10.1975
R18182 gnd.n3624 gnd.n2304 10.1975
R18183 gnd.n2220 gnd.n2218 10.1975
R18184 gnd.n3888 gnd.n3887 10.1975
R18185 gnd.n4049 gnd.n4048 10.1975
R18186 gnd.n6078 gnd.t157 9.87883
R18187 gnd.n3563 gnd.n2421 9.87883
R18188 gnd.n4370 gnd.n4369 9.87883
R18189 gnd.n7786 gnd.n66 9.73455
R18190 gnd.n6373 gnd.n6372 9.69747
R18191 gnd.n6341 gnd.n6340 9.69747
R18192 gnd.n6309 gnd.n6308 9.69747
R18193 gnd.n6278 gnd.n6277 9.69747
R18194 gnd.n6246 gnd.n6245 9.69747
R18195 gnd.n6214 gnd.n6213 9.69747
R18196 gnd.n6182 gnd.n6181 9.69747
R18197 gnd.n6151 gnd.n6150 9.69747
R18198 gnd.n3612 gnd.n3610 9.56018
R18199 gnd.n2455 gnd.n2328 9.56018
R18200 gnd.n3790 gnd.n3789 9.56018
R18201 gnd.t181 gnd.n2268 9.56018
R18202 gnd.n3740 gnd.n2242 9.56018
R18203 gnd.n3967 gnd.n3966 9.56018
R18204 gnd.n3916 gnd.t135 9.56018
R18205 gnd.n3917 gnd.n2155 9.56018
R18206 gnd.n4138 gnd.n4137 9.56018
R18207 gnd.n4205 gnd.t191 9.56018
R18208 gnd.n4896 gnd.n1326 9.45751
R18209 gnd.n1692 gnd.n1684 9.45599
R18210 gnd.n6379 gnd.n6378 9.45567
R18211 gnd.n6347 gnd.n6346 9.45567
R18212 gnd.n6315 gnd.n6314 9.45567
R18213 gnd.n6284 gnd.n6283 9.45567
R18214 gnd.n6252 gnd.n6251 9.45567
R18215 gnd.n6220 gnd.n6219 9.45567
R18216 gnd.n6188 gnd.n6187 9.45567
R18217 gnd.n6157 gnd.n6156 9.45567
R18218 gnd.n5342 gnd.n5341 9.39724
R18219 gnd.n6378 gnd.n6377 9.3005
R18220 gnd.n6351 gnd.n6350 9.3005
R18221 gnd.n6372 gnd.n6371 9.3005
R18222 gnd.n6370 gnd.n6369 9.3005
R18223 gnd.n6355 gnd.n6354 9.3005
R18224 gnd.n6364 gnd.n6363 9.3005
R18225 gnd.n6362 gnd.n6361 9.3005
R18226 gnd.n6346 gnd.n6345 9.3005
R18227 gnd.n6319 gnd.n6318 9.3005
R18228 gnd.n6340 gnd.n6339 9.3005
R18229 gnd.n6338 gnd.n6337 9.3005
R18230 gnd.n6323 gnd.n6322 9.3005
R18231 gnd.n6332 gnd.n6331 9.3005
R18232 gnd.n6330 gnd.n6329 9.3005
R18233 gnd.n6314 gnd.n6313 9.3005
R18234 gnd.n6287 gnd.n6286 9.3005
R18235 gnd.n6308 gnd.n6307 9.3005
R18236 gnd.n6306 gnd.n6305 9.3005
R18237 gnd.n6291 gnd.n6290 9.3005
R18238 gnd.n6300 gnd.n6299 9.3005
R18239 gnd.n6298 gnd.n6297 9.3005
R18240 gnd.n6283 gnd.n6282 9.3005
R18241 gnd.n6256 gnd.n6255 9.3005
R18242 gnd.n6277 gnd.n6276 9.3005
R18243 gnd.n6275 gnd.n6274 9.3005
R18244 gnd.n6260 gnd.n6259 9.3005
R18245 gnd.n6269 gnd.n6268 9.3005
R18246 gnd.n6267 gnd.n6266 9.3005
R18247 gnd.n6251 gnd.n6250 9.3005
R18248 gnd.n6224 gnd.n6223 9.3005
R18249 gnd.n6245 gnd.n6244 9.3005
R18250 gnd.n6243 gnd.n6242 9.3005
R18251 gnd.n6228 gnd.n6227 9.3005
R18252 gnd.n6237 gnd.n6236 9.3005
R18253 gnd.n6235 gnd.n6234 9.3005
R18254 gnd.n6219 gnd.n6218 9.3005
R18255 gnd.n6192 gnd.n6191 9.3005
R18256 gnd.n6213 gnd.n6212 9.3005
R18257 gnd.n6211 gnd.n6210 9.3005
R18258 gnd.n6196 gnd.n6195 9.3005
R18259 gnd.n6205 gnd.n6204 9.3005
R18260 gnd.n6203 gnd.n6202 9.3005
R18261 gnd.n6187 gnd.n6186 9.3005
R18262 gnd.n6160 gnd.n6159 9.3005
R18263 gnd.n6181 gnd.n6180 9.3005
R18264 gnd.n6179 gnd.n6178 9.3005
R18265 gnd.n6164 gnd.n6163 9.3005
R18266 gnd.n6173 gnd.n6172 9.3005
R18267 gnd.n6171 gnd.n6170 9.3005
R18268 gnd.n6156 gnd.n6155 9.3005
R18269 gnd.n6129 gnd.n6128 9.3005
R18270 gnd.n6150 gnd.n6149 9.3005
R18271 gnd.n6148 gnd.n6147 9.3005
R18272 gnd.n6133 gnd.n6132 9.3005
R18273 gnd.n6142 gnd.n6141 9.3005
R18274 gnd.n6140 gnd.n6139 9.3005
R18275 gnd.n964 gnd.n963 9.3005
R18276 gnd.n6487 gnd.n5147 9.3005
R18277 gnd.n6486 gnd.n5148 9.3005
R18278 gnd.n6485 gnd.n5149 9.3005
R18279 gnd.n6482 gnd.n5150 9.3005
R18280 gnd.n6481 gnd.n5151 9.3005
R18281 gnd.n6478 gnd.n5152 9.3005
R18282 gnd.n6477 gnd.n5153 9.3005
R18283 gnd.n6474 gnd.n5154 9.3005
R18284 gnd.n6473 gnd.n5155 9.3005
R18285 gnd.n6470 gnd.n5156 9.3005
R18286 gnd.n6469 gnd.n5157 9.3005
R18287 gnd.n6466 gnd.n5158 9.3005
R18288 gnd.n6465 gnd.n5159 9.3005
R18289 gnd.n6462 gnd.n6461 9.3005
R18290 gnd.n6460 gnd.n5160 9.3005
R18291 gnd.n6493 gnd.n6492 9.3005
R18292 gnd.n5765 gnd.n5764 9.3005
R18293 gnd.n5766 gnd.n5468 9.3005
R18294 gnd.n5768 gnd.n5767 9.3005
R18295 gnd.n5449 gnd.n5448 9.3005
R18296 gnd.n5795 gnd.n5794 9.3005
R18297 gnd.n5796 gnd.n5447 9.3005
R18298 gnd.n5800 gnd.n5797 9.3005
R18299 gnd.n5799 gnd.n5798 9.3005
R18300 gnd.n5423 gnd.n5422 9.3005
R18301 gnd.n5829 gnd.n5828 9.3005
R18302 gnd.n5830 gnd.n5421 9.3005
R18303 gnd.n5837 gnd.n5831 9.3005
R18304 gnd.n5836 gnd.n5832 9.3005
R18305 gnd.n5835 gnd.n5833 9.3005
R18306 gnd.n5390 gnd.n5389 9.3005
R18307 gnd.n5890 gnd.n5889 9.3005
R18308 gnd.n5891 gnd.n5388 9.3005
R18309 gnd.n5895 gnd.n5892 9.3005
R18310 gnd.n5894 gnd.n5893 9.3005
R18311 gnd.n5363 gnd.n5362 9.3005
R18312 gnd.n5930 gnd.n5929 9.3005
R18313 gnd.n5931 gnd.n5361 9.3005
R18314 gnd.n5935 gnd.n5932 9.3005
R18315 gnd.n5934 gnd.n5933 9.3005
R18316 gnd.n5288 gnd.n5287 9.3005
R18317 gnd.n5975 gnd.n5974 9.3005
R18318 gnd.n5976 gnd.n5286 9.3005
R18319 gnd.n5980 gnd.n5977 9.3005
R18320 gnd.n5979 gnd.n5978 9.3005
R18321 gnd.n5260 gnd.n5259 9.3005
R18322 gnd.n6014 gnd.n6013 9.3005
R18323 gnd.n6015 gnd.n5258 9.3005
R18324 gnd.n6022 gnd.n6016 9.3005
R18325 gnd.n6021 gnd.n6017 9.3005
R18326 gnd.n6020 gnd.n6018 9.3005
R18327 gnd.n5229 gnd.n5228 9.3005
R18328 gnd.n6069 gnd.n6068 9.3005
R18329 gnd.n6070 gnd.n5227 9.3005
R18330 gnd.n6075 gnd.n6071 9.3005
R18331 gnd.n6074 gnd.n6073 9.3005
R18332 gnd.n6072 gnd.n912 9.3005
R18333 gnd.n6524 gnd.n913 9.3005
R18334 gnd.n6523 gnd.n914 9.3005
R18335 gnd.n6522 gnd.n915 9.3005
R18336 gnd.n935 gnd.n916 9.3005
R18337 gnd.n936 gnd.n934 9.3005
R18338 gnd.n6510 gnd.n937 9.3005
R18339 gnd.n6509 gnd.n938 9.3005
R18340 gnd.n6508 gnd.n939 9.3005
R18341 gnd.n960 gnd.n940 9.3005
R18342 gnd.n961 gnd.n959 9.3005
R18343 gnd.n6496 gnd.n962 9.3005
R18344 gnd.n6495 gnd.n6494 9.3005
R18345 gnd.n5470 gnd.n5469 9.3005
R18346 gnd.n5710 gnd.n5709 9.3005
R18347 gnd.n5713 gnd.n5705 9.3005
R18348 gnd.n5714 gnd.n5704 9.3005
R18349 gnd.n5717 gnd.n5703 9.3005
R18350 gnd.n5718 gnd.n5702 9.3005
R18351 gnd.n5721 gnd.n5701 9.3005
R18352 gnd.n5722 gnd.n5700 9.3005
R18353 gnd.n5725 gnd.n5699 9.3005
R18354 gnd.n5726 gnd.n5698 9.3005
R18355 gnd.n5729 gnd.n5697 9.3005
R18356 gnd.n5730 gnd.n5696 9.3005
R18357 gnd.n5733 gnd.n5695 9.3005
R18358 gnd.n5735 gnd.n5694 9.3005
R18359 gnd.n5736 gnd.n5693 9.3005
R18360 gnd.n5737 gnd.n5692 9.3005
R18361 gnd.n5738 gnd.n5691 9.3005
R18362 gnd.n5706 gnd.n5487 9.3005
R18363 gnd.n5755 gnd.n5478 9.3005
R18364 gnd.n5757 gnd.n5756 9.3005
R18365 gnd.n5465 gnd.n5460 9.3005
R18366 gnd.n5778 gnd.n5459 9.3005
R18367 gnd.n5781 gnd.n5780 9.3005
R18368 gnd.n5783 gnd.n5782 9.3005
R18369 gnd.n5786 gnd.n5442 9.3005
R18370 gnd.n5784 gnd.n5440 9.3005
R18371 gnd.n5806 gnd.n5438 9.3005
R18372 gnd.n5810 gnd.n5809 9.3005
R18373 gnd.n5808 gnd.n5413 9.3005
R18374 gnd.n5844 gnd.n5412 9.3005
R18375 gnd.n5847 gnd.n5846 9.3005
R18376 gnd.n5410 gnd.n5409 9.3005
R18377 gnd.n5853 gnd.n5407 9.3005
R18378 gnd.n5855 gnd.n5854 9.3005
R18379 gnd.n5381 gnd.n5380 9.3005
R18380 gnd.n5904 gnd.n5903 9.3005
R18381 gnd.n5905 gnd.n5374 9.3005
R18382 gnd.n5913 gnd.n5373 9.3005
R18383 gnd.n5916 gnd.n5915 9.3005
R18384 gnd.n5918 gnd.n5917 9.3005
R18385 gnd.n5921 gnd.n5356 9.3005
R18386 gnd.n5919 gnd.n5354 9.3005
R18387 gnd.n5941 gnd.n5352 9.3005
R18388 gnd.n5943 gnd.n5942 9.3005
R18389 gnd.n5278 gnd.n5277 9.3005
R18390 gnd.n5989 gnd.n5988 9.3005
R18391 gnd.n5990 gnd.n5271 9.3005
R18392 gnd.n5998 gnd.n5270 9.3005
R18393 gnd.n6001 gnd.n6000 9.3005
R18394 gnd.n6003 gnd.n6002 9.3005
R18395 gnd.n6005 gnd.n5253 9.3005
R18396 gnd.n5250 gnd.n5248 9.3005
R18397 gnd.n6030 gnd.n6029 9.3005
R18398 gnd.n5251 gnd.n5234 9.3005
R18399 gnd.n6058 gnd.n5233 9.3005
R18400 gnd.n6062 gnd.n6060 9.3005
R18401 gnd.n6061 gnd.n5218 9.3005
R18402 gnd.n6083 gnd.n5217 9.3005
R18403 gnd.n6087 gnd.n6086 9.3005
R18404 gnd.n5210 gnd.n5209 9.3005
R18405 gnd.n6100 gnd.n6096 9.3005
R18406 gnd.n6099 gnd.n6098 9.3005
R18407 gnd.n5202 gnd.n5201 9.3005
R18408 gnd.n6122 gnd.n5203 9.3005
R18409 gnd.n6124 gnd.n6123 9.3005
R18410 gnd.n6126 gnd.n5200 9.3005
R18411 gnd.n6385 gnd.n6384 9.3005
R18412 gnd.n6387 gnd.n6386 9.3005
R18413 gnd.n6395 gnd.n6388 9.3005
R18414 gnd.n6394 gnd.n6390 9.3005
R18415 gnd.n6393 gnd.n5163 9.3005
R18416 gnd.n5754 gnd.n5481 9.3005
R18417 gnd.n6456 gnd.n5164 9.3005
R18418 gnd.n6455 gnd.n5166 9.3005
R18419 gnd.n6452 gnd.n5167 9.3005
R18420 gnd.n6451 gnd.n5168 9.3005
R18421 gnd.n6448 gnd.n5169 9.3005
R18422 gnd.n6447 gnd.n5170 9.3005
R18423 gnd.n6444 gnd.n5171 9.3005
R18424 gnd.n6443 gnd.n5172 9.3005
R18425 gnd.n6440 gnd.n5173 9.3005
R18426 gnd.n6439 gnd.n5174 9.3005
R18427 gnd.n6436 gnd.n5175 9.3005
R18428 gnd.n6435 gnd.n5176 9.3005
R18429 gnd.n6432 gnd.n5177 9.3005
R18430 gnd.n6431 gnd.n5178 9.3005
R18431 gnd.n6428 gnd.n5179 9.3005
R18432 gnd.n6427 gnd.n5180 9.3005
R18433 gnd.n6424 gnd.n5181 9.3005
R18434 gnd.n6423 gnd.n5182 9.3005
R18435 gnd.n6420 gnd.n5183 9.3005
R18436 gnd.n6419 gnd.n5184 9.3005
R18437 gnd.n6416 gnd.n5185 9.3005
R18438 gnd.n6415 gnd.n5186 9.3005
R18439 gnd.n6412 gnd.n5190 9.3005
R18440 gnd.n6411 gnd.n5191 9.3005
R18441 gnd.n6408 gnd.n5192 9.3005
R18442 gnd.n6407 gnd.n5193 9.3005
R18443 gnd.n6458 gnd.n6457 9.3005
R18444 gnd.n5951 gnd.n5950 9.3005
R18445 gnd.n5952 gnd.n5294 9.3005
R18446 gnd.n5969 gnd.n5953 9.3005
R18447 gnd.n5968 gnd.n5954 9.3005
R18448 gnd.n5967 gnd.n5955 9.3005
R18449 gnd.n5965 gnd.n5956 9.3005
R18450 gnd.n5964 gnd.n5957 9.3005
R18451 gnd.n5962 gnd.n5958 9.3005
R18452 gnd.n5961 gnd.n5959 9.3005
R18453 gnd.n5241 gnd.n5240 9.3005
R18454 gnd.n6037 gnd.n6036 9.3005
R18455 gnd.n6038 gnd.n5239 9.3005
R18456 gnd.n6052 gnd.n6039 9.3005
R18457 gnd.n6051 gnd.n6040 9.3005
R18458 gnd.n6050 gnd.n6041 9.3005
R18459 gnd.n6049 gnd.n6042 9.3005
R18460 gnd.n6047 gnd.n6043 9.3005
R18461 gnd.n6046 gnd.n6044 9.3005
R18462 gnd.n5207 gnd.n5206 9.3005
R18463 gnd.n6106 gnd.n6105 9.3005
R18464 gnd.n6107 gnd.n5205 9.3005
R18465 gnd.n6117 gnd.n6108 9.3005
R18466 gnd.n6116 gnd.n6109 9.3005
R18467 gnd.n6115 gnd.n6110 9.3005
R18468 gnd.n6112 gnd.n6111 9.3005
R18469 gnd.n5196 gnd.n5195 9.3005
R18470 gnd.n6401 gnd.n6400 9.3005
R18471 gnd.n6402 gnd.n5194 9.3005
R18472 gnd.n6404 gnd.n6403 9.3005
R18473 gnd.n5624 gnd.n5518 9.3005
R18474 gnd.n5626 gnd.n5625 9.3005
R18475 gnd.n5508 gnd.n5507 9.3005
R18476 gnd.n5639 gnd.n5638 9.3005
R18477 gnd.n5640 gnd.n5506 9.3005
R18478 gnd.n5642 gnd.n5641 9.3005
R18479 gnd.n5495 gnd.n5494 9.3005
R18480 gnd.n5655 gnd.n5654 9.3005
R18481 gnd.n5656 gnd.n5493 9.3005
R18482 gnd.n5680 gnd.n5657 9.3005
R18483 gnd.n5679 gnd.n5658 9.3005
R18484 gnd.n5678 gnd.n5659 9.3005
R18485 gnd.n5677 gnd.n5660 9.3005
R18486 gnd.n5675 gnd.n5661 9.3005
R18487 gnd.n5674 gnd.n5662 9.3005
R18488 gnd.n5672 gnd.n5663 9.3005
R18489 gnd.n5671 gnd.n5664 9.3005
R18490 gnd.n5669 gnd.n5665 9.3005
R18491 gnd.n5668 gnd.n5666 9.3005
R18492 gnd.n5430 gnd.n5429 9.3005
R18493 gnd.n5818 gnd.n5817 9.3005
R18494 gnd.n5819 gnd.n5428 9.3005
R18495 gnd.n5823 gnd.n5820 9.3005
R18496 gnd.n5822 gnd.n5821 9.3005
R18497 gnd.n5397 gnd.n5396 9.3005
R18498 gnd.n5865 gnd.n5864 9.3005
R18499 gnd.n5866 gnd.n5395 9.3005
R18500 gnd.n5868 gnd.n5867 9.3005
R18501 gnd.n5623 gnd.n5622 9.3005
R18502 gnd.n5563 gnd.n5562 9.3005
R18503 gnd.n5568 gnd.n5560 9.3005
R18504 gnd.n5569 gnd.n5559 9.3005
R18505 gnd.n5571 gnd.n5556 9.3005
R18506 gnd.n5555 gnd.n5553 9.3005
R18507 gnd.n5577 gnd.n5552 9.3005
R18508 gnd.n5578 gnd.n5551 9.3005
R18509 gnd.n5579 gnd.n5550 9.3005
R18510 gnd.n5549 gnd.n5547 9.3005
R18511 gnd.n5585 gnd.n5546 9.3005
R18512 gnd.n5586 gnd.n5545 9.3005
R18513 gnd.n5587 gnd.n5544 9.3005
R18514 gnd.n5543 gnd.n5541 9.3005
R18515 gnd.n5593 gnd.n5540 9.3005
R18516 gnd.n5594 gnd.n5539 9.3005
R18517 gnd.n5595 gnd.n5538 9.3005
R18518 gnd.n5537 gnd.n5535 9.3005
R18519 gnd.n5601 gnd.n5534 9.3005
R18520 gnd.n5602 gnd.n5533 9.3005
R18521 gnd.n5603 gnd.n5532 9.3005
R18522 gnd.n5531 gnd.n5529 9.3005
R18523 gnd.n5608 gnd.n5528 9.3005
R18524 gnd.n5609 gnd.n5527 9.3005
R18525 gnd.n5526 gnd.n5524 9.3005
R18526 gnd.n5614 gnd.n5523 9.3005
R18527 gnd.n5616 gnd.n5615 9.3005
R18528 gnd.n5561 gnd.n5519 9.3005
R18529 gnd.n5514 gnd.n5513 9.3005
R18530 gnd.n5631 gnd.n5630 9.3005
R18531 gnd.n5632 gnd.n5512 9.3005
R18532 gnd.n5634 gnd.n5633 9.3005
R18533 gnd.n5502 gnd.n5501 9.3005
R18534 gnd.n5647 gnd.n5646 9.3005
R18535 gnd.n5648 gnd.n5500 9.3005
R18536 gnd.n5650 gnd.n5649 9.3005
R18537 gnd.n5489 gnd.n5488 9.3005
R18538 gnd.n5745 gnd.n5744 9.3005
R18539 gnd.n5747 gnd.n5486 9.3005
R18540 gnd.n5749 gnd.n5748 9.3005
R18541 gnd.n5480 gnd.n5477 9.3005
R18542 gnd.n5759 gnd.n5758 9.3005
R18543 gnd.n5479 gnd.n5461 9.3005
R18544 gnd.n5777 gnd.n5776 9.3005
R18545 gnd.n5779 gnd.n5457 9.3005
R18546 gnd.n5789 gnd.n5458 9.3005
R18547 gnd.n5788 gnd.n5787 9.3005
R18548 gnd.n5785 gnd.n5436 9.3005
R18549 gnd.n5813 gnd.n5437 9.3005
R18550 gnd.n5812 gnd.n5811 9.3005
R18551 gnd.n5439 gnd.n5414 9.3005
R18552 gnd.n5843 gnd.n5842 9.3005
R18553 gnd.n5845 gnd.n5404 9.3005
R18554 gnd.n5860 gnd.n5405 9.3005
R18555 gnd.n5859 gnd.n5406 9.3005
R18556 gnd.n5858 gnd.n5856 9.3005
R18557 gnd.n5408 gnd.n5382 9.3005
R18558 gnd.n5901 gnd.n5900 9.3005
R18559 gnd.n5902 gnd.n5375 9.3005
R18560 gnd.n5912 gnd.n5911 9.3005
R18561 gnd.n5914 gnd.n5371 9.3005
R18562 gnd.n5924 gnd.n5372 9.3005
R18563 gnd.n5923 gnd.n5922 9.3005
R18564 gnd.n5920 gnd.n5350 9.3005
R18565 gnd.n5946 gnd.n5351 9.3005
R18566 gnd.n5945 gnd.n5944 9.3005
R18567 gnd.n5353 gnd.n5279 9.3005
R18568 gnd.n5986 gnd.n5985 9.3005
R18569 gnd.n5987 gnd.n5272 9.3005
R18570 gnd.n5997 gnd.n5996 9.3005
R18571 gnd.n5999 gnd.n5268 9.3005
R18572 gnd.n6008 gnd.n5269 9.3005
R18573 gnd.n6007 gnd.n6006 9.3005
R18574 gnd.n6004 gnd.n5247 9.3005
R18575 gnd.n6032 gnd.n6031 9.3005
R18576 gnd.n5249 gnd.n5235 9.3005
R18577 gnd.n6057 gnd.n6056 9.3005
R18578 gnd.n6059 gnd.n5219 9.3005
R18579 gnd.n6080 gnd.n5220 9.3005
R18580 gnd.n6082 gnd.n6081 9.3005
R18581 gnd.n6084 gnd.n5213 9.3005
R18582 gnd.n6085 gnd.n5211 9.3005
R18583 gnd.n6095 gnd.n6094 9.3005
R18584 gnd.n6097 gnd.n923 9.3005
R18585 gnd.n6517 gnd.n924 9.3005
R18586 gnd.n6516 gnd.n925 9.3005
R18587 gnd.n6515 gnd.n926 9.3005
R18588 gnd.n6125 gnd.n927 9.3005
R18589 gnd.n6383 gnd.n948 9.3005
R18590 gnd.n6503 gnd.n949 9.3005
R18591 gnd.n6502 gnd.n950 9.3005
R18592 gnd.n6501 gnd.n951 9.3005
R18593 gnd.n6389 gnd.n952 9.3005
R18594 gnd.n5618 gnd.n5617 9.3005
R18595 gnd.n738 gnd.n737 9.3005
R18596 gnd.n6700 gnd.n6699 9.3005
R18597 gnd.n6701 gnd.n736 9.3005
R18598 gnd.n6703 gnd.n6702 9.3005
R18599 gnd.n732 gnd.n731 9.3005
R18600 gnd.n6710 gnd.n6709 9.3005
R18601 gnd.n6711 gnd.n730 9.3005
R18602 gnd.n6713 gnd.n6712 9.3005
R18603 gnd.n726 gnd.n725 9.3005
R18604 gnd.n6720 gnd.n6719 9.3005
R18605 gnd.n6721 gnd.n724 9.3005
R18606 gnd.n6723 gnd.n6722 9.3005
R18607 gnd.n720 gnd.n719 9.3005
R18608 gnd.n6730 gnd.n6729 9.3005
R18609 gnd.n6731 gnd.n718 9.3005
R18610 gnd.n6733 gnd.n6732 9.3005
R18611 gnd.n714 gnd.n713 9.3005
R18612 gnd.n6740 gnd.n6739 9.3005
R18613 gnd.n6741 gnd.n712 9.3005
R18614 gnd.n6743 gnd.n6742 9.3005
R18615 gnd.n708 gnd.n707 9.3005
R18616 gnd.n6750 gnd.n6749 9.3005
R18617 gnd.n6751 gnd.n706 9.3005
R18618 gnd.n6753 gnd.n6752 9.3005
R18619 gnd.n702 gnd.n701 9.3005
R18620 gnd.n6760 gnd.n6759 9.3005
R18621 gnd.n6761 gnd.n700 9.3005
R18622 gnd.n6763 gnd.n6762 9.3005
R18623 gnd.n696 gnd.n695 9.3005
R18624 gnd.n6770 gnd.n6769 9.3005
R18625 gnd.n6771 gnd.n694 9.3005
R18626 gnd.n6773 gnd.n6772 9.3005
R18627 gnd.n690 gnd.n689 9.3005
R18628 gnd.n6780 gnd.n6779 9.3005
R18629 gnd.n6781 gnd.n688 9.3005
R18630 gnd.n6783 gnd.n6782 9.3005
R18631 gnd.n684 gnd.n683 9.3005
R18632 gnd.n6790 gnd.n6789 9.3005
R18633 gnd.n6791 gnd.n682 9.3005
R18634 gnd.n6793 gnd.n6792 9.3005
R18635 gnd.n678 gnd.n677 9.3005
R18636 gnd.n6800 gnd.n6799 9.3005
R18637 gnd.n6801 gnd.n676 9.3005
R18638 gnd.n6803 gnd.n6802 9.3005
R18639 gnd.n672 gnd.n671 9.3005
R18640 gnd.n6810 gnd.n6809 9.3005
R18641 gnd.n6811 gnd.n670 9.3005
R18642 gnd.n6813 gnd.n6812 9.3005
R18643 gnd.n666 gnd.n665 9.3005
R18644 gnd.n6820 gnd.n6819 9.3005
R18645 gnd.n6821 gnd.n664 9.3005
R18646 gnd.n6823 gnd.n6822 9.3005
R18647 gnd.n660 gnd.n659 9.3005
R18648 gnd.n6830 gnd.n6829 9.3005
R18649 gnd.n6831 gnd.n658 9.3005
R18650 gnd.n6833 gnd.n6832 9.3005
R18651 gnd.n654 gnd.n653 9.3005
R18652 gnd.n6840 gnd.n6839 9.3005
R18653 gnd.n6841 gnd.n652 9.3005
R18654 gnd.n6843 gnd.n6842 9.3005
R18655 gnd.n648 gnd.n647 9.3005
R18656 gnd.n6850 gnd.n6849 9.3005
R18657 gnd.n6851 gnd.n646 9.3005
R18658 gnd.n6853 gnd.n6852 9.3005
R18659 gnd.n642 gnd.n641 9.3005
R18660 gnd.n6860 gnd.n6859 9.3005
R18661 gnd.n6861 gnd.n640 9.3005
R18662 gnd.n6863 gnd.n6862 9.3005
R18663 gnd.n636 gnd.n635 9.3005
R18664 gnd.n6870 gnd.n6869 9.3005
R18665 gnd.n6871 gnd.n634 9.3005
R18666 gnd.n6873 gnd.n6872 9.3005
R18667 gnd.n630 gnd.n629 9.3005
R18668 gnd.n6880 gnd.n6879 9.3005
R18669 gnd.n6881 gnd.n628 9.3005
R18670 gnd.n6883 gnd.n6882 9.3005
R18671 gnd.n624 gnd.n623 9.3005
R18672 gnd.n6890 gnd.n6889 9.3005
R18673 gnd.n6891 gnd.n622 9.3005
R18674 gnd.n6893 gnd.n6892 9.3005
R18675 gnd.n618 gnd.n617 9.3005
R18676 gnd.n6900 gnd.n6899 9.3005
R18677 gnd.n6901 gnd.n616 9.3005
R18678 gnd.n6903 gnd.n6902 9.3005
R18679 gnd.n612 gnd.n611 9.3005
R18680 gnd.n6910 gnd.n6909 9.3005
R18681 gnd.n6911 gnd.n610 9.3005
R18682 gnd.n6913 gnd.n6912 9.3005
R18683 gnd.n606 gnd.n605 9.3005
R18684 gnd.n6920 gnd.n6919 9.3005
R18685 gnd.n6921 gnd.n604 9.3005
R18686 gnd.n6923 gnd.n6922 9.3005
R18687 gnd.n600 gnd.n599 9.3005
R18688 gnd.n6930 gnd.n6929 9.3005
R18689 gnd.n6931 gnd.n598 9.3005
R18690 gnd.n6933 gnd.n6932 9.3005
R18691 gnd.n594 gnd.n593 9.3005
R18692 gnd.n6940 gnd.n6939 9.3005
R18693 gnd.n6941 gnd.n592 9.3005
R18694 gnd.n6943 gnd.n6942 9.3005
R18695 gnd.n588 gnd.n587 9.3005
R18696 gnd.n6950 gnd.n6949 9.3005
R18697 gnd.n6951 gnd.n586 9.3005
R18698 gnd.n6953 gnd.n6952 9.3005
R18699 gnd.n582 gnd.n581 9.3005
R18700 gnd.n6960 gnd.n6959 9.3005
R18701 gnd.n6961 gnd.n580 9.3005
R18702 gnd.n6963 gnd.n6962 9.3005
R18703 gnd.n576 gnd.n575 9.3005
R18704 gnd.n6970 gnd.n6969 9.3005
R18705 gnd.n6971 gnd.n574 9.3005
R18706 gnd.n6973 gnd.n6972 9.3005
R18707 gnd.n570 gnd.n569 9.3005
R18708 gnd.n6980 gnd.n6979 9.3005
R18709 gnd.n6981 gnd.n568 9.3005
R18710 gnd.n6983 gnd.n6982 9.3005
R18711 gnd.n564 gnd.n563 9.3005
R18712 gnd.n6990 gnd.n6989 9.3005
R18713 gnd.n6991 gnd.n562 9.3005
R18714 gnd.n6993 gnd.n6992 9.3005
R18715 gnd.n558 gnd.n557 9.3005
R18716 gnd.n7000 gnd.n6999 9.3005
R18717 gnd.n7001 gnd.n556 9.3005
R18718 gnd.n7003 gnd.n7002 9.3005
R18719 gnd.n552 gnd.n551 9.3005
R18720 gnd.n7010 gnd.n7009 9.3005
R18721 gnd.n7011 gnd.n550 9.3005
R18722 gnd.n7013 gnd.n7012 9.3005
R18723 gnd.n546 gnd.n545 9.3005
R18724 gnd.n7020 gnd.n7019 9.3005
R18725 gnd.n7021 gnd.n544 9.3005
R18726 gnd.n7023 gnd.n7022 9.3005
R18727 gnd.n540 gnd.n539 9.3005
R18728 gnd.n7030 gnd.n7029 9.3005
R18729 gnd.n7031 gnd.n538 9.3005
R18730 gnd.n7033 gnd.n7032 9.3005
R18731 gnd.n534 gnd.n533 9.3005
R18732 gnd.n7040 gnd.n7039 9.3005
R18733 gnd.n7041 gnd.n532 9.3005
R18734 gnd.n7043 gnd.n7042 9.3005
R18735 gnd.n528 gnd.n527 9.3005
R18736 gnd.n7050 gnd.n7049 9.3005
R18737 gnd.n7051 gnd.n526 9.3005
R18738 gnd.n7053 gnd.n7052 9.3005
R18739 gnd.n522 gnd.n521 9.3005
R18740 gnd.n7060 gnd.n7059 9.3005
R18741 gnd.n7061 gnd.n520 9.3005
R18742 gnd.n7063 gnd.n7062 9.3005
R18743 gnd.n516 gnd.n515 9.3005
R18744 gnd.n7070 gnd.n7069 9.3005
R18745 gnd.n7071 gnd.n514 9.3005
R18746 gnd.n7073 gnd.n7072 9.3005
R18747 gnd.n510 gnd.n509 9.3005
R18748 gnd.n7080 gnd.n7079 9.3005
R18749 gnd.n7081 gnd.n508 9.3005
R18750 gnd.n7083 gnd.n7082 9.3005
R18751 gnd.n504 gnd.n503 9.3005
R18752 gnd.n7090 gnd.n7089 9.3005
R18753 gnd.n7091 gnd.n502 9.3005
R18754 gnd.n7093 gnd.n7092 9.3005
R18755 gnd.n498 gnd.n497 9.3005
R18756 gnd.n7100 gnd.n7099 9.3005
R18757 gnd.n7101 gnd.n496 9.3005
R18758 gnd.n7103 gnd.n7102 9.3005
R18759 gnd.n492 gnd.n491 9.3005
R18760 gnd.n7110 gnd.n7109 9.3005
R18761 gnd.n7111 gnd.n490 9.3005
R18762 gnd.n7113 gnd.n7112 9.3005
R18763 gnd.n486 gnd.n485 9.3005
R18764 gnd.n7120 gnd.n7119 9.3005
R18765 gnd.n7121 gnd.n484 9.3005
R18766 gnd.n7123 gnd.n7122 9.3005
R18767 gnd.n480 gnd.n479 9.3005
R18768 gnd.n7130 gnd.n7129 9.3005
R18769 gnd.n7131 gnd.n478 9.3005
R18770 gnd.n7133 gnd.n7132 9.3005
R18771 gnd.n474 gnd.n473 9.3005
R18772 gnd.n7140 gnd.n7139 9.3005
R18773 gnd.n7141 gnd.n472 9.3005
R18774 gnd.n7143 gnd.n7142 9.3005
R18775 gnd.n468 gnd.n467 9.3005
R18776 gnd.n7150 gnd.n7149 9.3005
R18777 gnd.n7151 gnd.n466 9.3005
R18778 gnd.n7153 gnd.n7152 9.3005
R18779 gnd.n462 gnd.n461 9.3005
R18780 gnd.n7160 gnd.n7159 9.3005
R18781 gnd.n7161 gnd.n460 9.3005
R18782 gnd.n7163 gnd.n7162 9.3005
R18783 gnd.n456 gnd.n455 9.3005
R18784 gnd.n7170 gnd.n7169 9.3005
R18785 gnd.n7171 gnd.n454 9.3005
R18786 gnd.n7174 gnd.n7173 9.3005
R18787 gnd.n7172 gnd.n450 9.3005
R18788 gnd.n7180 gnd.n449 9.3005
R18789 gnd.n7182 gnd.n7181 9.3005
R18790 gnd.n445 gnd.n444 9.3005
R18791 gnd.n7191 gnd.n7190 9.3005
R18792 gnd.n7192 gnd.n443 9.3005
R18793 gnd.n7194 gnd.n7193 9.3005
R18794 gnd.n439 gnd.n438 9.3005
R18795 gnd.n7201 gnd.n7200 9.3005
R18796 gnd.n7202 gnd.n437 9.3005
R18797 gnd.n7204 gnd.n7203 9.3005
R18798 gnd.n433 gnd.n432 9.3005
R18799 gnd.n7211 gnd.n7210 9.3005
R18800 gnd.n7212 gnd.n431 9.3005
R18801 gnd.n7214 gnd.n7213 9.3005
R18802 gnd.n427 gnd.n426 9.3005
R18803 gnd.n7221 gnd.n7220 9.3005
R18804 gnd.n7222 gnd.n425 9.3005
R18805 gnd.n7224 gnd.n7223 9.3005
R18806 gnd.n421 gnd.n420 9.3005
R18807 gnd.n7231 gnd.n7230 9.3005
R18808 gnd.n7232 gnd.n419 9.3005
R18809 gnd.n7234 gnd.n7233 9.3005
R18810 gnd.n415 gnd.n414 9.3005
R18811 gnd.n7241 gnd.n7240 9.3005
R18812 gnd.n7242 gnd.n413 9.3005
R18813 gnd.n7244 gnd.n7243 9.3005
R18814 gnd.n409 gnd.n408 9.3005
R18815 gnd.n7251 gnd.n7250 9.3005
R18816 gnd.n7252 gnd.n407 9.3005
R18817 gnd.n7254 gnd.n7253 9.3005
R18818 gnd.n403 gnd.n402 9.3005
R18819 gnd.n7261 gnd.n7260 9.3005
R18820 gnd.n7262 gnd.n401 9.3005
R18821 gnd.n7264 gnd.n7263 9.3005
R18822 gnd.n397 gnd.n396 9.3005
R18823 gnd.n7271 gnd.n7270 9.3005
R18824 gnd.n7272 gnd.n395 9.3005
R18825 gnd.n7274 gnd.n7273 9.3005
R18826 gnd.n391 gnd.n390 9.3005
R18827 gnd.n7281 gnd.n7280 9.3005
R18828 gnd.n7282 gnd.n389 9.3005
R18829 gnd.n7284 gnd.n7283 9.3005
R18830 gnd.n385 gnd.n384 9.3005
R18831 gnd.n7291 gnd.n7290 9.3005
R18832 gnd.n7292 gnd.n383 9.3005
R18833 gnd.n7294 gnd.n7293 9.3005
R18834 gnd.n379 gnd.n378 9.3005
R18835 gnd.n7301 gnd.n7300 9.3005
R18836 gnd.n7302 gnd.n377 9.3005
R18837 gnd.n7304 gnd.n7303 9.3005
R18838 gnd.n373 gnd.n372 9.3005
R18839 gnd.n7311 gnd.n7310 9.3005
R18840 gnd.n7312 gnd.n371 9.3005
R18841 gnd.n7314 gnd.n7313 9.3005
R18842 gnd.n367 gnd.n366 9.3005
R18843 gnd.n7321 gnd.n7320 9.3005
R18844 gnd.n7322 gnd.n365 9.3005
R18845 gnd.n7324 gnd.n7323 9.3005
R18846 gnd.n361 gnd.n360 9.3005
R18847 gnd.n7331 gnd.n7330 9.3005
R18848 gnd.n7332 gnd.n359 9.3005
R18849 gnd.n7334 gnd.n7333 9.3005
R18850 gnd.n355 gnd.n354 9.3005
R18851 gnd.n7341 gnd.n7340 9.3005
R18852 gnd.n7342 gnd.n353 9.3005
R18853 gnd.n7344 gnd.n7343 9.3005
R18854 gnd.n349 gnd.n348 9.3005
R18855 gnd.n7351 gnd.n7350 9.3005
R18856 gnd.n7352 gnd.n347 9.3005
R18857 gnd.n7354 gnd.n7353 9.3005
R18858 gnd.n343 gnd.n342 9.3005
R18859 gnd.n7361 gnd.n7360 9.3005
R18860 gnd.n7362 gnd.n341 9.3005
R18861 gnd.n7364 gnd.n7363 9.3005
R18862 gnd.n337 gnd.n336 9.3005
R18863 gnd.n7371 gnd.n7370 9.3005
R18864 gnd.n7372 gnd.n335 9.3005
R18865 gnd.n7374 gnd.n7373 9.3005
R18866 gnd.n331 gnd.n330 9.3005
R18867 gnd.n7381 gnd.n7380 9.3005
R18868 gnd.n7382 gnd.n329 9.3005
R18869 gnd.n7384 gnd.n7383 9.3005
R18870 gnd.n325 gnd.n324 9.3005
R18871 gnd.n7392 gnd.n7391 9.3005
R18872 gnd.n7393 gnd.n323 9.3005
R18873 gnd.n7395 gnd.n7394 9.3005
R18874 gnd.n7184 gnd.n7183 9.3005
R18875 gnd.n7737 gnd.n112 9.3005
R18876 gnd.n7736 gnd.n114 9.3005
R18877 gnd.n119 gnd.n115 9.3005
R18878 gnd.n7731 gnd.n120 9.3005
R18879 gnd.n7730 gnd.n121 9.3005
R18880 gnd.n7729 gnd.n122 9.3005
R18881 gnd.n126 gnd.n123 9.3005
R18882 gnd.n7724 gnd.n127 9.3005
R18883 gnd.n7723 gnd.n128 9.3005
R18884 gnd.n7722 gnd.n129 9.3005
R18885 gnd.n133 gnd.n130 9.3005
R18886 gnd.n7717 gnd.n134 9.3005
R18887 gnd.n7716 gnd.n135 9.3005
R18888 gnd.n7715 gnd.n136 9.3005
R18889 gnd.n140 gnd.n137 9.3005
R18890 gnd.n7710 gnd.n141 9.3005
R18891 gnd.n7709 gnd.n142 9.3005
R18892 gnd.n7705 gnd.n143 9.3005
R18893 gnd.n147 gnd.n144 9.3005
R18894 gnd.n7700 gnd.n148 9.3005
R18895 gnd.n7699 gnd.n149 9.3005
R18896 gnd.n7698 gnd.n150 9.3005
R18897 gnd.n154 gnd.n151 9.3005
R18898 gnd.n7693 gnd.n155 9.3005
R18899 gnd.n7692 gnd.n156 9.3005
R18900 gnd.n7691 gnd.n157 9.3005
R18901 gnd.n161 gnd.n158 9.3005
R18902 gnd.n7686 gnd.n162 9.3005
R18903 gnd.n7685 gnd.n163 9.3005
R18904 gnd.n7684 gnd.n164 9.3005
R18905 gnd.n168 gnd.n165 9.3005
R18906 gnd.n7679 gnd.n169 9.3005
R18907 gnd.n7678 gnd.n170 9.3005
R18908 gnd.n7677 gnd.n171 9.3005
R18909 gnd.n175 gnd.n172 9.3005
R18910 gnd.n7672 gnd.n176 9.3005
R18911 gnd.n7671 gnd.n7670 9.3005
R18912 gnd.n7669 gnd.n179 9.3005
R18913 gnd.n7739 gnd.n7738 9.3005
R18914 gnd.n1981 gnd.n1640 9.3005
R18915 gnd.n4489 gnd.n1639 9.3005
R18916 gnd.n4491 gnd.n4490 9.3005
R18917 gnd.n4492 gnd.n1638 9.3005
R18918 gnd.n4518 gnd.n4493 9.3005
R18919 gnd.n4517 gnd.n4494 9.3005
R18920 gnd.n4516 gnd.n4495 9.3005
R18921 gnd.n4515 gnd.n4496 9.3005
R18922 gnd.n4514 gnd.n4497 9.3005
R18923 gnd.n4512 gnd.n4498 9.3005
R18924 gnd.n4511 gnd.n4499 9.3005
R18925 gnd.n4509 gnd.n4500 9.3005
R18926 gnd.n4508 gnd.n4501 9.3005
R18927 gnd.n4507 gnd.n4502 9.3005
R18928 gnd.n4505 gnd.n4504 9.3005
R18929 gnd.n4503 gnd.n1558 9.3005
R18930 gnd.n4614 gnd.n1559 9.3005
R18931 gnd.n4615 gnd.n1557 9.3005
R18932 gnd.n4618 gnd.n4617 9.3005
R18933 gnd.n4619 gnd.n1556 9.3005
R18934 gnd.n4623 gnd.n4620 9.3005
R18935 gnd.n4622 gnd.n4621 9.3005
R18936 gnd.n1550 gnd.n1549 9.3005
R18937 gnd.n4641 gnd.n4640 9.3005
R18938 gnd.n4642 gnd.n1548 9.3005
R18939 gnd.n4644 gnd.n4643 9.3005
R18940 gnd.n300 gnd.n299 9.3005
R18941 gnd.n7478 gnd.n301 9.3005
R18942 gnd.n7477 gnd.n302 9.3005
R18943 gnd.n7476 gnd.n303 9.3005
R18944 gnd.n7405 gnd.n304 9.3005
R18945 gnd.n7409 gnd.n7408 9.3005
R18946 gnd.n7410 gnd.n7404 9.3005
R18947 gnd.n7415 gnd.n7411 9.3005
R18948 gnd.n7416 gnd.n7403 9.3005
R18949 gnd.n7420 gnd.n7419 9.3005
R18950 gnd.n7421 gnd.n7402 9.3005
R18951 gnd.n7454 gnd.n7422 9.3005
R18952 gnd.n7453 gnd.n7423 9.3005
R18953 gnd.n7452 gnd.n7424 9.3005
R18954 gnd.n7449 gnd.n7425 9.3005
R18955 gnd.n7448 gnd.n7426 9.3005
R18956 gnd.n7446 gnd.n7427 9.3005
R18957 gnd.n7445 gnd.n7428 9.3005
R18958 gnd.n7443 gnd.n7429 9.3005
R18959 gnd.n7442 gnd.n7430 9.3005
R18960 gnd.n7440 gnd.n7431 9.3005
R18961 gnd.n7439 gnd.n7432 9.3005
R18962 gnd.n7437 gnd.n7433 9.3005
R18963 gnd.n7436 gnd.n7435 9.3005
R18964 gnd.n7434 gnd.n183 9.3005
R18965 gnd.n7666 gnd.n182 9.3005
R18966 gnd.n7668 gnd.n7667 9.3005
R18967 gnd.n1983 gnd.n1982 9.3005
R18968 gnd.n1991 gnd.n1990 9.3005
R18969 gnd.n1980 gnd.n1975 9.3005
R18970 gnd.n1997 gnd.n1974 9.3005
R18971 gnd.n1998 gnd.n1973 9.3005
R18972 gnd.n1999 gnd.n1972 9.3005
R18973 gnd.n1971 gnd.n1969 9.3005
R18974 gnd.n2005 gnd.n1968 9.3005
R18975 gnd.n2006 gnd.n1967 9.3005
R18976 gnd.n2007 gnd.n1966 9.3005
R18977 gnd.n1965 gnd.n1963 9.3005
R18978 gnd.n2013 gnd.n1962 9.3005
R18979 gnd.n2014 gnd.n1961 9.3005
R18980 gnd.n2015 gnd.n1960 9.3005
R18981 gnd.n1959 gnd.n1957 9.3005
R18982 gnd.n2021 gnd.n1956 9.3005
R18983 gnd.n2022 gnd.n1955 9.3005
R18984 gnd.n2023 gnd.n1954 9.3005
R18985 gnd.n1953 gnd.n1951 9.3005
R18986 gnd.n2029 gnd.n1950 9.3005
R18987 gnd.n1946 gnd.n1889 9.3005
R18988 gnd.n1945 gnd.n1944 9.3005
R18989 gnd.n1892 gnd.n1891 9.3005
R18990 gnd.n1935 gnd.n1895 9.3005
R18991 gnd.n1937 gnd.n1936 9.3005
R18992 gnd.n1934 gnd.n1897 9.3005
R18993 gnd.n1933 gnd.n1932 9.3005
R18994 gnd.n1899 gnd.n1898 9.3005
R18995 gnd.n1926 gnd.n1925 9.3005
R18996 gnd.n1924 gnd.n1901 9.3005
R18997 gnd.n1923 gnd.n1922 9.3005
R18998 gnd.n1903 gnd.n1902 9.3005
R18999 gnd.n1916 gnd.n1915 9.3005
R19000 gnd.n1914 gnd.n1905 9.3005
R19001 gnd.n1913 gnd.n1912 9.3005
R19002 gnd.n1908 gnd.n1907 9.3005
R19003 gnd.n1989 gnd.n1979 9.3005
R19004 gnd.n1988 gnd.n1987 9.3005
R19005 gnd.n4722 gnd.n1485 9.3005
R19006 gnd.n4721 gnd.n1486 9.3005
R19007 gnd.n4720 gnd.n1487 9.3005
R19008 gnd.n4522 gnd.n1488 9.3005
R19009 gnd.n4526 gnd.n4523 9.3005
R19010 gnd.n4525 gnd.n4524 9.3005
R19011 gnd.n1603 gnd.n1602 9.3005
R19012 gnd.n4553 gnd.n4552 9.3005
R19013 gnd.n4554 gnd.n1601 9.3005
R19014 gnd.n4558 gnd.n4555 9.3005
R19015 gnd.n4557 gnd.n4556 9.3005
R19016 gnd.n1576 gnd.n1575 9.3005
R19017 gnd.n4592 gnd.n4591 9.3005
R19018 gnd.n4593 gnd.n1574 9.3005
R19019 gnd.n4597 gnd.n4594 9.3005
R19020 gnd.n4596 gnd.n4595 9.3005
R19021 gnd.n1524 gnd.n1523 9.3005
R19022 gnd.n4682 gnd.n4681 9.3005
R19023 gnd.n4683 gnd.n1522 9.3005
R19024 gnd.n4685 gnd.n4684 9.3005
R19025 gnd.n274 gnd.n267 9.3005
R19026 gnd.n253 gnd.n252 9.3005
R19027 gnd.n7519 gnd.n7518 9.3005
R19028 gnd.n7520 gnd.n251 9.3005
R19029 gnd.n7522 gnd.n7521 9.3005
R19030 gnd.n237 gnd.n236 9.3005
R19031 gnd.n7535 gnd.n7534 9.3005
R19032 gnd.n7536 gnd.n235 9.3005
R19033 gnd.n7538 gnd.n7537 9.3005
R19034 gnd.n223 gnd.n222 9.3005
R19035 gnd.n7551 gnd.n7550 9.3005
R19036 gnd.n7552 gnd.n221 9.3005
R19037 gnd.n7554 gnd.n7553 9.3005
R19038 gnd.n206 gnd.n205 9.3005
R19039 gnd.n7567 gnd.n7566 9.3005
R19040 gnd.n7568 gnd.n204 9.3005
R19041 gnd.n7570 gnd.n7569 9.3005
R19042 gnd.n191 gnd.n190 9.3005
R19043 gnd.n7658 gnd.n7657 9.3005
R19044 gnd.n7659 gnd.n189 9.3005
R19045 gnd.n7661 gnd.n7660 9.3005
R19046 gnd.n111 gnd.n110 9.3005
R19047 gnd.n7741 gnd.n7740 9.3005
R19048 gnd.n1906 gnd.n1484 9.3005
R19049 gnd.n7505 gnd.n272 9.3005
R19050 gnd.n7506 gnd.n7505 9.3005
R19051 gnd.n2977 gnd.n2941 9.3005
R19052 gnd.n2976 gnd.n2947 9.3005
R19053 gnd.n2950 gnd.n2948 9.3005
R19054 gnd.n2972 gnd.n2951 9.3005
R19055 gnd.n2971 gnd.n2952 9.3005
R19056 gnd.n2970 gnd.n2953 9.3005
R19057 gnd.n2956 gnd.n2954 9.3005
R19058 gnd.n2966 gnd.n2957 9.3005
R19059 gnd.n2965 gnd.n2958 9.3005
R19060 gnd.n2964 gnd.n2959 9.3005
R19061 gnd.n2961 gnd.n2960 9.3005
R19062 gnd.n2856 gnd.n2855 9.3005
R19063 gnd.n3303 gnd.n3302 9.3005
R19064 gnd.n3304 gnd.n2854 9.3005
R19065 gnd.n3306 gnd.n3305 9.3005
R19066 gnd.n2852 gnd.n2851 9.3005
R19067 gnd.n3311 gnd.n3310 9.3005
R19068 gnd.n3312 gnd.n2850 9.3005
R19069 gnd.n3314 gnd.n3313 9.3005
R19070 gnd.n2848 gnd.n2847 9.3005
R19071 gnd.n3319 gnd.n3318 9.3005
R19072 gnd.n3320 gnd.n2846 9.3005
R19073 gnd.n3322 gnd.n3321 9.3005
R19074 gnd.n2844 gnd.n2843 9.3005
R19075 gnd.n3330 gnd.n3329 9.3005
R19076 gnd.n3331 gnd.n2842 9.3005
R19077 gnd.n3333 gnd.n3332 9.3005
R19078 gnd.n2706 gnd.n2705 9.3005
R19079 gnd.n3343 gnd.n3342 9.3005
R19080 gnd.n3344 gnd.n2704 9.3005
R19081 gnd.n3346 gnd.n3345 9.3005
R19082 gnd.n2700 gnd.n2699 9.3005
R19083 gnd.n3359 gnd.n3358 9.3005
R19084 gnd.n3360 gnd.n2698 9.3005
R19085 gnd.n3362 gnd.n3361 9.3005
R19086 gnd.n2694 gnd.n2693 9.3005
R19087 gnd.n3375 gnd.n3374 9.3005
R19088 gnd.n3376 gnd.n2692 9.3005
R19089 gnd.n3378 gnd.n3377 9.3005
R19090 gnd.n2688 gnd.n2687 9.3005
R19091 gnd.n3391 gnd.n3390 9.3005
R19092 gnd.n3392 gnd.n2686 9.3005
R19093 gnd.n3394 gnd.n3393 9.3005
R19094 gnd.n2385 gnd.n2384 9.3005
R19095 gnd.n3567 gnd.n3566 9.3005
R19096 gnd.n3568 gnd.n2383 9.3005
R19097 gnd.n3570 gnd.n3569 9.3005
R19098 gnd.n2363 gnd.n2362 9.3005
R19099 gnd.n3595 gnd.n3594 9.3005
R19100 gnd.n3596 gnd.n2361 9.3005
R19101 gnd.n3600 gnd.n3597 9.3005
R19102 gnd.n3599 gnd.n3598 9.3005
R19103 gnd.n2335 gnd.n2334 9.3005
R19104 gnd.n3669 gnd.n3668 9.3005
R19105 gnd.n3670 gnd.n2333 9.3005
R19106 gnd.n3672 gnd.n3671 9.3005
R19107 gnd.n2315 gnd.n2314 9.3005
R19108 gnd.n3694 gnd.n3693 9.3005
R19109 gnd.n3695 gnd.n2313 9.3005
R19110 gnd.n3697 gnd.n3696 9.3005
R19111 gnd.n2295 gnd.n2294 9.3005
R19112 gnd.n3728 gnd.n3727 9.3005
R19113 gnd.n3729 gnd.n2293 9.3005
R19114 gnd.n3731 gnd.n3730 9.3005
R19115 gnd.n2278 gnd.n2277 9.3005
R19116 gnd.n3773 gnd.n3772 9.3005
R19117 gnd.n3774 gnd.n2276 9.3005
R19118 gnd.n3778 gnd.n3775 9.3005
R19119 gnd.n3777 gnd.n3776 9.3005
R19120 gnd.n2250 gnd.n2249 9.3005
R19121 gnd.n3846 gnd.n3845 9.3005
R19122 gnd.n3847 gnd.n2248 9.3005
R19123 gnd.n3849 gnd.n3848 9.3005
R19124 gnd.n2230 gnd.n2229 9.3005
R19125 gnd.n3872 gnd.n3871 9.3005
R19126 gnd.n3873 gnd.n2228 9.3005
R19127 gnd.n3875 gnd.n3874 9.3005
R19128 gnd.n2207 gnd.n2206 9.3005
R19129 gnd.n3905 gnd.n3904 9.3005
R19130 gnd.n3906 gnd.n2205 9.3005
R19131 gnd.n3908 gnd.n3907 9.3005
R19132 gnd.n2190 gnd.n2189 9.3005
R19133 gnd.n3951 gnd.n3950 9.3005
R19134 gnd.n3952 gnd.n2188 9.3005
R19135 gnd.n3956 gnd.n3953 9.3005
R19136 gnd.n3955 gnd.n3954 9.3005
R19137 gnd.n2163 gnd.n2162 9.3005
R19138 gnd.n4008 gnd.n4007 9.3005
R19139 gnd.n4009 gnd.n2161 9.3005
R19140 gnd.n4011 gnd.n4010 9.3005
R19141 gnd.n2142 gnd.n2141 9.3005
R19142 gnd.n4033 gnd.n4032 9.3005
R19143 gnd.n4034 gnd.n2140 9.3005
R19144 gnd.n4036 gnd.n4035 9.3005
R19145 gnd.n2120 gnd.n2119 9.3005
R19146 gnd.n4093 gnd.n4092 9.3005
R19147 gnd.n4094 gnd.n2118 9.3005
R19148 gnd.n4096 gnd.n4095 9.3005
R19149 gnd.n2098 gnd.n2097 9.3005
R19150 gnd.n4122 gnd.n4121 9.3005
R19151 gnd.n4123 gnd.n2096 9.3005
R19152 gnd.n4127 gnd.n4124 9.3005
R19153 gnd.n4126 gnd.n4125 9.3005
R19154 gnd.n2070 gnd.n2069 9.3005
R19155 gnd.n4172 gnd.n4171 9.3005
R19156 gnd.n4173 gnd.n2068 9.3005
R19157 gnd.n4175 gnd.n4174 9.3005
R19158 gnd.n2049 gnd.n2048 9.3005
R19159 gnd.n4198 gnd.n4197 9.3005
R19160 gnd.n4199 gnd.n2047 9.3005
R19161 gnd.n4203 gnd.n4200 9.3005
R19162 gnd.n4202 gnd.n4201 9.3005
R19163 gnd.n1845 gnd.n1844 9.3005
R19164 gnd.n4383 gnd.n4382 9.3005
R19165 gnd.n4384 gnd.n1843 9.3005
R19166 gnd.n4386 gnd.n4385 9.3005
R19167 gnd.n1832 gnd.n1831 9.3005
R19168 gnd.n4403 gnd.n4402 9.3005
R19169 gnd.n4404 gnd.n1830 9.3005
R19170 gnd.n4406 gnd.n4405 9.3005
R19171 gnd.n1819 gnd.n1818 9.3005
R19172 gnd.n4423 gnd.n4422 9.3005
R19173 gnd.n4424 gnd.n1817 9.3005
R19174 gnd.n4426 gnd.n4425 9.3005
R19175 gnd.n1806 gnd.n1805 9.3005
R19176 gnd.n4446 gnd.n4445 9.3005
R19177 gnd.n4447 gnd.n1804 9.3005
R19178 gnd.n4450 gnd.n4449 9.3005
R19179 gnd.n4448 gnd.n1461 9.3005
R19180 gnd.n4737 gnd.n1462 9.3005
R19181 gnd.n4736 gnd.n1463 9.3005
R19182 gnd.n4735 gnd.n1464 9.3005
R19183 gnd.n1470 gnd.n1465 9.3005
R19184 gnd.n4729 gnd.n1471 9.3005
R19185 gnd.n4728 gnd.n1472 9.3005
R19186 gnd.n4727 gnd.n1473 9.3005
R19187 gnd.n1626 gnd.n1474 9.3005
R19188 gnd.n1629 gnd.n1628 9.3005
R19189 gnd.n1630 gnd.n1625 9.3005
R19190 gnd.n1632 gnd.n1631 9.3005
R19191 gnd.n1614 gnd.n1613 9.3005
R19192 gnd.n4541 gnd.n4540 9.3005
R19193 gnd.n4542 gnd.n1612 9.3005
R19194 gnd.n4546 gnd.n4543 9.3005
R19195 gnd.n4545 gnd.n4544 9.3005
R19196 gnd.n1587 gnd.n1586 9.3005
R19197 gnd.n4574 gnd.n4573 9.3005
R19198 gnd.n4575 gnd.n1585 9.3005
R19199 gnd.n4586 gnd.n4576 9.3005
R19200 gnd.n4585 gnd.n4577 9.3005
R19201 gnd.n4584 gnd.n4578 9.3005
R19202 gnd.n4581 gnd.n4580 9.3005
R19203 gnd.n4579 gnd.n1532 9.3005
R19204 gnd.n4676 gnd.n1533 9.3005
R19205 gnd.n4675 gnd.n1534 9.3005
R19206 gnd.n4674 gnd.n1535 9.3005
R19207 gnd.n1537 gnd.n1536 9.3005
R19208 gnd.n7468 gnd.n309 9.3005
R19209 gnd.n312 gnd.n310 9.3005
R19210 gnd.n7464 gnd.n313 9.3005
R19211 gnd.n7463 gnd.n314 9.3005
R19212 gnd.n7462 gnd.n315 9.3005
R19213 gnd.n318 gnd.n316 9.3005
R19214 gnd.n7401 gnd.n319 9.3005
R19215 gnd.n7400 gnd.n320 9.3005
R19216 gnd.n7399 gnd.n321 9.3005
R19217 gnd.n2548 gnd.n2544 9.3005
R19218 gnd.n2581 gnd.n2578 9.3005
R19219 gnd.n2582 gnd.n2577 9.3005
R19220 gnd.n2585 gnd.n2576 9.3005
R19221 gnd.n2586 gnd.n2575 9.3005
R19222 gnd.n2589 gnd.n2574 9.3005
R19223 gnd.n2590 gnd.n2573 9.3005
R19224 gnd.n2593 gnd.n2572 9.3005
R19225 gnd.n2594 gnd.n2571 9.3005
R19226 gnd.n2597 gnd.n2570 9.3005
R19227 gnd.n2598 gnd.n2569 9.3005
R19228 gnd.n2601 gnd.n2568 9.3005
R19229 gnd.n2602 gnd.n2567 9.3005
R19230 gnd.n2603 gnd.n2566 9.3005
R19231 gnd.n2565 gnd.n2562 9.3005
R19232 gnd.n2564 gnd.n2563 9.3005
R19233 gnd.n3492 gnd.n3491 9.3005
R19234 gnd.n2550 gnd.n2549 9.3005
R19235 gnd.n2609 gnd.n2607 9.3005
R19236 gnd.n3484 gnd.n2610 9.3005
R19237 gnd.n3483 gnd.n2611 9.3005
R19238 gnd.n3482 gnd.n2612 9.3005
R19239 gnd.n2616 gnd.n2613 9.3005
R19240 gnd.n3477 gnd.n2617 9.3005
R19241 gnd.n3476 gnd.n2618 9.3005
R19242 gnd.n3475 gnd.n2619 9.3005
R19243 gnd.n2623 gnd.n2620 9.3005
R19244 gnd.n3470 gnd.n2624 9.3005
R19245 gnd.n3469 gnd.n2625 9.3005
R19246 gnd.n3468 gnd.n2626 9.3005
R19247 gnd.n2630 gnd.n2627 9.3005
R19248 gnd.n3463 gnd.n2631 9.3005
R19249 gnd.n3462 gnd.n2632 9.3005
R19250 gnd.n3461 gnd.n2633 9.3005
R19251 gnd.n2638 gnd.n2636 9.3005
R19252 gnd.n3456 gnd.n3455 9.3005
R19253 gnd.n3493 gnd.n2543 9.3005
R19254 gnd.n3044 gnd.n3018 9.3005
R19255 gnd.n3103 gnd.n3019 9.3005
R19256 gnd.n3104 gnd.n3017 9.3005
R19257 gnd.n3107 gnd.n3106 9.3005
R19258 gnd.n3108 gnd.n3016 9.3005
R19259 gnd.n3111 gnd.n3109 9.3005
R19260 gnd.n3112 gnd.n3015 9.3005
R19261 gnd.n3115 gnd.n3114 9.3005
R19262 gnd.n3116 gnd.n3014 9.3005
R19263 gnd.n3119 gnd.n3117 9.3005
R19264 gnd.n3120 gnd.n3013 9.3005
R19265 gnd.n3144 gnd.n3143 9.3005
R19266 gnd.n3145 gnd.n3012 9.3005
R19267 gnd.n3147 gnd.n3146 9.3005
R19268 gnd.n3008 gnd.n3007 9.3005
R19269 gnd.n3160 gnd.n3159 9.3005
R19270 gnd.n3161 gnd.n3006 9.3005
R19271 gnd.n3163 gnd.n3162 9.3005
R19272 gnd.n2910 gnd.n2909 9.3005
R19273 gnd.n3176 gnd.n3175 9.3005
R19274 gnd.n3177 gnd.n2908 9.3005
R19275 gnd.n3179 gnd.n3178 9.3005
R19276 gnd.n2904 gnd.n2903 9.3005
R19277 gnd.n3192 gnd.n3191 9.3005
R19278 gnd.n3193 gnd.n2902 9.3005
R19279 gnd.n3196 gnd.n3195 9.3005
R19280 gnd.n3046 gnd.n3045 9.3005
R19281 gnd.n3051 gnd.n3050 9.3005
R19282 gnd.n3054 gnd.n3039 9.3005
R19283 gnd.n3055 gnd.n3038 9.3005
R19284 gnd.n3058 gnd.n3037 9.3005
R19285 gnd.n3059 gnd.n3036 9.3005
R19286 gnd.n3062 gnd.n3035 9.3005
R19287 gnd.n3063 gnd.n3034 9.3005
R19288 gnd.n3066 gnd.n3033 9.3005
R19289 gnd.n3067 gnd.n3032 9.3005
R19290 gnd.n3070 gnd.n3031 9.3005
R19291 gnd.n3071 gnd.n3030 9.3005
R19292 gnd.n3074 gnd.n3029 9.3005
R19293 gnd.n3075 gnd.n3028 9.3005
R19294 gnd.n3078 gnd.n3027 9.3005
R19295 gnd.n3079 gnd.n3026 9.3005
R19296 gnd.n3082 gnd.n3025 9.3005
R19297 gnd.n3085 gnd.n3084 9.3005
R19298 gnd.n3049 gnd.n3043 9.3005
R19299 gnd.n3048 gnd.n3047 9.3005
R19300 gnd.n3092 gnd.n3091 9.3005
R19301 gnd.n3090 gnd.n3024 9.3005
R19302 gnd.n3089 gnd.n3088 9.3005
R19303 gnd.n3087 gnd.n1080 9.3005
R19304 gnd.n5043 gnd.n1081 9.3005
R19305 gnd.n5042 gnd.n1082 9.3005
R19306 gnd.n5041 gnd.n1083 9.3005
R19307 gnd.n1099 gnd.n1084 9.3005
R19308 gnd.n5031 gnd.n1100 9.3005
R19309 gnd.n5030 gnd.n1101 9.3005
R19310 gnd.n5029 gnd.n1102 9.3005
R19311 gnd.n1121 gnd.n1103 9.3005
R19312 gnd.n5019 gnd.n1122 9.3005
R19313 gnd.n5018 gnd.n1123 9.3005
R19314 gnd.n5017 gnd.n1124 9.3005
R19315 gnd.n1142 gnd.n1125 9.3005
R19316 gnd.n5007 gnd.n1143 9.3005
R19317 gnd.n5006 gnd.n1144 9.3005
R19318 gnd.n5005 gnd.n1145 9.3005
R19319 gnd.n1163 gnd.n1146 9.3005
R19320 gnd.n4995 gnd.n1164 9.3005
R19321 gnd.n4994 gnd.n1165 9.3005
R19322 gnd.n4993 gnd.n1166 9.3005
R19323 gnd.n1182 gnd.n1167 9.3005
R19324 gnd.n4983 gnd.n1183 9.3005
R19325 gnd.n4982 gnd.n1184 9.3005
R19326 gnd.n4981 gnd.n1185 9.3005
R19327 gnd.n1200 gnd.n1186 9.3005
R19328 gnd.n4970 gnd.n1201 9.3005
R19329 gnd.n4969 gnd.n1202 9.3005
R19330 gnd.n4968 gnd.n1203 9.3005
R19331 gnd.n1220 gnd.n1204 9.3005
R19332 gnd.n4958 gnd.n1221 9.3005
R19333 gnd.n4957 gnd.n1222 9.3005
R19334 gnd.n4956 gnd.n1223 9.3005
R19335 gnd.n1241 gnd.n1224 9.3005
R19336 gnd.n4946 gnd.n1242 9.3005
R19337 gnd.n4945 gnd.n1243 9.3005
R19338 gnd.n4944 gnd.n1244 9.3005
R19339 gnd.n1262 gnd.n1245 9.3005
R19340 gnd.n4934 gnd.n1263 9.3005
R19341 gnd.n4933 gnd.n1264 9.3005
R19342 gnd.n4932 gnd.n1265 9.3005
R19343 gnd.n1283 gnd.n1266 9.3005
R19344 gnd.n4922 gnd.n1284 9.3005
R19345 gnd.n4921 gnd.n1285 9.3005
R19346 gnd.n4920 gnd.n1286 9.3005
R19347 gnd.n1305 gnd.n1287 9.3005
R19348 gnd.n4910 gnd.n1306 9.3005
R19349 gnd.n4909 gnd.n1307 9.3005
R19350 gnd.n4908 gnd.n1308 9.3005
R19351 gnd.n1325 gnd.n1309 9.3005
R19352 gnd.n4898 gnd.n4897 9.3005
R19353 gnd.n3086 gnd.n3023 9.3005
R19354 gnd.n5057 gnd.n5056 9.3005
R19355 gnd.n5055 gnd.n1058 9.3005
R19356 gnd.n5054 gnd.n5053 9.3005
R19357 gnd.n1060 gnd.n1059 9.3005
R19358 gnd.n3125 gnd.n3124 9.3005
R19359 gnd.n3128 gnd.n3127 9.3005
R19360 gnd.n3129 gnd.n3123 9.3005
R19361 gnd.n3132 gnd.n3130 9.3005
R19362 gnd.n3133 gnd.n3122 9.3005
R19363 gnd.n3136 gnd.n3135 9.3005
R19364 gnd.n3137 gnd.n3121 9.3005
R19365 gnd.n3139 gnd.n3138 9.3005
R19366 gnd.n3011 gnd.n3010 9.3005
R19367 gnd.n3152 gnd.n3151 9.3005
R19368 gnd.n3153 gnd.n3009 9.3005
R19369 gnd.n3155 gnd.n3154 9.3005
R19370 gnd.n2914 gnd.n2913 9.3005
R19371 gnd.n3168 gnd.n3167 9.3005
R19372 gnd.n3169 gnd.n2912 9.3005
R19373 gnd.n3171 gnd.n3170 9.3005
R19374 gnd.n2907 gnd.n2906 9.3005
R19375 gnd.n3184 gnd.n3183 9.3005
R19376 gnd.n3185 gnd.n2905 9.3005
R19377 gnd.n3187 gnd.n3186 9.3005
R19378 gnd.n2900 gnd.n2899 9.3005
R19379 gnd.n3201 gnd.n3200 9.3005
R19380 gnd.n3203 gnd.n2897 9.3005
R19381 gnd.n3205 gnd.n3204 9.3005
R19382 gnd.n2892 gnd.n2891 9.3005
R19383 gnd.n3218 gnd.n3217 9.3005
R19384 gnd.n3219 gnd.n2890 9.3005
R19385 gnd.n3221 gnd.n3220 9.3005
R19386 gnd.n2885 gnd.n2884 9.3005
R19387 gnd.n3234 gnd.n3233 9.3005
R19388 gnd.n3235 gnd.n2883 9.3005
R19389 gnd.n3237 gnd.n3236 9.3005
R19390 gnd.n2878 gnd.n2877 9.3005
R19391 gnd.n3250 gnd.n3249 9.3005
R19392 gnd.n3251 gnd.n2876 9.3005
R19393 gnd.n3254 gnd.n3253 9.3005
R19394 gnd.n3252 gnd.n2870 9.3005
R19395 gnd.n3266 gnd.n2871 9.3005
R19396 gnd.n3267 gnd.n2869 9.3005
R19397 gnd.n3269 gnd.n3268 9.3005
R19398 gnd.n3270 gnd.n2868 9.3005
R19399 gnd.n3274 gnd.n3271 9.3005
R19400 gnd.n3275 gnd.n2867 9.3005
R19401 gnd.n3279 gnd.n3278 9.3005
R19402 gnd.n3280 gnd.n2866 9.3005
R19403 gnd.n3283 gnd.n3282 9.3005
R19404 gnd.n3281 gnd.n2640 9.3005
R19405 gnd.n3452 gnd.n2639 9.3005
R19406 gnd.n3454 gnd.n3453 9.3005
R19407 gnd.n5058 gnd.n1056 9.3005
R19408 gnd.n5065 gnd.n5064 9.3005
R19409 gnd.n5066 gnd.n1050 9.3005
R19410 gnd.n5069 gnd.n1049 9.3005
R19411 gnd.n5070 gnd.n1048 9.3005
R19412 gnd.n5073 gnd.n1047 9.3005
R19413 gnd.n5074 gnd.n1046 9.3005
R19414 gnd.n5077 gnd.n1045 9.3005
R19415 gnd.n5078 gnd.n1044 9.3005
R19416 gnd.n5081 gnd.n1043 9.3005
R19417 gnd.n5082 gnd.n1042 9.3005
R19418 gnd.n5085 gnd.n1041 9.3005
R19419 gnd.n5086 gnd.n1040 9.3005
R19420 gnd.n5089 gnd.n1039 9.3005
R19421 gnd.n5090 gnd.n1038 9.3005
R19422 gnd.n5093 gnd.n1037 9.3005
R19423 gnd.n5094 gnd.n1036 9.3005
R19424 gnd.n5097 gnd.n1035 9.3005
R19425 gnd.n5098 gnd.n1034 9.3005
R19426 gnd.n5101 gnd.n1033 9.3005
R19427 gnd.n5103 gnd.n1030 9.3005
R19428 gnd.n5106 gnd.n1029 9.3005
R19429 gnd.n5107 gnd.n1028 9.3005
R19430 gnd.n5110 gnd.n1027 9.3005
R19431 gnd.n5111 gnd.n1026 9.3005
R19432 gnd.n5114 gnd.n1025 9.3005
R19433 gnd.n5115 gnd.n1024 9.3005
R19434 gnd.n5118 gnd.n1023 9.3005
R19435 gnd.n5119 gnd.n1022 9.3005
R19436 gnd.n5122 gnd.n1021 9.3005
R19437 gnd.n5123 gnd.n1020 9.3005
R19438 gnd.n5126 gnd.n1019 9.3005
R19439 gnd.n5127 gnd.n1018 9.3005
R19440 gnd.n5130 gnd.n1017 9.3005
R19441 gnd.n5132 gnd.n1016 9.3005
R19442 gnd.n5133 gnd.n1015 9.3005
R19443 gnd.n5134 gnd.n1014 9.3005
R19444 gnd.n5135 gnd.n1013 9.3005
R19445 gnd.n5063 gnd.n1055 9.3005
R19446 gnd.n5062 gnd.n5061 9.3005
R19447 gnd.n3098 gnd.n3097 9.3005
R19448 gnd.n3096 gnd.n1069 9.3005
R19449 gnd.n5049 gnd.n1070 9.3005
R19450 gnd.n5048 gnd.n1071 9.3005
R19451 gnd.n5047 gnd.n1072 9.3005
R19452 gnd.n1090 gnd.n1073 9.3005
R19453 gnd.n5037 gnd.n1091 9.3005
R19454 gnd.n5036 gnd.n1092 9.3005
R19455 gnd.n5035 gnd.n1093 9.3005
R19456 gnd.n1110 gnd.n1094 9.3005
R19457 gnd.n5025 gnd.n1111 9.3005
R19458 gnd.n5024 gnd.n1112 9.3005
R19459 gnd.n5023 gnd.n1113 9.3005
R19460 gnd.n1132 gnd.n1114 9.3005
R19461 gnd.n5013 gnd.n1133 9.3005
R19462 gnd.n5012 gnd.n1134 9.3005
R19463 gnd.n5011 gnd.n1135 9.3005
R19464 gnd.n1152 gnd.n1136 9.3005
R19465 gnd.n5001 gnd.n1153 9.3005
R19466 gnd.n5000 gnd.n1154 9.3005
R19467 gnd.n4999 gnd.n1155 9.3005
R19468 gnd.n4963 gnd.n1212 9.3005
R19469 gnd.n4962 gnd.n1213 9.3005
R19470 gnd.n1230 gnd.n1214 9.3005
R19471 gnd.n4952 gnd.n1231 9.3005
R19472 gnd.n4951 gnd.n1232 9.3005
R19473 gnd.n4950 gnd.n1233 9.3005
R19474 gnd.n1252 gnd.n1234 9.3005
R19475 gnd.n4940 gnd.n1253 9.3005
R19476 gnd.n4939 gnd.n1254 9.3005
R19477 gnd.n4938 gnd.n1255 9.3005
R19478 gnd.n1272 gnd.n1256 9.3005
R19479 gnd.n4928 gnd.n1273 9.3005
R19480 gnd.n4927 gnd.n1274 9.3005
R19481 gnd.n4926 gnd.n1275 9.3005
R19482 gnd.n1294 gnd.n1276 9.3005
R19483 gnd.n4916 gnd.n1295 9.3005
R19484 gnd.n4915 gnd.n1296 9.3005
R19485 gnd.n4914 gnd.n1297 9.3005
R19486 gnd.n1315 gnd.n1298 9.3005
R19487 gnd.n4904 gnd.n1316 9.3005
R19488 gnd.n4903 gnd.n1317 9.3005
R19489 gnd.n4902 gnd.n1318 9.3005
R19490 gnd.n3095 gnd.n3094 9.3005
R19491 gnd.n4988 gnd.n1175 9.3005
R19492 gnd.n4964 gnd.n1175 9.3005
R19493 gnd.n2928 gnd.n2927 9.3005
R19494 gnd.n2919 gnd.n2918 9.3005
R19495 gnd.n2933 gnd.n2932 9.3005
R19496 gnd.n2934 gnd.n2917 9.3005
R19497 gnd.n3003 gnd.n2935 9.3005
R19498 gnd.n3002 gnd.n2936 9.3005
R19499 gnd.n3001 gnd.n2937 9.3005
R19500 gnd.n2994 gnd.n2938 9.3005
R19501 gnd.n2926 gnd.n2921 9.3005
R19502 gnd.n2922 gnd.n905 9.3005
R19503 gnd.n6531 gnd.n904 9.3005
R19504 gnd.n6532 gnd.n903 9.3005
R19505 gnd.n6533 gnd.n902 9.3005
R19506 gnd.n901 gnd.n897 9.3005
R19507 gnd.n6539 gnd.n896 9.3005
R19508 gnd.n6540 gnd.n895 9.3005
R19509 gnd.n6541 gnd.n894 9.3005
R19510 gnd.n893 gnd.n889 9.3005
R19511 gnd.n6547 gnd.n888 9.3005
R19512 gnd.n6548 gnd.n887 9.3005
R19513 gnd.n6549 gnd.n886 9.3005
R19514 gnd.n885 gnd.n881 9.3005
R19515 gnd.n6555 gnd.n880 9.3005
R19516 gnd.n6556 gnd.n879 9.3005
R19517 gnd.n6557 gnd.n878 9.3005
R19518 gnd.n877 gnd.n873 9.3005
R19519 gnd.n6563 gnd.n872 9.3005
R19520 gnd.n6564 gnd.n871 9.3005
R19521 gnd.n6565 gnd.n870 9.3005
R19522 gnd.n869 gnd.n865 9.3005
R19523 gnd.n6571 gnd.n864 9.3005
R19524 gnd.n6572 gnd.n863 9.3005
R19525 gnd.n6573 gnd.n862 9.3005
R19526 gnd.n861 gnd.n857 9.3005
R19527 gnd.n6579 gnd.n856 9.3005
R19528 gnd.n6580 gnd.n855 9.3005
R19529 gnd.n6581 gnd.n854 9.3005
R19530 gnd.n853 gnd.n849 9.3005
R19531 gnd.n6587 gnd.n848 9.3005
R19532 gnd.n6588 gnd.n847 9.3005
R19533 gnd.n6589 gnd.n846 9.3005
R19534 gnd.n845 gnd.n841 9.3005
R19535 gnd.n6595 gnd.n840 9.3005
R19536 gnd.n6596 gnd.n839 9.3005
R19537 gnd.n6597 gnd.n838 9.3005
R19538 gnd.n837 gnd.n833 9.3005
R19539 gnd.n6603 gnd.n832 9.3005
R19540 gnd.n6604 gnd.n831 9.3005
R19541 gnd.n6605 gnd.n830 9.3005
R19542 gnd.n829 gnd.n825 9.3005
R19543 gnd.n6611 gnd.n824 9.3005
R19544 gnd.n6612 gnd.n823 9.3005
R19545 gnd.n6613 gnd.n822 9.3005
R19546 gnd.n821 gnd.n817 9.3005
R19547 gnd.n6619 gnd.n816 9.3005
R19548 gnd.n6620 gnd.n815 9.3005
R19549 gnd.n6621 gnd.n814 9.3005
R19550 gnd.n813 gnd.n809 9.3005
R19551 gnd.n6627 gnd.n808 9.3005
R19552 gnd.n6628 gnd.n807 9.3005
R19553 gnd.n6629 gnd.n806 9.3005
R19554 gnd.n805 gnd.n801 9.3005
R19555 gnd.n6635 gnd.n800 9.3005
R19556 gnd.n6636 gnd.n799 9.3005
R19557 gnd.n6637 gnd.n798 9.3005
R19558 gnd.n797 gnd.n793 9.3005
R19559 gnd.n6643 gnd.n792 9.3005
R19560 gnd.n6644 gnd.n791 9.3005
R19561 gnd.n6645 gnd.n790 9.3005
R19562 gnd.n789 gnd.n785 9.3005
R19563 gnd.n6651 gnd.n784 9.3005
R19564 gnd.n6652 gnd.n783 9.3005
R19565 gnd.n6653 gnd.n782 9.3005
R19566 gnd.n781 gnd.n777 9.3005
R19567 gnd.n6659 gnd.n776 9.3005
R19568 gnd.n6660 gnd.n775 9.3005
R19569 gnd.n6661 gnd.n774 9.3005
R19570 gnd.n773 gnd.n769 9.3005
R19571 gnd.n6667 gnd.n768 9.3005
R19572 gnd.n6668 gnd.n767 9.3005
R19573 gnd.n6669 gnd.n766 9.3005
R19574 gnd.n765 gnd.n761 9.3005
R19575 gnd.n6675 gnd.n760 9.3005
R19576 gnd.n6676 gnd.n759 9.3005
R19577 gnd.n6677 gnd.n758 9.3005
R19578 gnd.n757 gnd.n753 9.3005
R19579 gnd.n6683 gnd.n752 9.3005
R19580 gnd.n6684 gnd.n751 9.3005
R19581 gnd.n6685 gnd.n750 9.3005
R19582 gnd.n749 gnd.n745 9.3005
R19583 gnd.n6691 gnd.n744 9.3005
R19584 gnd.n6692 gnd.n743 9.3005
R19585 gnd.n6693 gnd.n742 9.3005
R19586 gnd.n2925 gnd.n2924 9.3005
R19587 gnd.n1702 gnd.n1701 9.3005
R19588 gnd.n1680 gnd.n1679 9.3005
R19589 gnd.n1714 gnd.n1713 9.3005
R19590 gnd.n1677 gnd.n1675 9.3005
R19591 gnd.n1721 gnd.n1720 9.3005
R19592 gnd.n1671 gnd.n1670 9.3005
R19593 gnd.n1733 gnd.n1732 9.3005
R19594 gnd.n1668 gnd.n1666 9.3005
R19595 gnd.n1740 gnd.n1739 9.3005
R19596 gnd.n1662 gnd.n1661 9.3005
R19597 gnd.n1752 gnd.n1751 9.3005
R19598 gnd.n1659 gnd.n1657 9.3005
R19599 gnd.n1759 gnd.n1758 9.3005
R19600 gnd.n1653 gnd.n1652 9.3005
R19601 gnd.n1771 gnd.n1770 9.3005
R19602 gnd.n1650 gnd.n1648 9.3005
R19603 gnd.n4475 gnd.n4474 9.3005
R19604 gnd.n4473 gnd.n1649 9.3005
R19605 gnd.n1697 gnd.n1695 9.3005
R19606 gnd.n1768 gnd.n1767 9.3005
R19607 gnd.n1658 gnd.n1654 9.3005
R19608 gnd.n1761 gnd.n1760 9.3005
R19609 gnd.n1750 gnd.n1656 9.3005
R19610 gnd.n1749 gnd.n1748 9.3005
R19611 gnd.n1667 gnd.n1663 9.3005
R19612 gnd.n1742 gnd.n1741 9.3005
R19613 gnd.n1731 gnd.n1665 9.3005
R19614 gnd.n1730 gnd.n1729 9.3005
R19615 gnd.n1676 gnd.n1672 9.3005
R19616 gnd.n1723 gnd.n1722 9.3005
R19617 gnd.n1712 gnd.n1674 9.3005
R19618 gnd.n1711 gnd.n1710 9.3005
R19619 gnd.n1696 gnd.n1681 9.3005
R19620 gnd.n1704 gnd.n1703 9.3005
R19621 gnd.n1694 gnd.n1683 9.3005
R19622 gnd.n1769 gnd.n1647 9.3005
R19623 gnd.n4477 gnd.n4476 9.3005
R19624 gnd.n4472 gnd.n4471 9.3005
R19625 gnd.n4470 gnd.n1779 9.3005
R19626 gnd.n4469 gnd.n4468 9.3005
R19627 gnd.n4467 gnd.n1780 9.3005
R19628 gnd.n4466 gnd.n4465 9.3005
R19629 gnd.n4464 gnd.n1787 9.3005
R19630 gnd.n4463 gnd.n4462 9.3005
R19631 gnd.n4461 gnd.n1788 9.3005
R19632 gnd.n4460 gnd.n4459 9.3005
R19633 gnd.n4458 gnd.n1799 9.3005
R19634 gnd.n3425 gnd.n2664 9.3005
R19635 gnd.n3424 gnd.n3423 9.3005
R19636 gnd.n3422 gnd.n2668 9.3005
R19637 gnd.n3421 gnd.n3420 9.3005
R19638 gnd.n3419 gnd.n2669 9.3005
R19639 gnd.n3418 gnd.n3417 9.3005
R19640 gnd.n3416 gnd.n2673 9.3005
R19641 gnd.n3415 gnd.n3414 9.3005
R19642 gnd.n3413 gnd.n2674 9.3005
R19643 gnd.n3412 gnd.n3411 9.3005
R19644 gnd.n3410 gnd.n2678 9.3005
R19645 gnd.n3409 gnd.n3408 9.3005
R19646 gnd.n3407 gnd.n2679 9.3005
R19647 gnd.n3406 gnd.n3405 9.3005
R19648 gnd.n3404 gnd.n2683 9.3005
R19649 gnd.n3403 gnd.n3402 9.3005
R19650 gnd.n2378 gnd.n2377 9.3005
R19651 gnd.n3576 gnd.n3575 9.3005
R19652 gnd.n3577 gnd.n2375 9.3005
R19653 gnd.n3580 gnd.n3579 9.3005
R19654 gnd.n3578 gnd.n2376 9.3005
R19655 gnd.n2349 gnd.n2348 9.3005
R19656 gnd.n3615 gnd.n3614 9.3005
R19657 gnd.n3616 gnd.n2346 9.3005
R19658 gnd.n3655 gnd.n3654 9.3005
R19659 gnd.n3653 gnd.n2347 9.3005
R19660 gnd.n3652 gnd.n3651 9.3005
R19661 gnd.n3650 gnd.n3617 9.3005
R19662 gnd.n3649 gnd.n3648 9.3005
R19663 gnd.n3647 gnd.n3621 9.3005
R19664 gnd.n3646 gnd.n3645 9.3005
R19665 gnd.n3644 gnd.n3622 9.3005
R19666 gnd.n3643 gnd.n3642 9.3005
R19667 gnd.n3641 gnd.n3627 9.3005
R19668 gnd.n3640 gnd.n3639 9.3005
R19669 gnd.n3638 gnd.n3628 9.3005
R19670 gnd.n3637 gnd.n3636 9.3005
R19671 gnd.n3635 gnd.n3634 9.3005
R19672 gnd.n2264 gnd.n2263 9.3005
R19673 gnd.n3793 gnd.n3792 9.3005
R19674 gnd.n3794 gnd.n2261 9.3005
R19675 gnd.n3831 gnd.n3830 9.3005
R19676 gnd.n3829 gnd.n2262 9.3005
R19677 gnd.n3828 gnd.n3827 9.3005
R19678 gnd.n3826 gnd.n3795 9.3005
R19679 gnd.n3825 gnd.n3824 9.3005
R19680 gnd.n3823 gnd.n3799 9.3005
R19681 gnd.n3822 gnd.n3821 9.3005
R19682 gnd.n3820 gnd.n3800 9.3005
R19683 gnd.n3819 gnd.n3818 9.3005
R19684 gnd.n3817 gnd.n3803 9.3005
R19685 gnd.n3816 gnd.n3815 9.3005
R19686 gnd.n3814 gnd.n3804 9.3005
R19687 gnd.n3813 gnd.n3812 9.3005
R19688 gnd.n3811 gnd.n3810 9.3005
R19689 gnd.n2177 gnd.n2176 9.3005
R19690 gnd.n3970 gnd.n3969 9.3005
R19691 gnd.n3971 gnd.n2174 9.3005
R19692 gnd.n3993 gnd.n3992 9.3005
R19693 gnd.n3991 gnd.n2175 9.3005
R19694 gnd.n3990 gnd.n3989 9.3005
R19695 gnd.n3988 gnd.n3972 9.3005
R19696 gnd.n3987 gnd.n3986 9.3005
R19697 gnd.n3985 gnd.n3976 9.3005
R19698 gnd.n3984 gnd.n3983 9.3005
R19699 gnd.n3982 gnd.n3977 9.3005
R19700 gnd.n3981 gnd.n3980 9.3005
R19701 gnd.n2112 gnd.n2111 9.3005
R19702 gnd.n4102 gnd.n4101 9.3005
R19703 gnd.n4103 gnd.n2109 9.3005
R19704 gnd.n4106 gnd.n4105 9.3005
R19705 gnd.n4104 gnd.n2110 9.3005
R19706 gnd.n2085 gnd.n2084 9.3005
R19707 gnd.n4141 gnd.n4140 9.3005
R19708 gnd.n4142 gnd.n2082 9.3005
R19709 gnd.n4158 gnd.n4157 9.3005
R19710 gnd.n4156 gnd.n2083 9.3005
R19711 gnd.n4155 gnd.n4154 9.3005
R19712 gnd.n4153 gnd.n4143 9.3005
R19713 gnd.n4152 gnd.n4151 9.3005
R19714 gnd.n4150 gnd.n4147 9.3005
R19715 gnd.n4149 gnd.n4148 9.3005
R19716 gnd.n1850 gnd.n1849 9.3005
R19717 gnd.n4373 gnd.n4372 9.3005
R19718 gnd.n4374 gnd.n1848 9.3005
R19719 gnd.n4376 gnd.n4375 9.3005
R19720 gnd.n1838 gnd.n1837 9.3005
R19721 gnd.n4393 gnd.n4392 9.3005
R19722 gnd.n4394 gnd.n1836 9.3005
R19723 gnd.n4396 gnd.n4395 9.3005
R19724 gnd.n1825 gnd.n1824 9.3005
R19725 gnd.n4413 gnd.n4412 9.3005
R19726 gnd.n4414 gnd.n1823 9.3005
R19727 gnd.n4416 gnd.n4415 9.3005
R19728 gnd.n1812 gnd.n1811 9.3005
R19729 gnd.n4433 gnd.n4432 9.3005
R19730 gnd.n4434 gnd.n1810 9.3005
R19731 gnd.n4437 gnd.n4436 9.3005
R19732 gnd.n4435 gnd.n1801 9.3005
R19733 gnd.n4455 gnd.n1800 9.3005
R19734 gnd.n4457 gnd.n4456 9.3005
R19735 gnd.n3427 gnd.n3426 9.3005
R19736 gnd.n3430 gnd.n3429 9.3005
R19737 gnd.n3431 gnd.n2659 9.3005
R19738 gnd.n3433 gnd.n3432 9.3005
R19739 gnd.n3435 gnd.n3434 9.3005
R19740 gnd.n3436 gnd.n2652 9.3005
R19741 gnd.n3438 gnd.n3437 9.3005
R19742 gnd.n3439 gnd.n2651 9.3005
R19743 gnd.n3441 gnd.n3440 9.3005
R19744 gnd.n3442 gnd.n2645 9.3005
R19745 gnd.n3428 gnd.n2663 9.3005
R19746 gnd.n2895 gnd.n2894 9.3005
R19747 gnd.n3210 gnd.n3209 9.3005
R19748 gnd.n3211 gnd.n2893 9.3005
R19749 gnd.n3213 gnd.n3212 9.3005
R19750 gnd.n2889 gnd.n2888 9.3005
R19751 gnd.n3226 gnd.n3225 9.3005
R19752 gnd.n3227 gnd.n2887 9.3005
R19753 gnd.n3229 gnd.n3228 9.3005
R19754 gnd.n2881 gnd.n2880 9.3005
R19755 gnd.n3242 gnd.n3241 9.3005
R19756 gnd.n3243 gnd.n2879 9.3005
R19757 gnd.n3245 gnd.n3244 9.3005
R19758 gnd.n2875 gnd.n2874 9.3005
R19759 gnd.n3259 gnd.n3258 9.3005
R19760 gnd.n3260 gnd.n2873 9.3005
R19761 gnd.n3262 gnd.n3261 9.3005
R19762 gnd.n2861 gnd.n2859 9.3005
R19763 gnd.n3297 gnd.n3296 9.3005
R19764 gnd.n3295 gnd.n2860 9.3005
R19765 gnd.n3294 gnd.n3293 9.3005
R19766 gnd.n3292 gnd.n2862 9.3005
R19767 gnd.n3291 gnd.n3290 9.3005
R19768 gnd.n3289 gnd.n2865 9.3005
R19769 gnd.n3288 gnd.n3287 9.3005
R19770 gnd.n2644 gnd.n2642 9.3005
R19771 gnd.n3448 gnd.n3447 9.3005
R19772 gnd.n3446 gnd.n2643 9.3005
R19773 gnd.n3444 gnd.n3443 9.3005
R19774 gnd.n2647 gnd.n2646 9.3005
R19775 gnd.n2796 gnd.n2795 9.3005
R19776 gnd.n2798 gnd.n2797 9.3005
R19777 gnd.n2776 gnd.n2775 9.3005
R19778 gnd.n2804 gnd.n2803 9.3005
R19779 gnd.n2806 gnd.n2805 9.3005
R19780 gnd.n2766 gnd.n2765 9.3005
R19781 gnd.n2812 gnd.n2811 9.3005
R19782 gnd.n2814 gnd.n2813 9.3005
R19783 gnd.n2753 gnd.n2752 9.3005
R19784 gnd.n2820 gnd.n2819 9.3005
R19785 gnd.n2822 gnd.n2821 9.3005
R19786 gnd.n2743 gnd.n2742 9.3005
R19787 gnd.n2828 gnd.n2827 9.3005
R19788 gnd.n2830 gnd.n2829 9.3005
R19789 gnd.n2728 gnd.n2726 9.3005
R19790 gnd.n2836 gnd.n2835 9.3005
R19791 gnd.n2837 gnd.n2725 9.3005
R19792 gnd.n2730 gnd.n1327 9.3005
R19793 gnd.n2729 gnd.n2727 9.3005
R19794 gnd.n2834 gnd.n2833 9.3005
R19795 gnd.n2832 gnd.n2831 9.3005
R19796 gnd.n2738 gnd.n2737 9.3005
R19797 gnd.n2826 gnd.n2825 9.3005
R19798 gnd.n2824 gnd.n2823 9.3005
R19799 gnd.n2749 gnd.n2748 9.3005
R19800 gnd.n2818 gnd.n2817 9.3005
R19801 gnd.n2816 gnd.n2815 9.3005
R19802 gnd.n2760 gnd.n2759 9.3005
R19803 gnd.n2810 gnd.n2809 9.3005
R19804 gnd.n2808 gnd.n2807 9.3005
R19805 gnd.n2772 gnd.n2771 9.3005
R19806 gnd.n2802 gnd.n2801 9.3005
R19807 gnd.n2800 gnd.n2799 9.3005
R19808 gnd.n2785 gnd.n2784 9.3005
R19809 gnd.n2794 gnd.n2793 9.3005
R19810 gnd.n4892 gnd.n1328 9.3005
R19811 gnd.n4891 gnd.n4890 9.3005
R19812 gnd.n4889 gnd.n1332 9.3005
R19813 gnd.n4888 gnd.n4887 9.3005
R19814 gnd.n4886 gnd.n1333 9.3005
R19815 gnd.n4885 gnd.n4884 9.3005
R19816 gnd.n4883 gnd.n1337 9.3005
R19817 gnd.n4882 gnd.n4881 9.3005
R19818 gnd.n4880 gnd.n1338 9.3005
R19819 gnd.n4879 gnd.n4878 9.3005
R19820 gnd.n4877 gnd.n1342 9.3005
R19821 gnd.n4876 gnd.n4875 9.3005
R19822 gnd.n4874 gnd.n1343 9.3005
R19823 gnd.n4873 gnd.n4872 9.3005
R19824 gnd.n4871 gnd.n1347 9.3005
R19825 gnd.n4870 gnd.n4869 9.3005
R19826 gnd.n4868 gnd.n1348 9.3005
R19827 gnd.n4867 gnd.n4866 9.3005
R19828 gnd.n4865 gnd.n1352 9.3005
R19829 gnd.n4864 gnd.n4863 9.3005
R19830 gnd.n4862 gnd.n1353 9.3005
R19831 gnd.n4861 gnd.n4860 9.3005
R19832 gnd.n4859 gnd.n1357 9.3005
R19833 gnd.n4858 gnd.n4857 9.3005
R19834 gnd.n4856 gnd.n1358 9.3005
R19835 gnd.n4855 gnd.n4854 9.3005
R19836 gnd.n4853 gnd.n1362 9.3005
R19837 gnd.n4852 gnd.n4851 9.3005
R19838 gnd.n4850 gnd.n1363 9.3005
R19839 gnd.n4849 gnd.n4848 9.3005
R19840 gnd.n4847 gnd.n1367 9.3005
R19841 gnd.n4846 gnd.n4845 9.3005
R19842 gnd.n4844 gnd.n1368 9.3005
R19843 gnd.n4843 gnd.n4842 9.3005
R19844 gnd.n4841 gnd.n1372 9.3005
R19845 gnd.n4840 gnd.n4839 9.3005
R19846 gnd.n4838 gnd.n1373 9.3005
R19847 gnd.n4837 gnd.n4836 9.3005
R19848 gnd.n4835 gnd.n1377 9.3005
R19849 gnd.n4834 gnd.n4833 9.3005
R19850 gnd.n4832 gnd.n1378 9.3005
R19851 gnd.n4831 gnd.n4830 9.3005
R19852 gnd.n4829 gnd.n1382 9.3005
R19853 gnd.n4828 gnd.n4827 9.3005
R19854 gnd.n4826 gnd.n1383 9.3005
R19855 gnd.n4825 gnd.n4824 9.3005
R19856 gnd.n4823 gnd.n1387 9.3005
R19857 gnd.n4822 gnd.n4821 9.3005
R19858 gnd.n4820 gnd.n1388 9.3005
R19859 gnd.n4819 gnd.n4818 9.3005
R19860 gnd.n4817 gnd.n1392 9.3005
R19861 gnd.n4816 gnd.n4815 9.3005
R19862 gnd.n4814 gnd.n1393 9.3005
R19863 gnd.n4813 gnd.n4812 9.3005
R19864 gnd.n4811 gnd.n1397 9.3005
R19865 gnd.n4810 gnd.n4809 9.3005
R19866 gnd.n4808 gnd.n1398 9.3005
R19867 gnd.n4807 gnd.n4806 9.3005
R19868 gnd.n4805 gnd.n1402 9.3005
R19869 gnd.n4804 gnd.n4803 9.3005
R19870 gnd.n4802 gnd.n1403 9.3005
R19871 gnd.n4801 gnd.n4800 9.3005
R19872 gnd.n4799 gnd.n1407 9.3005
R19873 gnd.n4798 gnd.n4797 9.3005
R19874 gnd.n4796 gnd.n1408 9.3005
R19875 gnd.n4795 gnd.n4794 9.3005
R19876 gnd.n4793 gnd.n1412 9.3005
R19877 gnd.n4792 gnd.n4791 9.3005
R19878 gnd.n4790 gnd.n1413 9.3005
R19879 gnd.n4789 gnd.n4788 9.3005
R19880 gnd.n4787 gnd.n1417 9.3005
R19881 gnd.n4786 gnd.n4785 9.3005
R19882 gnd.n4784 gnd.n1418 9.3005
R19883 gnd.n4783 gnd.n4782 9.3005
R19884 gnd.n4781 gnd.n1422 9.3005
R19885 gnd.n4780 gnd.n4779 9.3005
R19886 gnd.n4778 gnd.n1423 9.3005
R19887 gnd.n4777 gnd.n4776 9.3005
R19888 gnd.n4775 gnd.n1427 9.3005
R19889 gnd.n4774 gnd.n4773 9.3005
R19890 gnd.n4772 gnd.n1428 9.3005
R19891 gnd.n4771 gnd.n4770 9.3005
R19892 gnd.n4769 gnd.n1432 9.3005
R19893 gnd.n4768 gnd.n4767 9.3005
R19894 gnd.n4766 gnd.n1433 9.3005
R19895 gnd.n4765 gnd.n4764 9.3005
R19896 gnd.n4763 gnd.n1437 9.3005
R19897 gnd.n4762 gnd.n4761 9.3005
R19898 gnd.n4760 gnd.n1438 9.3005
R19899 gnd.n4759 gnd.n4758 9.3005
R19900 gnd.n4757 gnd.n1442 9.3005
R19901 gnd.n4756 gnd.n4755 9.3005
R19902 gnd.n4754 gnd.n1443 9.3005
R19903 gnd.n4753 gnd.n4752 9.3005
R19904 gnd.n4751 gnd.n1447 9.3005
R19905 gnd.n4750 gnd.n4749 9.3005
R19906 gnd.n4748 gnd.n1448 9.3005
R19907 gnd.n4747 gnd.n4746 9.3005
R19908 gnd.n4745 gnd.n1452 9.3005
R19909 gnd.n4744 gnd.n4743 9.3005
R19910 gnd.n4742 gnd.n1453 9.3005
R19911 gnd.n4894 gnd.n4893 9.3005
R19912 gnd.n1689 gnd.n1685 9.3005
R19913 gnd.n1498 gnd.n1496 9.3005
R19914 gnd.n4716 gnd.n4715 9.3005
R19915 gnd.n4714 gnd.n1497 9.3005
R19916 gnd.n4713 gnd.n4712 9.3005
R19917 gnd.n4711 gnd.n1499 9.3005
R19918 gnd.n4710 gnd.n4709 9.3005
R19919 gnd.n4708 gnd.n1503 9.3005
R19920 gnd.n4707 gnd.n4706 9.3005
R19921 gnd.n4705 gnd.n1504 9.3005
R19922 gnd.n4704 gnd.n4703 9.3005
R19923 gnd.n4702 gnd.n1508 9.3005
R19924 gnd.n4701 gnd.n4700 9.3005
R19925 gnd.n4699 gnd.n1509 9.3005
R19926 gnd.n4698 gnd.n4697 9.3005
R19927 gnd.n4696 gnd.n1513 9.3005
R19928 gnd.n4695 gnd.n4694 9.3005
R19929 gnd.n4693 gnd.n1514 9.3005
R19930 gnd.n4692 gnd.n4691 9.3005
R19931 gnd.n4690 gnd.n4689 9.3005
R19932 gnd.n285 gnd.n283 9.3005
R19933 gnd.n7499 gnd.n7498 9.3005
R19934 gnd.n7497 gnd.n284 9.3005
R19935 gnd.n7496 gnd.n7495 9.3005
R19936 gnd.n7494 gnd.n286 9.3005
R19937 gnd.n7493 gnd.n7492 9.3005
R19938 gnd.n7490 gnd.n290 9.3005
R19939 gnd.n7489 gnd.n7488 9.3005
R19940 gnd.n7487 gnd.n292 9.3005
R19941 gnd.n261 gnd.n260 9.3005
R19942 gnd.n7511 gnd.n7510 9.3005
R19943 gnd.n7512 gnd.n259 9.3005
R19944 gnd.n7514 gnd.n7513 9.3005
R19945 gnd.n245 gnd.n244 9.3005
R19946 gnd.n7527 gnd.n7526 9.3005
R19947 gnd.n7528 gnd.n243 9.3005
R19948 gnd.n7530 gnd.n7529 9.3005
R19949 gnd.n230 gnd.n229 9.3005
R19950 gnd.n7543 gnd.n7542 9.3005
R19951 gnd.n7544 gnd.n228 9.3005
R19952 gnd.n7546 gnd.n7545 9.3005
R19953 gnd.n215 gnd.n214 9.3005
R19954 gnd.n7559 gnd.n7558 9.3005
R19955 gnd.n7560 gnd.n213 9.3005
R19956 gnd.n7562 gnd.n7561 9.3005
R19957 gnd.n200 gnd.n199 9.3005
R19958 gnd.n7575 gnd.n7574 9.3005
R19959 gnd.n7576 gnd.n197 9.3005
R19960 gnd.n7653 gnd.n7652 9.3005
R19961 gnd.n7651 gnd.n198 9.3005
R19962 gnd.n7650 gnd.n7649 9.3005
R19963 gnd.n7648 gnd.n7577 9.3005
R19964 gnd.n7647 gnd.n7646 9.3005
R19965 gnd.n1691 gnd.n1690 9.3005
R19966 gnd.n7643 gnd.n7579 9.3005
R19967 gnd.n7642 gnd.n7641 9.3005
R19968 gnd.n7640 gnd.n7584 9.3005
R19969 gnd.n7639 gnd.n7638 9.3005
R19970 gnd.n7637 gnd.n7585 9.3005
R19971 gnd.n7636 gnd.n7635 9.3005
R19972 gnd.n7634 gnd.n7592 9.3005
R19973 gnd.n7633 gnd.n7632 9.3005
R19974 gnd.n7631 gnd.n7593 9.3005
R19975 gnd.n7630 gnd.n7629 9.3005
R19976 gnd.n7628 gnd.n7600 9.3005
R19977 gnd.n7627 gnd.n7626 9.3005
R19978 gnd.n7625 gnd.n7601 9.3005
R19979 gnd.n7624 gnd.n7623 9.3005
R19980 gnd.n7622 gnd.n7608 9.3005
R19981 gnd.n7621 gnd.n7620 9.3005
R19982 gnd.n7619 gnd.n7609 9.3005
R19983 gnd.n7618 gnd.n7617 9.3005
R19984 gnd.n7645 gnd.n7644 9.3005
R19985 gnd.n4482 gnd.n1641 9.3005
R19986 gnd.n4485 gnd.n4484 9.3005
R19987 gnd.n4483 gnd.n1642 9.3005
R19988 gnd.n1622 gnd.n1621 9.3005
R19989 gnd.n4531 gnd.n4530 9.3005
R19990 gnd.n4532 gnd.n1619 9.3005
R19991 gnd.n4535 gnd.n4534 9.3005
R19992 gnd.n4533 gnd.n1620 9.3005
R19993 gnd.n1595 gnd.n1594 9.3005
R19994 gnd.n4563 gnd.n4562 9.3005
R19995 gnd.n4564 gnd.n1592 9.3005
R19996 gnd.n4567 gnd.n4566 9.3005
R19997 gnd.n4565 gnd.n1593 9.3005
R19998 gnd.n1566 gnd.n1565 9.3005
R19999 gnd.n4602 gnd.n4601 9.3005
R20000 gnd.n4603 gnd.n1563 9.3005
R20001 gnd.n4609 gnd.n4608 9.3005
R20002 gnd.n4607 gnd.n1564 9.3005
R20003 gnd.n4606 gnd.n4605 9.3005
R20004 gnd.n1555 gnd.n1554 9.3005
R20005 gnd.n4628 gnd.n4627 9.3005
R20006 gnd.n4629 gnd.n1552 9.3005
R20007 gnd.n4634 gnd.n4633 9.3005
R20008 gnd.n4632 gnd.n1553 9.3005
R20009 gnd.n4631 gnd.n4630 9.3005
R20010 gnd.n69 gnd.n67 9.3005
R20011 gnd.n7784 gnd.n7783 9.3005
R20012 gnd.n7782 gnd.n68 9.3005
R20013 gnd.n7781 gnd.n7780 9.3005
R20014 gnd.n7779 gnd.n73 9.3005
R20015 gnd.n7778 gnd.n7777 9.3005
R20016 gnd.n7776 gnd.n74 9.3005
R20017 gnd.n7775 gnd.n7774 9.3005
R20018 gnd.n7773 gnd.n78 9.3005
R20019 gnd.n7772 gnd.n7771 9.3005
R20020 gnd.n7770 gnd.n79 9.3005
R20021 gnd.n7769 gnd.n7768 9.3005
R20022 gnd.n7767 gnd.n83 9.3005
R20023 gnd.n7766 gnd.n7765 9.3005
R20024 gnd.n7764 gnd.n84 9.3005
R20025 gnd.n7763 gnd.n7762 9.3005
R20026 gnd.n7761 gnd.n88 9.3005
R20027 gnd.n7760 gnd.n7759 9.3005
R20028 gnd.n7758 gnd.n89 9.3005
R20029 gnd.n7757 gnd.n7756 9.3005
R20030 gnd.n7755 gnd.n93 9.3005
R20031 gnd.n7754 gnd.n7753 9.3005
R20032 gnd.n7752 gnd.n94 9.3005
R20033 gnd.n7751 gnd.n7750 9.3005
R20034 gnd.n7749 gnd.n98 9.3005
R20035 gnd.n7748 gnd.n7747 9.3005
R20036 gnd.n7746 gnd.n99 9.3005
R20037 gnd.n7745 gnd.n102 9.3005
R20038 gnd.n4481 gnd.n4480 9.3005
R20039 gnd.t158 gnd.n5262 9.24152
R20040 gnd.t187 gnd.n945 9.24152
R20041 gnd.n6397 gnd.t206 9.24152
R20042 gnd.t194 gnd.n1063 9.24152
R20043 gnd.n4906 gnd.t202 9.24152
R20044 gnd.t91 gnd.n3690 9.24152
R20045 gnd.n4109 gnd.t68 9.24152
R20046 gnd.n4487 gnd.t221 9.24152
R20047 gnd.n7663 gnd.t210 9.24152
R20048 gnd.t2 gnd.t158 8.92286
R20049 gnd.n3703 gnd.n2309 8.92286
R20050 gnd.n3763 gnd.n3762 8.92286
R20051 gnd.n3880 gnd.n2224 8.92286
R20052 gnd.n3941 gnd.n3940 8.92286
R20053 gnd.n4041 gnd.n2136 8.92286
R20054 gnd.n4112 gnd.n4111 8.92286
R20055 gnd.n4208 gnd.n2042 8.92286
R20056 gnd.n6376 gnd.n6351 8.92171
R20057 gnd.n6344 gnd.n6319 8.92171
R20058 gnd.n6312 gnd.n6287 8.92171
R20059 gnd.n6281 gnd.n6256 8.92171
R20060 gnd.n6249 gnd.n6224 8.92171
R20061 gnd.n6217 gnd.n6192 8.92171
R20062 gnd.n6185 gnd.n6160 8.92171
R20063 gnd.n6154 gnd.n6129 8.92171
R20064 gnd.n4230 gnd.n4212 8.72777
R20065 gnd.t144 gnd.n5357 8.60421
R20066 gnd.n3338 gnd.t241 8.60421
R20067 gnd.n3384 gnd.t323 8.60421
R20068 gnd.t10 gnd.n3878 8.60421
R20069 gnd.n3911 gnd.t120 8.60421
R20070 gnd.n4400 gnd.t128 8.60421
R20071 gnd.n4452 gnd.t198 8.60421
R20072 gnd.n5325 gnd.n5309 8.43467
R20073 gnd.n50 gnd.n34 8.43467
R20074 gnd.n3194 gnd.n0 8.41456
R20075 gnd.n7786 gnd.n7785 8.41456
R20076 gnd.n2470 gnd.t245 8.28555
R20077 gnd.n3682 gnd.n2322 8.28555
R20078 gnd.n3755 gnd.n2282 8.28555
R20079 gnd.n3859 gnd.n2237 8.28555
R20080 gnd.n3933 gnd.n2195 8.28555
R20081 gnd.n4021 gnd.n2150 8.28555
R20082 gnd.n4077 gnd.n2101 8.28555
R20083 gnd.n4185 gnd.n2056 8.28555
R20084 gnd.n6377 gnd.n6349 8.14595
R20085 gnd.n6345 gnd.n6317 8.14595
R20086 gnd.n6313 gnd.n6285 8.14595
R20087 gnd.n6282 gnd.n6254 8.14595
R20088 gnd.n6250 gnd.n6222 8.14595
R20089 gnd.n6218 gnd.n6190 8.14595
R20090 gnd.n6186 gnd.n6158 8.14595
R20091 gnd.n6155 gnd.n6127 8.14595
R20092 gnd.n6382 gnd.n6381 7.97301
R20093 gnd.n5850 gnd.t150 7.9669
R20094 gnd.n3335 gnd.n2840 7.9669
R20095 gnd.t57 gnd.n2337 7.9669
R20096 gnd.n4161 gnd.t61 7.9669
R20097 gnd.n1467 gnd.n1458 7.9669
R20098 gnd.n7619 gnd.n7618 7.75808
R20099 gnd.n4477 gnd.n1647 7.75808
R20100 gnd.n2793 gnd.n2784 7.75808
R20101 gnd.n3047 gnd.n3043 7.75808
R20102 gnd.n3682 gnd.t298 7.64824
R20103 gnd.n3840 gnd.t54 7.64824
R20104 gnd.n3739 gnd.t54 7.64824
R20105 gnd.t87 gnd.n3924 7.64824
R20106 gnd.n3926 gnd.t87 7.64824
R20107 gnd.n4077 gnd.t180 7.64824
R20108 gnd.t156 gnd.n5443 7.32958
R20109 gnd.t241 gnd.n2702 7.32958
R20110 gnd.t323 gnd.n3383 7.32958
R20111 gnd.t128 gnd.n4399 7.32958
R20112 gnd.n4440 gnd.t198 7.32958
R20113 gnd.n2443 gnd.n2442 7.30353
R20114 gnd.n4229 gnd.n4228 7.30353
R20115 gnd.n5752 gnd.n5751 7.01093
R20116 gnd.n5762 gnd.n5472 7.01093
R20117 gnd.n5761 gnd.n5475 7.01093
R20118 gnd.n5770 gnd.n5466 7.01093
R20119 gnd.n5774 gnd.n5773 7.01093
R20120 gnd.n5792 gnd.n5451 7.01093
R20121 gnd.n5791 gnd.n5454 7.01093
R20122 gnd.n5802 gnd.n5443 7.01093
R20123 gnd.n5444 gnd.n5432 7.01093
R20124 gnd.n5815 gnd.n5433 7.01093
R20125 gnd.n5826 gnd.n5425 7.01093
R20126 gnd.n5825 gnd.n5416 7.01093
R20127 gnd.n5418 gnd.n5400 7.01093
R20128 gnd.n5862 gnd.n5401 7.01093
R20129 gnd.n5851 gnd.n5850 7.01093
R20130 gnd.n5887 gnd.n5392 7.01093
R20131 gnd.n5898 gnd.n5897 7.01093
R20132 gnd.n5385 gnd.n5377 7.01093
R20133 gnd.n5927 gnd.n5365 7.01093
R20134 gnd.n5926 gnd.n5368 7.01093
R20135 gnd.n5937 gnd.n5357 7.01093
R20136 gnd.n5358 gnd.n5346 7.01093
R20137 gnd.n5948 gnd.n5347 7.01093
R20138 gnd.n5972 gnd.n5290 7.01093
R20139 gnd.n5971 gnd.n5281 7.01093
R20140 gnd.n5283 gnd.n5274 7.01093
R20141 gnd.n5994 gnd.n5993 7.01093
R20142 gnd.n6011 gnd.n5262 7.01093
R20143 gnd.n6010 gnd.n5265 7.01093
R20144 gnd.n6024 gnd.n5254 7.01093
R20145 gnd.n5255 gnd.n5243 7.01093
R20146 gnd.n6034 gnd.n5245 7.01093
R20147 gnd.n6065 gnd.n6064 7.01093
R20148 gnd.n6078 gnd.n6077 7.01093
R20149 gnd.n5224 gnd.n5214 7.01093
R20150 gnd.n6090 gnd.n6089 7.01093
R20151 gnd.n6102 gnd.n909 7.01093
R20152 gnd.n6519 gnd.n920 7.01093
R20153 gnd.n6120 gnd.n6119 7.01093
R20154 gnd.n6513 gnd.n6512 7.01093
R20155 gnd.n5198 gnd.n931 7.01093
R20156 gnd.n6506 gnd.n942 7.01093
R20157 gnd.n6505 gnd.n945 7.01093
R20158 gnd.n6398 gnd.n6397 7.01093
R20159 gnd.n6499 gnd.n6498 7.01093
R20160 gnd.n966 gnd.n956 7.01093
R20161 gnd.n3585 gnd.n2370 7.01093
R20162 gnd.n3763 gnd.n2286 7.01093
R20163 gnd.n2244 gnd.t45 7.01093
R20164 gnd.n3880 gnd.n3879 7.01093
R20165 gnd.n3941 gnd.n2199 7.01093
R20166 gnd.t301 gnd.n2184 7.01093
R20167 gnd.n4041 gnd.n4040 7.01093
R20168 gnd.n4208 gnd.n4207 7.01093
R20169 gnd.n5433 gnd.t154 6.69227
R20170 gnd.n5993 gnd.t2 6.69227
R20171 gnd.n6520 gnd.t149 6.69227
R20172 gnd.n5033 gnd.t106 6.69227
R20173 gnd.n3691 gnd.t91 6.69227
R20174 gnd.n4119 gnd.t68 6.69227
R20175 gnd.t6 gnd.n208 6.69227
R20176 gnd.n4362 gnd.n4361 6.5566
R20177 gnd.n2538 gnd.n2537 6.5566
R20178 gnd.n3504 gnd.n2449 6.5566
R20179 gnd.n4240 gnd.n4239 6.5566
R20180 gnd.n3610 gnd.n2352 6.37362
R20181 gnd.n2455 gnd.n2454 6.37362
R20182 gnd.n3789 gnd.n2268 6.37362
R20183 gnd.n3917 gnd.n3916 6.37362
R20184 gnd.n4137 gnd.n2089 6.37362
R20185 gnd.n4061 gnd.n2075 6.37362
R20186 gnd.t191 gnd.n2037 6.37362
R20187 gnd.n3432 gnd.n2658 6.20656
R20188 gnd.n7708 gnd.n7705 6.20656
R20189 gnd.n5102 gnd.n5101 6.20656
R20190 gnd.n4462 gnd.n1791 6.20656
R20191 gnd.n5886 gnd.t316 6.05496
R20192 gnd.n5885 gnd.t153 6.05496
R20193 gnd.t163 gnd.n5358 6.05496
R20194 gnd.t152 gnd.n5237 6.05496
R20195 gnd.n5027 gnd.n1108 6.05496
R20196 gnd.n5009 gnd.t303 6.05496
R20197 gnd.n3564 gnd.n3563 6.05496
R20198 gnd.n7417 gnd.t27 6.05496
R20199 gnd.n7396 gnd.n218 6.05496
R20200 gnd.n6379 gnd.n6349 5.81868
R20201 gnd.n6347 gnd.n6317 5.81868
R20202 gnd.n6315 gnd.n6285 5.81868
R20203 gnd.n6284 gnd.n6254 5.81868
R20204 gnd.n6252 gnd.n6222 5.81868
R20205 gnd.n6220 gnd.n6190 5.81868
R20206 gnd.n6188 gnd.n6158 5.81868
R20207 gnd.n6157 gnd.n6127 5.81868
R20208 gnd.n2420 gnd.t218 5.73631
R20209 gnd.t218 gnd.n2380 5.73631
R20210 gnd.t225 gnd.n2343 5.73631
R20211 gnd.n3703 gnd.t299 5.73631
R20212 gnd.n3625 gnd.n3624 5.73631
R20213 gnd.n3711 gnd.n2298 5.73631
R20214 gnd.n3748 gnd.t181 5.73631
R20215 gnd.n3879 gnd.t18 5.73631
R20216 gnd.n2220 gnd.n2209 5.73631
R20217 gnd.n3888 gnd.n2212 5.73631
R20218 gnd.t117 gnd.n2199 5.73631
R20219 gnd.n4003 gnd.t135 5.73631
R20220 gnd.n2132 gnd.n2123 5.73631
R20221 gnd.n4049 gnd.n4047 5.73631
R20222 gnd.n4112 gnd.t296 5.73631
R20223 gnd.t252 gnd.n2061 5.73631
R20224 gnd.n4366 gnd.n2031 5.62001
R20225 gnd.n3499 gnd.n2542 5.62001
R20226 gnd.n3500 gnd.n3499 5.62001
R20227 gnd.n4235 gnd.n2031 5.62001
R20228 gnd.n5570 gnd.n5569 5.4308
R20229 gnd.n6412 gnd.n5189 5.4308
R20230 gnd.n5347 gnd.t151 5.41765
R20231 gnd.t143 gnd.n5982 5.41765
R20232 gnd.n6066 gnd.t167 5.41765
R20233 gnd.n4985 gnd.t50 5.41765
R20234 gnd.t59 gnd.n3710 5.41765
R20235 gnd.t33 gnd.n2130 5.41765
R20236 gnd.n7480 gnd.t130 5.41765
R20237 gnd.t258 gnd.n3584 5.09899
R20238 gnd.n3658 gnd.n2343 5.09899
R20239 gnd.n3666 gnd.n2337 5.09899
R20240 gnd.t16 gnd.n2272 5.09899
R20241 gnd.n3834 gnd.n2258 5.09899
R20242 gnd.n3843 gnd.n2252 5.09899
R20243 gnd.n3997 gnd.n2171 5.09899
R20244 gnd.n4005 gnd.n2165 5.09899
R20245 gnd.n2157 gnd.t295 5.09899
R20246 gnd.n4161 gnd.n2079 5.09899
R20247 gnd.n4169 gnd.n2072 5.09899
R20248 gnd.n6377 gnd.n6376 5.04292
R20249 gnd.n6345 gnd.n6344 5.04292
R20250 gnd.n6313 gnd.n6312 5.04292
R20251 gnd.n6282 gnd.n6281 5.04292
R20252 gnd.n6250 gnd.n6249 5.04292
R20253 gnd.n6218 gnd.n6217 5.04292
R20254 gnd.n6186 gnd.n6185 5.04292
R20255 gnd.n6155 gnd.n6154 5.04292
R20256 gnd.n5341 gnd.n5340 4.82753
R20257 gnd.n66 gnd.n65 4.82753
R20258 gnd.t146 gnd.n5908 4.78034
R20259 gnd.n6024 gnd.t147 4.78034
R20260 gnd.n4960 gnd.t133 4.78034
R20261 gnd.t55 gnd.n2387 4.78034
R20262 gnd.n3711 gnd.t59 4.78034
R20263 gnd.n2132 gnd.t33 4.78034
R20264 gnd.n4369 gnd.t264 4.78034
R20265 gnd.n1870 gnd.t161 4.78034
R20266 gnd.n4687 gnd.t109 4.78034
R20267 gnd.n5882 gnd.n5881 4.74817
R20268 gnd.n5877 gnd.n5876 4.74817
R20269 gnd.n5873 gnd.n5872 4.74817
R20270 gnd.n5869 gnd.n5344 4.74817
R20271 gnd.n5881 gnd.n5880 4.74817
R20272 gnd.n5879 gnd.n5877 4.74817
R20273 gnd.n5875 gnd.n5873 4.74817
R20274 gnd.n5871 gnd.n5869 4.74817
R20275 gnd.n7504 gnd.n7503 4.74817
R20276 gnd.n1547 gnd.n271 4.74817
R20277 gnd.n7482 gnd.n270 4.74817
R20278 gnd.n269 gnd.n266 4.74817
R20279 gnd.n7504 gnd.n273 4.74817
R20280 gnd.n4662 gnd.n271 4.74817
R20281 gnd.n1546 gnd.n270 4.74817
R20282 gnd.n7483 gnd.n269 4.74817
R20283 gnd.n2997 gnd.n2996 4.74817
R20284 gnd.n2993 gnd.n2945 4.74817
R20285 gnd.n2986 gnd.n2944 4.74817
R20286 gnd.n2982 gnd.n2943 4.74817
R20287 gnd.n2978 gnd.n2942 4.74817
R20288 gnd.n4669 gnd.n4668 4.74817
R20289 gnd.n4651 gnd.n1539 4.74817
R20290 gnd.n4656 gnd.n4655 4.74817
R20291 gnd.n4652 gnd.n308 4.74817
R20292 gnd.n7470 gnd.n7469 4.74817
R20293 gnd.n4670 gnd.n4669 4.74817
R20294 gnd.n4667 gnd.n1539 4.74817
R20295 gnd.n4657 gnd.n4656 4.74817
R20296 gnd.n4654 gnd.n4652 4.74817
R20297 gnd.n7471 gnd.n7470 4.74817
R20298 gnd.n1174 gnd.n1156 4.74817
R20299 gnd.n1192 gnd.n1176 4.74817
R20300 gnd.n4976 gnd.n4975 4.74817
R20301 gnd.n1211 gnd.n1193 4.74817
R20302 gnd.n4989 gnd.n1174 4.74817
R20303 gnd.n4987 gnd.n1176 4.74817
R20304 gnd.n4977 gnd.n4976 4.74817
R20305 gnd.n4974 gnd.n1193 4.74817
R20306 gnd.n2996 gnd.n2940 4.74817
R20307 gnd.n2993 gnd.n2992 4.74817
R20308 gnd.n2988 gnd.n2944 4.74817
R20309 gnd.n2985 gnd.n2943 4.74817
R20310 gnd.n2981 gnd.n2942 4.74817
R20311 gnd.n5325 gnd.n5324 4.7074
R20312 gnd.n50 gnd.n49 4.7074
R20313 gnd.n5341 gnd.n5325 4.65959
R20314 gnd.n66 gnd.n50 4.65959
R20315 gnd.n2030 gnd.n1947 4.6132
R20316 gnd.n3495 gnd.n3494 4.6132
R20317 gnd.n3573 gnd.n2380 4.46168
R20318 gnd.n2470 gnd.t214 4.46168
R20319 gnd.n3718 gnd.n2303 4.46168
R20320 gnd.n3709 gnd.n2291 4.46168
R20321 gnd.n3895 gnd.n2217 4.46168
R20322 gnd.n3886 gnd.n2203 4.46168
R20323 gnd.n4056 gnd.n2129 4.46168
R20324 gnd.n4099 gnd.n2114 4.46168
R20325 gnd.n4185 gnd.t248 4.46168
R20326 gnd.n4301 gnd.n2037 4.46168
R20327 gnd.n4225 gnd.n4212 4.46111
R20328 gnd.n6362 gnd.n6358 4.38594
R20329 gnd.n6330 gnd.n6326 4.38594
R20330 gnd.n6298 gnd.n6294 4.38594
R20331 gnd.n6267 gnd.n6263 4.38594
R20332 gnd.n6235 gnd.n6231 4.38594
R20333 gnd.n6203 gnd.n6199 4.38594
R20334 gnd.n6171 gnd.n6167 4.38594
R20335 gnd.n6140 gnd.n6136 4.38594
R20336 gnd.n6373 gnd.n6351 4.26717
R20337 gnd.n6341 gnd.n6319 4.26717
R20338 gnd.n6309 gnd.n6287 4.26717
R20339 gnd.n6278 gnd.n6256 4.26717
R20340 gnd.n6246 gnd.n6224 4.26717
R20341 gnd.n6214 gnd.n6192 4.26717
R20342 gnd.n6182 gnd.n6160 4.26717
R20343 gnd.n6151 gnd.n6129 4.26717
R20344 gnd.t148 gnd.n5839 4.14303
R20345 gnd.n6089 gnd.t145 4.14303
R20346 gnd.n3141 gnd.t46 4.14303
R20347 gnd.n4936 gnd.t48 4.14303
R20348 gnd.n3300 gnd.t39 4.14303
R20349 gnd.n3740 gnd.t321 4.14303
R20350 gnd.n3966 gnd.t93 4.14303
R20351 gnd.n1610 gnd.t88 4.14303
R20352 gnd.t31 gnd.n4570 4.14303
R20353 gnd.n7548 gnd.t78 4.14303
R20354 gnd.n6381 gnd.n6380 4.08274
R20355 gnd.n4361 gnd.n4360 4.05904
R20356 gnd.n2537 gnd.n2536 4.05904
R20357 gnd.n3507 gnd.n2449 4.05904
R20358 gnd.n4241 gnd.n4240 4.05904
R20359 gnd.n19 gnd.n9 3.99943
R20360 gnd.n3325 gnd.n2606 3.82437
R20361 gnd.n3585 gnd.t258 3.82437
R20362 gnd.n3602 gnd.n2358 3.82437
R20363 gnd.n3675 gnd.n3674 3.82437
R20364 gnd.t44 gnd.n2286 3.82437
R20365 gnd.n3780 gnd.n2266 3.82437
R20366 gnd.n3852 gnd.n3851 3.82437
R20367 gnd.n3958 gnd.n2179 3.82437
R20368 gnd.n4014 gnd.n4013 3.82437
R20369 gnd.n4040 gnd.t19 3.82437
R20370 gnd.n4129 gnd.n2087 3.82437
R20371 gnd.n4061 gnd.t252 3.82437
R20372 gnd.n4178 gnd.n4177 3.82437
R20373 gnd.n4731 gnd.n1468 3.82437
R20374 gnd.n6381 gnd.n6253 3.70378
R20375 gnd.n5343 gnd.n5342 3.65935
R20376 gnd.n19 gnd.n18 3.60163
R20377 gnd.n6527 gnd.n907 3.50571
R20378 gnd.n6527 gnd.n6526 3.50571
R20379 gnd.n2882 gnd.t20 3.50571
R20380 gnd.t159 gnd.n3364 3.50571
R20381 gnd.t12 gnd.n4418 3.50571
R20382 gnd.n4611 gnd.t4 3.50571
R20383 gnd.n6372 gnd.n6353 3.49141
R20384 gnd.n6340 gnd.n6321 3.49141
R20385 gnd.n6308 gnd.n6289 3.49141
R20386 gnd.n6277 gnd.n6258 3.49141
R20387 gnd.n6245 gnd.n6226 3.49141
R20388 gnd.n6213 gnd.n6194 3.49141
R20389 gnd.n6181 gnd.n6162 3.49141
R20390 gnd.n6150 gnd.n6131 3.49141
R20391 gnd.n3583 gnd.n3582 3.18706
R20392 gnd.t214 gnd.n2356 3.18706
R20393 gnd.n3690 gnd.n3689 3.18706
R20394 gnd.n3761 gnd.n2280 3.18706
R20395 gnd.n3868 gnd.n3866 3.18706
R20396 gnd.n3939 gnd.n2192 3.18706
R20397 gnd.n4029 gnd.n4028 3.18706
R20398 gnd.n4110 gnd.n4109 3.18706
R20399 gnd.n2063 gnd.t248 3.18706
R20400 gnd.n4194 gnd.n4193 3.18706
R20401 gnd.n5840 gnd.t148 2.8684
R20402 gnd.n2896 gnd.t52 2.8684
R20403 gnd.n3657 gnd.t57 2.8684
R20404 gnd.t61 gnd.n4160 2.8684
R20405 gnd.t70 gnd.n1544 2.8684
R20406 gnd.n5326 gnd.t142 2.82907
R20407 gnd.n5326 gnd.t122 2.82907
R20408 gnd.n5328 gnd.t112 2.82907
R20409 gnd.n5328 gnd.t179 2.82907
R20410 gnd.n5330 gnd.t124 2.82907
R20411 gnd.n5330 gnd.t134 2.82907
R20412 gnd.n5332 gnd.t178 2.82907
R20413 gnd.n5332 gnd.t177 2.82907
R20414 gnd.n5334 gnd.t77 2.82907
R20415 gnd.n5334 gnd.t176 2.82907
R20416 gnd.n5336 gnd.t81 2.82907
R20417 gnd.n5336 gnd.t304 2.82907
R20418 gnd.n5338 gnd.t175 2.82907
R20419 gnd.n5338 gnd.t185 2.82907
R20420 gnd.n5295 gnd.t49 2.82907
R20421 gnd.n5295 gnd.t100 2.82907
R20422 gnd.n5297 gnd.t21 2.82907
R20423 gnd.n5297 gnd.t30 2.82907
R20424 gnd.n5299 gnd.t174 2.82907
R20425 gnd.n5299 gnd.t311 2.82907
R20426 gnd.n5301 gnd.t101 2.82907
R20427 gnd.n5301 gnd.t66 2.82907
R20428 gnd.n5303 gnd.t125 2.82907
R20429 gnd.n5303 gnd.t38 2.82907
R20430 gnd.n5305 gnd.t138 2.82907
R20431 gnd.n5305 gnd.t318 2.82907
R20432 gnd.n5307 gnd.t107 2.82907
R20433 gnd.n5307 gnd.t313 2.82907
R20434 gnd.n5310 gnd.t172 2.82907
R20435 gnd.n5310 gnd.t40 2.82907
R20436 gnd.n5312 gnd.t308 2.82907
R20437 gnd.n5312 gnd.t104 2.82907
R20438 gnd.n5314 gnd.t170 2.82907
R20439 gnd.n5314 gnd.t173 2.82907
R20440 gnd.n5316 gnd.t51 2.82907
R20441 gnd.n5316 gnd.t53 2.82907
R20442 gnd.n5318 gnd.t108 2.82907
R20443 gnd.n5318 gnd.t43 2.82907
R20444 gnd.n5320 gnd.t99 2.82907
R20445 gnd.n5320 gnd.t312 2.82907
R20446 gnd.n5322 gnd.t183 2.82907
R20447 gnd.n5322 gnd.t47 2.82907
R20448 gnd.n63 gnd.t79 2.82907
R20449 gnd.n63 gnd.t116 2.82907
R20450 gnd.n61 gnd.t127 2.82907
R20451 gnd.n61 gnd.t83 2.82907
R20452 gnd.n59 gnd.t26 2.82907
R20453 gnd.n59 gnd.t113 2.82907
R20454 gnd.n57 gnd.t114 2.82907
R20455 gnd.n57 gnd.t320 2.82907
R20456 gnd.n55 gnd.t110 2.82907
R20457 gnd.n55 gnd.t126 2.82907
R20458 gnd.n53 gnd.t67 2.82907
R20459 gnd.n53 gnd.t84 2.82907
R20460 gnd.n51 gnd.t115 2.82907
R20461 gnd.n51 gnd.t32 2.82907
R20462 gnd.n32 gnd.t139 2.82907
R20463 gnd.n32 gnd.t169 2.82907
R20464 gnd.n30 gnd.t182 2.82907
R20465 gnd.n30 gnd.t141 2.82907
R20466 gnd.n28 gnd.t137 2.82907
R20467 gnd.n28 gnd.t36 2.82907
R20468 gnd.n26 gnd.t75 2.82907
R20469 gnd.n26 gnd.t132 2.82907
R20470 gnd.n24 gnd.t302 2.82907
R20471 gnd.n24 gnd.t74 2.82907
R20472 gnd.n22 gnd.t72 2.82907
R20473 gnd.n22 gnd.t315 2.82907
R20474 gnd.n20 gnd.t90 2.82907
R20475 gnd.n20 gnd.t103 2.82907
R20476 gnd.n47 gnd.t136 2.82907
R20477 gnd.n47 gnd.t7 2.82907
R20478 gnd.n45 gnd.t28 2.82907
R20479 gnd.n45 gnd.t305 2.82907
R20480 gnd.n43 gnd.t309 2.82907
R20481 gnd.n43 gnd.t171 2.82907
R20482 gnd.n41 gnd.t71 2.82907
R20483 gnd.n41 gnd.t131 2.82907
R20484 gnd.n39 gnd.t314 2.82907
R20485 gnd.n39 gnd.t184 2.82907
R20486 gnd.n37 gnd.t64 2.82907
R20487 gnd.n37 gnd.t5 2.82907
R20488 gnd.n35 gnd.t89 2.82907
R20489 gnd.n35 gnd.t310 2.82907
R20490 gnd.n6369 gnd.n6368 2.71565
R20491 gnd.n6337 gnd.n6336 2.71565
R20492 gnd.n6305 gnd.n6304 2.71565
R20493 gnd.n6274 gnd.n6273 2.71565
R20494 gnd.n6242 gnd.n6241 2.71565
R20495 gnd.n6210 gnd.n6209 2.71565
R20496 gnd.n6178 gnd.n6177 2.71565
R20497 gnd.n6147 gnd.n6146 2.71565
R20498 gnd.n5021 gnd.n1116 2.54975
R20499 gnd.n3149 gnd.n1119 2.54975
R20500 gnd.n5015 gnd.n1127 2.54975
R20501 gnd.n3157 gnd.n1130 2.54975
R20502 gnd.n5009 gnd.n1138 2.54975
R20503 gnd.n3165 gnd.n3005 2.54975
R20504 gnd.n5003 gnd.n1148 2.54975
R20505 gnd.n3173 gnd.n2911 2.54975
R20506 gnd.n4997 gnd.n1158 2.54975
R20507 gnd.n3181 gnd.n1161 2.54975
R20508 gnd.n4991 gnd.n1169 2.54975
R20509 gnd.n3189 gnd.n1172 2.54975
R20510 gnd.n4985 gnd.n1178 2.54975
R20511 gnd.n3198 gnd.n2901 2.54975
R20512 gnd.n4979 gnd.n1188 2.54975
R20513 gnd.n3207 gnd.n2896 2.54975
R20514 gnd.n4972 gnd.n1195 2.54975
R20515 gnd.n3215 gnd.n1198 2.54975
R20516 gnd.n4966 gnd.n1206 2.54975
R20517 gnd.n3223 gnd.n1209 2.54975
R20518 gnd.n4960 gnd.n1216 2.54975
R20519 gnd.n3231 gnd.n2886 2.54975
R20520 gnd.n4954 gnd.n1226 2.54975
R20521 gnd.n3239 gnd.n2882 2.54975
R20522 gnd.n4948 gnd.n1236 2.54975
R20523 gnd.n3247 gnd.n1239 2.54975
R20524 gnd.n4942 gnd.n1247 2.54975
R20525 gnd.n3256 gnd.n1250 2.54975
R20526 gnd.n4936 gnd.n1258 2.54975
R20527 gnd.n3264 gnd.n2872 2.54975
R20528 gnd.n4930 gnd.n1268 2.54975
R20529 gnd.n3300 gnd.n3299 2.54975
R20530 gnd.n4924 gnd.n1278 2.54975
R20531 gnd.n3272 gnd.n1281 2.54975
R20532 gnd.n4918 gnd.n1289 2.54975
R20533 gnd.n3276 gnd.n1292 2.54975
R20534 gnd.n4912 gnd.n1300 2.54975
R20535 gnd.n3285 gnd.n1303 2.54975
R20536 gnd.n4906 gnd.n1311 2.54975
R20537 gnd.n3450 gnd.n2641 2.54975
R20538 gnd.n4900 gnd.n1320 2.54975
R20539 gnd.n3592 gnd.n3591 2.54975
R20540 gnd.n3691 gnd.n2317 2.54975
R20541 gnd.n3725 gnd.t17 2.54975
R20542 gnd.n3770 gnd.n3769 2.54975
R20543 gnd.n3755 gnd.t16 2.54975
R20544 gnd.n3869 gnd.n2232 2.54975
R20545 gnd.n3948 gnd.n3947 2.54975
R20546 gnd.n4021 gnd.t295 2.54975
R20547 gnd.n4030 gnd.n2144 2.54975
R20548 gnd.n4090 gnd.t297 2.54975
R20549 gnd.n4119 gnd.n4118 2.54975
R20550 gnd.n4195 gnd.n2051 2.54975
R20551 gnd.n4725 gnd.n1477 2.54975
R20552 gnd.n4724 gnd.n1480 2.54975
R20553 gnd.n4487 gnd.n1490 2.54975
R20554 gnd.n4718 gnd.n1493 2.54975
R20555 gnd.n1635 gnd.n1634 2.54975
R20556 gnd.n4528 gnd.n4520 2.54975
R20557 gnd.n4538 gnd.n1616 2.54975
R20558 gnd.n4537 gnd.n1605 2.54975
R20559 gnd.n4550 gnd.n4548 2.54975
R20560 gnd.n1610 gnd.n1608 2.54975
R20561 gnd.n4560 gnd.n1598 2.54975
R20562 gnd.n4571 gnd.n1589 2.54975
R20563 gnd.n4570 gnd.n1578 2.54975
R20564 gnd.n4589 gnd.n4588 2.54975
R20565 gnd.n1583 gnd.n1581 2.54975
R20566 gnd.n4599 gnd.n1569 2.54975
R20567 gnd.n1572 gnd.n1561 2.54975
R20568 gnd.n4612 gnd.n4611 2.54975
R20569 gnd.n4679 gnd.n4678 2.54975
R20570 gnd.n1530 gnd.n1528 2.54975
R20571 gnd.n4687 gnd.n1520 2.54975
R20572 gnd.n4625 gnd.n277 2.54975
R20573 gnd.n7501 gnd.n280 2.54975
R20574 gnd.n4637 gnd.n4636 2.54975
R20575 gnd.n4665 gnd.n1541 2.54975
R20576 gnd.n4664 gnd.n1544 2.54975
R20577 gnd.n4660 gnd.n4659 2.54975
R20578 gnd.n4649 gnd.n4648 2.54975
R20579 gnd.n7480 gnd.n294 2.54975
R20580 gnd.n7485 gnd.n296 2.54975
R20581 gnd.n7474 gnd.n7473 2.54975
R20582 gnd.n7508 gnd.n264 2.54975
R20583 gnd.n7406 gnd.n255 2.54975
R20584 gnd.n7516 gnd.n257 2.54975
R20585 gnd.n7413 gnd.n247 2.54975
R20586 gnd.n7524 gnd.n249 2.54975
R20587 gnd.n7417 gnd.n239 2.54975
R20588 gnd.n7532 gnd.n241 2.54975
R20589 gnd.n7458 gnd.n7457 2.54975
R20590 gnd.n7540 gnd.n233 2.54975
R20591 gnd.n7450 gnd.n225 2.54975
R20592 gnd.n5881 gnd.n5343 2.27742
R20593 gnd.n5877 gnd.n5343 2.27742
R20594 gnd.n5873 gnd.n5343 2.27742
R20595 gnd.n5869 gnd.n5343 2.27742
R20596 gnd.n7505 gnd.n7504 2.27742
R20597 gnd.n7505 gnd.n271 2.27742
R20598 gnd.n7505 gnd.n270 2.27742
R20599 gnd.n7505 gnd.n269 2.27742
R20600 gnd.n4669 gnd.n268 2.27742
R20601 gnd.n1539 gnd.n268 2.27742
R20602 gnd.n4656 gnd.n268 2.27742
R20603 gnd.n4652 gnd.n268 2.27742
R20604 gnd.n7470 gnd.n268 2.27742
R20605 gnd.n1175 gnd.n1174 2.27742
R20606 gnd.n1176 gnd.n1175 2.27742
R20607 gnd.n4976 gnd.n1175 2.27742
R20608 gnd.n1193 gnd.n1175 2.27742
R20609 gnd.n2996 gnd.n2995 2.27742
R20610 gnd.n2995 gnd.n2993 2.27742
R20611 gnd.n2995 gnd.n2944 2.27742
R20612 gnd.n2995 gnd.n2943 2.27742
R20613 gnd.n2995 gnd.n2942 2.27742
R20614 gnd.t279 gnd.n5761 2.23109
R20615 gnd.n5909 gnd.t146 2.23109
R20616 gnd.n2911 gnd.t76 2.23109
R20617 gnd.t321 gnd.n3739 2.23109
R20618 gnd.n3924 gnd.t93 2.23109
R20619 gnd.t35 gnd.n257 2.23109
R20620 gnd.n6365 gnd.n6355 1.93989
R20621 gnd.n6333 gnd.n6323 1.93989
R20622 gnd.n6301 gnd.n6291 1.93989
R20623 gnd.n6270 gnd.n6260 1.93989
R20624 gnd.n6238 gnd.n6228 1.93989
R20625 gnd.n6206 gnd.n6196 1.93989
R20626 gnd.n6174 gnd.n6164 1.93989
R20627 gnd.n6143 gnd.n6133 1.93989
R20628 gnd.n3604 gnd.n3603 1.91244
R20629 gnd.n2331 gnd.n2330 1.91244
R20630 gnd.n2246 gnd.n2245 1.91244
R20631 gnd.n3960 gnd.n3959 1.91244
R20632 gnd.n4131 gnd.n4130 1.91244
R20633 gnd.n2066 gnd.n2064 1.91244
R20634 gnd.n5774 gnd.t14 1.59378
R20635 gnd.n5983 gnd.t143 1.59378
R20636 gnd.n6054 gnd.t167 1.59378
R20637 gnd.t165 gnd.n3782 1.59378
R20638 gnd.n2159 gnd.t306 1.59378
R20639 gnd.n3572 gnd.n2381 1.27512
R20640 gnd.n2358 gnd.t276 1.27512
R20641 gnd.t299 gnd.n3702 1.27512
R20642 gnd.n3700 gnd.n3699 1.27512
R20643 gnd.n3734 gnd.n3733 1.27512
R20644 gnd.n3878 gnd.n3877 1.27512
R20645 gnd.n3911 gnd.n3910 1.27512
R20646 gnd.n4039 gnd.n4038 1.27512
R20647 gnd.n4098 gnd.n2116 1.27512
R20648 gnd.n2115 gnd.t296 1.27512
R20649 gnd.n4193 gnd.t255 1.27512
R20650 gnd.n4206 gnd.n4205 1.27512
R20651 gnd.t264 gnd.n1871 1.27512
R20652 gnd.n5571 gnd.n5570 1.16414
R20653 gnd.n6415 gnd.n5189 1.16414
R20654 gnd.n6364 gnd.n6357 1.16414
R20655 gnd.n6332 gnd.n6325 1.16414
R20656 gnd.n6300 gnd.n6293 1.16414
R20657 gnd.n6269 gnd.n6262 1.16414
R20658 gnd.n6237 gnd.n6230 1.16414
R20659 gnd.n6205 gnd.n6198 1.16414
R20660 gnd.n6173 gnd.n6166 1.16414
R20661 gnd.n6142 gnd.n6135 1.16414
R20662 gnd.n2030 gnd.n2029 0.970197
R20663 gnd.n3495 gnd.n2543 0.970197
R20664 gnd.n6348 gnd.n6316 0.962709
R20665 gnd.n6380 gnd.n6348 0.962709
R20666 gnd.n6221 gnd.n6189 0.962709
R20667 gnd.n6253 gnd.n6221 0.962709
R20668 gnd.t316 gnd.n5885 0.956468
R20669 gnd.n5244 gnd.t152 0.956468
R20670 gnd.n3592 gnd.t95 0.956468
R20671 gnd.n4195 gnd.t97 0.956468
R20672 gnd.n5335 gnd.n5333 0.773756
R20673 gnd.n60 gnd.n58 0.773756
R20674 gnd.n5340 gnd.n5339 0.773756
R20675 gnd.n5339 gnd.n5337 0.773756
R20676 gnd.n5337 gnd.n5335 0.773756
R20677 gnd.n5333 gnd.n5331 0.773756
R20678 gnd.n5331 gnd.n5329 0.773756
R20679 gnd.n5329 gnd.n5327 0.773756
R20680 gnd.n54 gnd.n52 0.773756
R20681 gnd.n56 gnd.n54 0.773756
R20682 gnd.n58 gnd.n56 0.773756
R20683 gnd.n62 gnd.n60 0.773756
R20684 gnd.n64 gnd.n62 0.773756
R20685 gnd.n65 gnd.n64 0.773756
R20686 gnd.n2 gnd.n1 0.672012
R20687 gnd.n3 gnd.n2 0.672012
R20688 gnd.n4 gnd.n3 0.672012
R20689 gnd.n5 gnd.n4 0.672012
R20690 gnd.n6 gnd.n5 0.672012
R20691 gnd.n7 gnd.n6 0.672012
R20692 gnd.n8 gnd.n7 0.672012
R20693 gnd.n9 gnd.n8 0.672012
R20694 gnd.n11 gnd.n10 0.672012
R20695 gnd.n12 gnd.n11 0.672012
R20696 gnd.n13 gnd.n12 0.672012
R20697 gnd.n14 gnd.n13 0.672012
R20698 gnd.n15 gnd.n14 0.672012
R20699 gnd.n16 gnd.n15 0.672012
R20700 gnd.n17 gnd.n16 0.672012
R20701 gnd.n18 gnd.n17 0.672012
R20702 gnd gnd.n0 0.665707
R20703 gnd.n2463 gnd.n2462 0.637812
R20704 gnd.n3665 gnd.n3664 0.637812
R20705 gnd.n3664 gnd.t300 0.637812
R20706 gnd.n3748 gnd.n3747 0.637812
R20707 gnd.n3842 gnd.n3840 0.637812
R20708 gnd.n3859 gnd.t45 0.637812
R20709 gnd.n3933 gnd.t301 0.637812
R20710 gnd.n3926 gnd.n3925 0.637812
R20711 gnd.n4004 gnd.n4003 0.637812
R20712 gnd.n4070 gnd.t294 0.637812
R20713 gnd.n4070 gnd.n4069 0.637812
R20714 gnd.n4168 gnd.n4167 0.637812
R20715 gnd.t238 gnd.n2063 0.637812
R20716 gnd.n5309 gnd.n5308 0.573776
R20717 gnd.n5308 gnd.n5306 0.573776
R20718 gnd.n5306 gnd.n5304 0.573776
R20719 gnd.n5304 gnd.n5302 0.573776
R20720 gnd.n5302 gnd.n5300 0.573776
R20721 gnd.n5300 gnd.n5298 0.573776
R20722 gnd.n5298 gnd.n5296 0.573776
R20723 gnd.n5324 gnd.n5323 0.573776
R20724 gnd.n5323 gnd.n5321 0.573776
R20725 gnd.n5321 gnd.n5319 0.573776
R20726 gnd.n5319 gnd.n5317 0.573776
R20727 gnd.n5317 gnd.n5315 0.573776
R20728 gnd.n5315 gnd.n5313 0.573776
R20729 gnd.n5313 gnd.n5311 0.573776
R20730 gnd.n23 gnd.n21 0.573776
R20731 gnd.n25 gnd.n23 0.573776
R20732 gnd.n27 gnd.n25 0.573776
R20733 gnd.n29 gnd.n27 0.573776
R20734 gnd.n31 gnd.n29 0.573776
R20735 gnd.n33 gnd.n31 0.573776
R20736 gnd.n34 gnd.n33 0.573776
R20737 gnd.n38 gnd.n36 0.573776
R20738 gnd.n40 gnd.n38 0.573776
R20739 gnd.n42 gnd.n40 0.573776
R20740 gnd.n44 gnd.n42 0.573776
R20741 gnd.n46 gnd.n44 0.573776
R20742 gnd.n48 gnd.n46 0.573776
R20743 gnd.n49 gnd.n48 0.573776
R20744 gnd.n7787 gnd.n7786 0.553847
R20745 gnd.n7505 gnd.n268 0.548625
R20746 gnd.n2995 gnd.n1175 0.548625
R20747 gnd.n3048 gnd.n3046 0.505073
R20748 gnd.n3086 gnd.n3085 0.505073
R20749 gnd.n7646 gnd.n7645 0.505073
R20750 gnd.n7617 gnd.n102 0.505073
R20751 gnd.n7740 gnd.n7739 0.492878
R20752 gnd.n7669 gnd.n7668 0.492878
R20753 gnd.n1988 gnd.n1982 0.492878
R20754 gnd.n1907 gnd.n1906 0.492878
R20755 gnd.n2564 gnd.n1318 0.492878
R20756 gnd.n3455 gnd.n3454 0.492878
R20757 gnd.n5062 gnd.n1056 0.492878
R20758 gnd.n3095 gnd.n1013 0.492878
R20759 gnd.n6403 gnd.n5193 0.486781
R20760 gnd.n1693 gnd.n1453 0.486781
R20761 gnd.n5623 gnd.n5519 0.48678
R20762 gnd.n4895 gnd.n4894 0.485256
R20763 gnd.n6494 gnd.n6493 0.480683
R20764 gnd.n5691 gnd.n5469 0.480683
R20765 gnd.n4458 gnd.n4457 0.451719
R20766 gnd.n3428 gnd.n3427 0.451719
R20767 gnd.n742 gnd.n737 0.447146
R20768 gnd.n7183 gnd.n7182 0.447146
R20769 gnd.n7394 gnd.n321 0.447146
R20770 gnd.n2926 gnd.n2925 0.447146
R20771 gnd.n4897 gnd.n4896 0.406268
R20772 gnd.n1692 gnd.n1691 0.404992
R20773 gnd.n3435 gnd.n2658 0.388379
R20774 gnd.n6361 gnd.n6360 0.388379
R20775 gnd.n6329 gnd.n6328 0.388379
R20776 gnd.n6297 gnd.n6296 0.388379
R20777 gnd.n6266 gnd.n6265 0.388379
R20778 gnd.n6234 gnd.n6233 0.388379
R20779 gnd.n6202 gnd.n6201 0.388379
R20780 gnd.n6170 gnd.n6169 0.388379
R20781 gnd.n6139 gnd.n6138 0.388379
R20782 gnd.n7709 gnd.n7708 0.388379
R20783 gnd.n5103 gnd.n5102 0.388379
R20784 gnd.n1791 gnd.n1787 0.388379
R20785 gnd.n7787 gnd.n19 0.374463
R20786 gnd gnd.n7787 0.367492
R20787 gnd.n6103 gnd.t149 0.319156
R20788 gnd.n3783 gnd.t165 0.319156
R20789 gnd.t18 gnd.t10 0.319156
R20790 gnd.t120 gnd.t117 0.319156
R20791 gnd.t306 gnd.n2158 0.319156
R20792 gnd.n5617 gnd.n5616 0.311721
R20793 gnd.n3446 gnd.n3445 0.27489
R20794 gnd.n4481 gnd.n1643 0.27489
R20795 gnd.n6460 gnd.n6459 0.268793
R20796 gnd.n6459 gnd.n6458 0.241354
R20797 gnd.n1947 gnd.n1946 0.229039
R20798 gnd.n1950 gnd.n1947 0.229039
R20799 gnd.n3494 gnd.n2548 0.229039
R20800 gnd.n3494 gnd.n3493 0.229039
R20801 gnd.n5746 gnd.n5487 0.206293
R20802 gnd.n5342 gnd.n0 0.169152
R20803 gnd.n6378 gnd.n6350 0.155672
R20804 gnd.n6371 gnd.n6350 0.155672
R20805 gnd.n6371 gnd.n6370 0.155672
R20806 gnd.n6370 gnd.n6354 0.155672
R20807 gnd.n6363 gnd.n6354 0.155672
R20808 gnd.n6363 gnd.n6362 0.155672
R20809 gnd.n6346 gnd.n6318 0.155672
R20810 gnd.n6339 gnd.n6318 0.155672
R20811 gnd.n6339 gnd.n6338 0.155672
R20812 gnd.n6338 gnd.n6322 0.155672
R20813 gnd.n6331 gnd.n6322 0.155672
R20814 gnd.n6331 gnd.n6330 0.155672
R20815 gnd.n6314 gnd.n6286 0.155672
R20816 gnd.n6307 gnd.n6286 0.155672
R20817 gnd.n6307 gnd.n6306 0.155672
R20818 gnd.n6306 gnd.n6290 0.155672
R20819 gnd.n6299 gnd.n6290 0.155672
R20820 gnd.n6299 gnd.n6298 0.155672
R20821 gnd.n6283 gnd.n6255 0.155672
R20822 gnd.n6276 gnd.n6255 0.155672
R20823 gnd.n6276 gnd.n6275 0.155672
R20824 gnd.n6275 gnd.n6259 0.155672
R20825 gnd.n6268 gnd.n6259 0.155672
R20826 gnd.n6268 gnd.n6267 0.155672
R20827 gnd.n6251 gnd.n6223 0.155672
R20828 gnd.n6244 gnd.n6223 0.155672
R20829 gnd.n6244 gnd.n6243 0.155672
R20830 gnd.n6243 gnd.n6227 0.155672
R20831 gnd.n6236 gnd.n6227 0.155672
R20832 gnd.n6236 gnd.n6235 0.155672
R20833 gnd.n6219 gnd.n6191 0.155672
R20834 gnd.n6212 gnd.n6191 0.155672
R20835 gnd.n6212 gnd.n6211 0.155672
R20836 gnd.n6211 gnd.n6195 0.155672
R20837 gnd.n6204 gnd.n6195 0.155672
R20838 gnd.n6204 gnd.n6203 0.155672
R20839 gnd.n6187 gnd.n6159 0.155672
R20840 gnd.n6180 gnd.n6159 0.155672
R20841 gnd.n6180 gnd.n6179 0.155672
R20842 gnd.n6179 gnd.n6163 0.155672
R20843 gnd.n6172 gnd.n6163 0.155672
R20844 gnd.n6172 gnd.n6171 0.155672
R20845 gnd.n6156 gnd.n6128 0.155672
R20846 gnd.n6149 gnd.n6128 0.155672
R20847 gnd.n6149 gnd.n6148 0.155672
R20848 gnd.n6148 gnd.n6132 0.155672
R20849 gnd.n6141 gnd.n6132 0.155672
R20850 gnd.n6141 gnd.n6140 0.155672
R20851 gnd.n6493 gnd.n963 0.152939
R20852 gnd.n5147 gnd.n963 0.152939
R20853 gnd.n5148 gnd.n5147 0.152939
R20854 gnd.n5149 gnd.n5148 0.152939
R20855 gnd.n5150 gnd.n5149 0.152939
R20856 gnd.n5151 gnd.n5150 0.152939
R20857 gnd.n5152 gnd.n5151 0.152939
R20858 gnd.n5153 gnd.n5152 0.152939
R20859 gnd.n5154 gnd.n5153 0.152939
R20860 gnd.n5155 gnd.n5154 0.152939
R20861 gnd.n5156 gnd.n5155 0.152939
R20862 gnd.n5157 gnd.n5156 0.152939
R20863 gnd.n5158 gnd.n5157 0.152939
R20864 gnd.n5159 gnd.n5158 0.152939
R20865 gnd.n6461 gnd.n5159 0.152939
R20866 gnd.n6461 gnd.n6460 0.152939
R20867 gnd.n5765 gnd.n5469 0.152939
R20868 gnd.n5766 gnd.n5765 0.152939
R20869 gnd.n5767 gnd.n5766 0.152939
R20870 gnd.n5767 gnd.n5448 0.152939
R20871 gnd.n5795 gnd.n5448 0.152939
R20872 gnd.n5796 gnd.n5795 0.152939
R20873 gnd.n5797 gnd.n5796 0.152939
R20874 gnd.n5798 gnd.n5797 0.152939
R20875 gnd.n5798 gnd.n5422 0.152939
R20876 gnd.n5829 gnd.n5422 0.152939
R20877 gnd.n5830 gnd.n5829 0.152939
R20878 gnd.n5831 gnd.n5830 0.152939
R20879 gnd.n5832 gnd.n5831 0.152939
R20880 gnd.n5833 gnd.n5832 0.152939
R20881 gnd.n5833 gnd.n5389 0.152939
R20882 gnd.n5890 gnd.n5389 0.152939
R20883 gnd.n5891 gnd.n5890 0.152939
R20884 gnd.n5892 gnd.n5891 0.152939
R20885 gnd.n5893 gnd.n5892 0.152939
R20886 gnd.n5893 gnd.n5362 0.152939
R20887 gnd.n5930 gnd.n5362 0.152939
R20888 gnd.n5931 gnd.n5930 0.152939
R20889 gnd.n5932 gnd.n5931 0.152939
R20890 gnd.n5933 gnd.n5932 0.152939
R20891 gnd.n5933 gnd.n5287 0.152939
R20892 gnd.n5975 gnd.n5287 0.152939
R20893 gnd.n5976 gnd.n5975 0.152939
R20894 gnd.n5977 gnd.n5976 0.152939
R20895 gnd.n5978 gnd.n5977 0.152939
R20896 gnd.n5978 gnd.n5259 0.152939
R20897 gnd.n6014 gnd.n5259 0.152939
R20898 gnd.n6015 gnd.n6014 0.152939
R20899 gnd.n6016 gnd.n6015 0.152939
R20900 gnd.n6017 gnd.n6016 0.152939
R20901 gnd.n6018 gnd.n6017 0.152939
R20902 gnd.n6018 gnd.n5228 0.152939
R20903 gnd.n6069 gnd.n5228 0.152939
R20904 gnd.n6070 gnd.n6069 0.152939
R20905 gnd.n6071 gnd.n6070 0.152939
R20906 gnd.n6073 gnd.n6071 0.152939
R20907 gnd.n6073 gnd.n6072 0.152939
R20908 gnd.n6072 gnd.n913 0.152939
R20909 gnd.n914 gnd.n913 0.152939
R20910 gnd.n915 gnd.n914 0.152939
R20911 gnd.n935 gnd.n915 0.152939
R20912 gnd.n936 gnd.n935 0.152939
R20913 gnd.n937 gnd.n936 0.152939
R20914 gnd.n938 gnd.n937 0.152939
R20915 gnd.n939 gnd.n938 0.152939
R20916 gnd.n960 gnd.n939 0.152939
R20917 gnd.n961 gnd.n960 0.152939
R20918 gnd.n962 gnd.n961 0.152939
R20919 gnd.n6494 gnd.n962 0.152939
R20920 gnd.n5692 gnd.n5691 0.152939
R20921 gnd.n5693 gnd.n5692 0.152939
R20922 gnd.n5694 gnd.n5693 0.152939
R20923 gnd.n5695 gnd.n5694 0.152939
R20924 gnd.n5696 gnd.n5695 0.152939
R20925 gnd.n5697 gnd.n5696 0.152939
R20926 gnd.n5698 gnd.n5697 0.152939
R20927 gnd.n5699 gnd.n5698 0.152939
R20928 gnd.n5700 gnd.n5699 0.152939
R20929 gnd.n5701 gnd.n5700 0.152939
R20930 gnd.n5702 gnd.n5701 0.152939
R20931 gnd.n5703 gnd.n5702 0.152939
R20932 gnd.n5704 gnd.n5703 0.152939
R20933 gnd.n5705 gnd.n5704 0.152939
R20934 gnd.n5709 gnd.n5705 0.152939
R20935 gnd.n5709 gnd.n5487 0.152939
R20936 gnd.n6458 gnd.n5164 0.152939
R20937 gnd.n5166 gnd.n5164 0.152939
R20938 gnd.n5167 gnd.n5166 0.152939
R20939 gnd.n5168 gnd.n5167 0.152939
R20940 gnd.n5169 gnd.n5168 0.152939
R20941 gnd.n5170 gnd.n5169 0.152939
R20942 gnd.n5171 gnd.n5170 0.152939
R20943 gnd.n5172 gnd.n5171 0.152939
R20944 gnd.n5173 gnd.n5172 0.152939
R20945 gnd.n5174 gnd.n5173 0.152939
R20946 gnd.n5175 gnd.n5174 0.152939
R20947 gnd.n5176 gnd.n5175 0.152939
R20948 gnd.n5177 gnd.n5176 0.152939
R20949 gnd.n5178 gnd.n5177 0.152939
R20950 gnd.n5179 gnd.n5178 0.152939
R20951 gnd.n5180 gnd.n5179 0.152939
R20952 gnd.n5181 gnd.n5180 0.152939
R20953 gnd.n5182 gnd.n5181 0.152939
R20954 gnd.n5183 gnd.n5182 0.152939
R20955 gnd.n5184 gnd.n5183 0.152939
R20956 gnd.n5185 gnd.n5184 0.152939
R20957 gnd.n5186 gnd.n5185 0.152939
R20958 gnd.n5190 gnd.n5186 0.152939
R20959 gnd.n5191 gnd.n5190 0.152939
R20960 gnd.n5192 gnd.n5191 0.152939
R20961 gnd.n5193 gnd.n5192 0.152939
R20962 gnd.n5952 gnd.n5951 0.152939
R20963 gnd.n5953 gnd.n5952 0.152939
R20964 gnd.n5954 gnd.n5953 0.152939
R20965 gnd.n5955 gnd.n5954 0.152939
R20966 gnd.n5956 gnd.n5955 0.152939
R20967 gnd.n5957 gnd.n5956 0.152939
R20968 gnd.n5958 gnd.n5957 0.152939
R20969 gnd.n5959 gnd.n5958 0.152939
R20970 gnd.n5959 gnd.n5240 0.152939
R20971 gnd.n6037 gnd.n5240 0.152939
R20972 gnd.n6038 gnd.n6037 0.152939
R20973 gnd.n6039 gnd.n6038 0.152939
R20974 gnd.n6040 gnd.n6039 0.152939
R20975 gnd.n6041 gnd.n6040 0.152939
R20976 gnd.n6042 gnd.n6041 0.152939
R20977 gnd.n6043 gnd.n6042 0.152939
R20978 gnd.n6044 gnd.n6043 0.152939
R20979 gnd.n6044 gnd.n5206 0.152939
R20980 gnd.n6106 gnd.n5206 0.152939
R20981 gnd.n6107 gnd.n6106 0.152939
R20982 gnd.n6108 gnd.n6107 0.152939
R20983 gnd.n6109 gnd.n6108 0.152939
R20984 gnd.n6110 gnd.n6109 0.152939
R20985 gnd.n6111 gnd.n6110 0.152939
R20986 gnd.n6111 gnd.n5195 0.152939
R20987 gnd.n6401 gnd.n5195 0.152939
R20988 gnd.n6402 gnd.n6401 0.152939
R20989 gnd.n6403 gnd.n6402 0.152939
R20990 gnd.n5624 gnd.n5623 0.152939
R20991 gnd.n5625 gnd.n5624 0.152939
R20992 gnd.n5625 gnd.n5507 0.152939
R20993 gnd.n5639 gnd.n5507 0.152939
R20994 gnd.n5640 gnd.n5639 0.152939
R20995 gnd.n5641 gnd.n5640 0.152939
R20996 gnd.n5641 gnd.n5494 0.152939
R20997 gnd.n5655 gnd.n5494 0.152939
R20998 gnd.n5656 gnd.n5655 0.152939
R20999 gnd.n5657 gnd.n5656 0.152939
R21000 gnd.n5658 gnd.n5657 0.152939
R21001 gnd.n5659 gnd.n5658 0.152939
R21002 gnd.n5660 gnd.n5659 0.152939
R21003 gnd.n5661 gnd.n5660 0.152939
R21004 gnd.n5662 gnd.n5661 0.152939
R21005 gnd.n5663 gnd.n5662 0.152939
R21006 gnd.n5664 gnd.n5663 0.152939
R21007 gnd.n5665 gnd.n5664 0.152939
R21008 gnd.n5666 gnd.n5665 0.152939
R21009 gnd.n5666 gnd.n5429 0.152939
R21010 gnd.n5818 gnd.n5429 0.152939
R21011 gnd.n5819 gnd.n5818 0.152939
R21012 gnd.n5820 gnd.n5819 0.152939
R21013 gnd.n5821 gnd.n5820 0.152939
R21014 gnd.n5821 gnd.n5396 0.152939
R21015 gnd.n5865 gnd.n5396 0.152939
R21016 gnd.n5866 gnd.n5865 0.152939
R21017 gnd.n5867 gnd.n5866 0.152939
R21018 gnd.n5616 gnd.n5523 0.152939
R21019 gnd.n5526 gnd.n5523 0.152939
R21020 gnd.n5527 gnd.n5526 0.152939
R21021 gnd.n5528 gnd.n5527 0.152939
R21022 gnd.n5531 gnd.n5528 0.152939
R21023 gnd.n5532 gnd.n5531 0.152939
R21024 gnd.n5533 gnd.n5532 0.152939
R21025 gnd.n5534 gnd.n5533 0.152939
R21026 gnd.n5537 gnd.n5534 0.152939
R21027 gnd.n5538 gnd.n5537 0.152939
R21028 gnd.n5539 gnd.n5538 0.152939
R21029 gnd.n5540 gnd.n5539 0.152939
R21030 gnd.n5543 gnd.n5540 0.152939
R21031 gnd.n5544 gnd.n5543 0.152939
R21032 gnd.n5545 gnd.n5544 0.152939
R21033 gnd.n5546 gnd.n5545 0.152939
R21034 gnd.n5549 gnd.n5546 0.152939
R21035 gnd.n5550 gnd.n5549 0.152939
R21036 gnd.n5551 gnd.n5550 0.152939
R21037 gnd.n5552 gnd.n5551 0.152939
R21038 gnd.n5555 gnd.n5552 0.152939
R21039 gnd.n5556 gnd.n5555 0.152939
R21040 gnd.n5559 gnd.n5556 0.152939
R21041 gnd.n5560 gnd.n5559 0.152939
R21042 gnd.n5562 gnd.n5560 0.152939
R21043 gnd.n5562 gnd.n5519 0.152939
R21044 gnd.n6700 gnd.n737 0.152939
R21045 gnd.n6701 gnd.n6700 0.152939
R21046 gnd.n6702 gnd.n6701 0.152939
R21047 gnd.n6702 gnd.n731 0.152939
R21048 gnd.n6710 gnd.n731 0.152939
R21049 gnd.n6711 gnd.n6710 0.152939
R21050 gnd.n6712 gnd.n6711 0.152939
R21051 gnd.n6712 gnd.n725 0.152939
R21052 gnd.n6720 gnd.n725 0.152939
R21053 gnd.n6721 gnd.n6720 0.152939
R21054 gnd.n6722 gnd.n6721 0.152939
R21055 gnd.n6722 gnd.n719 0.152939
R21056 gnd.n6730 gnd.n719 0.152939
R21057 gnd.n6731 gnd.n6730 0.152939
R21058 gnd.n6732 gnd.n6731 0.152939
R21059 gnd.n6732 gnd.n713 0.152939
R21060 gnd.n6740 gnd.n713 0.152939
R21061 gnd.n6741 gnd.n6740 0.152939
R21062 gnd.n6742 gnd.n6741 0.152939
R21063 gnd.n6742 gnd.n707 0.152939
R21064 gnd.n6750 gnd.n707 0.152939
R21065 gnd.n6751 gnd.n6750 0.152939
R21066 gnd.n6752 gnd.n6751 0.152939
R21067 gnd.n6752 gnd.n701 0.152939
R21068 gnd.n6760 gnd.n701 0.152939
R21069 gnd.n6761 gnd.n6760 0.152939
R21070 gnd.n6762 gnd.n6761 0.152939
R21071 gnd.n6762 gnd.n695 0.152939
R21072 gnd.n6770 gnd.n695 0.152939
R21073 gnd.n6771 gnd.n6770 0.152939
R21074 gnd.n6772 gnd.n6771 0.152939
R21075 gnd.n6772 gnd.n689 0.152939
R21076 gnd.n6780 gnd.n689 0.152939
R21077 gnd.n6781 gnd.n6780 0.152939
R21078 gnd.n6782 gnd.n6781 0.152939
R21079 gnd.n6782 gnd.n683 0.152939
R21080 gnd.n6790 gnd.n683 0.152939
R21081 gnd.n6791 gnd.n6790 0.152939
R21082 gnd.n6792 gnd.n6791 0.152939
R21083 gnd.n6792 gnd.n677 0.152939
R21084 gnd.n6800 gnd.n677 0.152939
R21085 gnd.n6801 gnd.n6800 0.152939
R21086 gnd.n6802 gnd.n6801 0.152939
R21087 gnd.n6802 gnd.n671 0.152939
R21088 gnd.n6810 gnd.n671 0.152939
R21089 gnd.n6811 gnd.n6810 0.152939
R21090 gnd.n6812 gnd.n6811 0.152939
R21091 gnd.n6812 gnd.n665 0.152939
R21092 gnd.n6820 gnd.n665 0.152939
R21093 gnd.n6821 gnd.n6820 0.152939
R21094 gnd.n6822 gnd.n6821 0.152939
R21095 gnd.n6822 gnd.n659 0.152939
R21096 gnd.n6830 gnd.n659 0.152939
R21097 gnd.n6831 gnd.n6830 0.152939
R21098 gnd.n6832 gnd.n6831 0.152939
R21099 gnd.n6832 gnd.n653 0.152939
R21100 gnd.n6840 gnd.n653 0.152939
R21101 gnd.n6841 gnd.n6840 0.152939
R21102 gnd.n6842 gnd.n6841 0.152939
R21103 gnd.n6842 gnd.n647 0.152939
R21104 gnd.n6850 gnd.n647 0.152939
R21105 gnd.n6851 gnd.n6850 0.152939
R21106 gnd.n6852 gnd.n6851 0.152939
R21107 gnd.n6852 gnd.n641 0.152939
R21108 gnd.n6860 gnd.n641 0.152939
R21109 gnd.n6861 gnd.n6860 0.152939
R21110 gnd.n6862 gnd.n6861 0.152939
R21111 gnd.n6862 gnd.n635 0.152939
R21112 gnd.n6870 gnd.n635 0.152939
R21113 gnd.n6871 gnd.n6870 0.152939
R21114 gnd.n6872 gnd.n6871 0.152939
R21115 gnd.n6872 gnd.n629 0.152939
R21116 gnd.n6880 gnd.n629 0.152939
R21117 gnd.n6881 gnd.n6880 0.152939
R21118 gnd.n6882 gnd.n6881 0.152939
R21119 gnd.n6882 gnd.n623 0.152939
R21120 gnd.n6890 gnd.n623 0.152939
R21121 gnd.n6891 gnd.n6890 0.152939
R21122 gnd.n6892 gnd.n6891 0.152939
R21123 gnd.n6892 gnd.n617 0.152939
R21124 gnd.n6900 gnd.n617 0.152939
R21125 gnd.n6901 gnd.n6900 0.152939
R21126 gnd.n6902 gnd.n6901 0.152939
R21127 gnd.n6902 gnd.n611 0.152939
R21128 gnd.n6910 gnd.n611 0.152939
R21129 gnd.n6911 gnd.n6910 0.152939
R21130 gnd.n6912 gnd.n6911 0.152939
R21131 gnd.n6912 gnd.n605 0.152939
R21132 gnd.n6920 gnd.n605 0.152939
R21133 gnd.n6921 gnd.n6920 0.152939
R21134 gnd.n6922 gnd.n6921 0.152939
R21135 gnd.n6922 gnd.n599 0.152939
R21136 gnd.n6930 gnd.n599 0.152939
R21137 gnd.n6931 gnd.n6930 0.152939
R21138 gnd.n6932 gnd.n6931 0.152939
R21139 gnd.n6932 gnd.n593 0.152939
R21140 gnd.n6940 gnd.n593 0.152939
R21141 gnd.n6941 gnd.n6940 0.152939
R21142 gnd.n6942 gnd.n6941 0.152939
R21143 gnd.n6942 gnd.n587 0.152939
R21144 gnd.n6950 gnd.n587 0.152939
R21145 gnd.n6951 gnd.n6950 0.152939
R21146 gnd.n6952 gnd.n6951 0.152939
R21147 gnd.n6952 gnd.n581 0.152939
R21148 gnd.n6960 gnd.n581 0.152939
R21149 gnd.n6961 gnd.n6960 0.152939
R21150 gnd.n6962 gnd.n6961 0.152939
R21151 gnd.n6962 gnd.n575 0.152939
R21152 gnd.n6970 gnd.n575 0.152939
R21153 gnd.n6971 gnd.n6970 0.152939
R21154 gnd.n6972 gnd.n6971 0.152939
R21155 gnd.n6972 gnd.n569 0.152939
R21156 gnd.n6980 gnd.n569 0.152939
R21157 gnd.n6981 gnd.n6980 0.152939
R21158 gnd.n6982 gnd.n6981 0.152939
R21159 gnd.n6982 gnd.n563 0.152939
R21160 gnd.n6990 gnd.n563 0.152939
R21161 gnd.n6991 gnd.n6990 0.152939
R21162 gnd.n6992 gnd.n6991 0.152939
R21163 gnd.n6992 gnd.n557 0.152939
R21164 gnd.n7000 gnd.n557 0.152939
R21165 gnd.n7001 gnd.n7000 0.152939
R21166 gnd.n7002 gnd.n7001 0.152939
R21167 gnd.n7002 gnd.n551 0.152939
R21168 gnd.n7010 gnd.n551 0.152939
R21169 gnd.n7011 gnd.n7010 0.152939
R21170 gnd.n7012 gnd.n7011 0.152939
R21171 gnd.n7012 gnd.n545 0.152939
R21172 gnd.n7020 gnd.n545 0.152939
R21173 gnd.n7021 gnd.n7020 0.152939
R21174 gnd.n7022 gnd.n7021 0.152939
R21175 gnd.n7022 gnd.n539 0.152939
R21176 gnd.n7030 gnd.n539 0.152939
R21177 gnd.n7031 gnd.n7030 0.152939
R21178 gnd.n7032 gnd.n7031 0.152939
R21179 gnd.n7032 gnd.n533 0.152939
R21180 gnd.n7040 gnd.n533 0.152939
R21181 gnd.n7041 gnd.n7040 0.152939
R21182 gnd.n7042 gnd.n7041 0.152939
R21183 gnd.n7042 gnd.n527 0.152939
R21184 gnd.n7050 gnd.n527 0.152939
R21185 gnd.n7051 gnd.n7050 0.152939
R21186 gnd.n7052 gnd.n7051 0.152939
R21187 gnd.n7052 gnd.n521 0.152939
R21188 gnd.n7060 gnd.n521 0.152939
R21189 gnd.n7061 gnd.n7060 0.152939
R21190 gnd.n7062 gnd.n7061 0.152939
R21191 gnd.n7062 gnd.n515 0.152939
R21192 gnd.n7070 gnd.n515 0.152939
R21193 gnd.n7071 gnd.n7070 0.152939
R21194 gnd.n7072 gnd.n7071 0.152939
R21195 gnd.n7072 gnd.n509 0.152939
R21196 gnd.n7080 gnd.n509 0.152939
R21197 gnd.n7081 gnd.n7080 0.152939
R21198 gnd.n7082 gnd.n7081 0.152939
R21199 gnd.n7082 gnd.n503 0.152939
R21200 gnd.n7090 gnd.n503 0.152939
R21201 gnd.n7091 gnd.n7090 0.152939
R21202 gnd.n7092 gnd.n7091 0.152939
R21203 gnd.n7092 gnd.n497 0.152939
R21204 gnd.n7100 gnd.n497 0.152939
R21205 gnd.n7101 gnd.n7100 0.152939
R21206 gnd.n7102 gnd.n7101 0.152939
R21207 gnd.n7102 gnd.n491 0.152939
R21208 gnd.n7110 gnd.n491 0.152939
R21209 gnd.n7111 gnd.n7110 0.152939
R21210 gnd.n7112 gnd.n7111 0.152939
R21211 gnd.n7112 gnd.n485 0.152939
R21212 gnd.n7120 gnd.n485 0.152939
R21213 gnd.n7121 gnd.n7120 0.152939
R21214 gnd.n7122 gnd.n7121 0.152939
R21215 gnd.n7122 gnd.n479 0.152939
R21216 gnd.n7130 gnd.n479 0.152939
R21217 gnd.n7131 gnd.n7130 0.152939
R21218 gnd.n7132 gnd.n7131 0.152939
R21219 gnd.n7132 gnd.n473 0.152939
R21220 gnd.n7140 gnd.n473 0.152939
R21221 gnd.n7141 gnd.n7140 0.152939
R21222 gnd.n7142 gnd.n7141 0.152939
R21223 gnd.n7142 gnd.n467 0.152939
R21224 gnd.n7150 gnd.n467 0.152939
R21225 gnd.n7151 gnd.n7150 0.152939
R21226 gnd.n7152 gnd.n7151 0.152939
R21227 gnd.n7152 gnd.n461 0.152939
R21228 gnd.n7160 gnd.n461 0.152939
R21229 gnd.n7161 gnd.n7160 0.152939
R21230 gnd.n7162 gnd.n7161 0.152939
R21231 gnd.n7162 gnd.n455 0.152939
R21232 gnd.n7170 gnd.n455 0.152939
R21233 gnd.n7171 gnd.n7170 0.152939
R21234 gnd.n7173 gnd.n7171 0.152939
R21235 gnd.n7173 gnd.n7172 0.152939
R21236 gnd.n7172 gnd.n449 0.152939
R21237 gnd.n7182 gnd.n449 0.152939
R21238 gnd.n7183 gnd.n444 0.152939
R21239 gnd.n7191 gnd.n444 0.152939
R21240 gnd.n7192 gnd.n7191 0.152939
R21241 gnd.n7193 gnd.n7192 0.152939
R21242 gnd.n7193 gnd.n438 0.152939
R21243 gnd.n7201 gnd.n438 0.152939
R21244 gnd.n7202 gnd.n7201 0.152939
R21245 gnd.n7203 gnd.n7202 0.152939
R21246 gnd.n7203 gnd.n432 0.152939
R21247 gnd.n7211 gnd.n432 0.152939
R21248 gnd.n7212 gnd.n7211 0.152939
R21249 gnd.n7213 gnd.n7212 0.152939
R21250 gnd.n7213 gnd.n426 0.152939
R21251 gnd.n7221 gnd.n426 0.152939
R21252 gnd.n7222 gnd.n7221 0.152939
R21253 gnd.n7223 gnd.n7222 0.152939
R21254 gnd.n7223 gnd.n420 0.152939
R21255 gnd.n7231 gnd.n420 0.152939
R21256 gnd.n7232 gnd.n7231 0.152939
R21257 gnd.n7233 gnd.n7232 0.152939
R21258 gnd.n7233 gnd.n414 0.152939
R21259 gnd.n7241 gnd.n414 0.152939
R21260 gnd.n7242 gnd.n7241 0.152939
R21261 gnd.n7243 gnd.n7242 0.152939
R21262 gnd.n7243 gnd.n408 0.152939
R21263 gnd.n7251 gnd.n408 0.152939
R21264 gnd.n7252 gnd.n7251 0.152939
R21265 gnd.n7253 gnd.n7252 0.152939
R21266 gnd.n7253 gnd.n402 0.152939
R21267 gnd.n7261 gnd.n402 0.152939
R21268 gnd.n7262 gnd.n7261 0.152939
R21269 gnd.n7263 gnd.n7262 0.152939
R21270 gnd.n7263 gnd.n396 0.152939
R21271 gnd.n7271 gnd.n396 0.152939
R21272 gnd.n7272 gnd.n7271 0.152939
R21273 gnd.n7273 gnd.n7272 0.152939
R21274 gnd.n7273 gnd.n390 0.152939
R21275 gnd.n7281 gnd.n390 0.152939
R21276 gnd.n7282 gnd.n7281 0.152939
R21277 gnd.n7283 gnd.n7282 0.152939
R21278 gnd.n7283 gnd.n384 0.152939
R21279 gnd.n7291 gnd.n384 0.152939
R21280 gnd.n7292 gnd.n7291 0.152939
R21281 gnd.n7293 gnd.n7292 0.152939
R21282 gnd.n7293 gnd.n378 0.152939
R21283 gnd.n7301 gnd.n378 0.152939
R21284 gnd.n7302 gnd.n7301 0.152939
R21285 gnd.n7303 gnd.n7302 0.152939
R21286 gnd.n7303 gnd.n372 0.152939
R21287 gnd.n7311 gnd.n372 0.152939
R21288 gnd.n7312 gnd.n7311 0.152939
R21289 gnd.n7313 gnd.n7312 0.152939
R21290 gnd.n7313 gnd.n366 0.152939
R21291 gnd.n7321 gnd.n366 0.152939
R21292 gnd.n7322 gnd.n7321 0.152939
R21293 gnd.n7323 gnd.n7322 0.152939
R21294 gnd.n7323 gnd.n360 0.152939
R21295 gnd.n7331 gnd.n360 0.152939
R21296 gnd.n7332 gnd.n7331 0.152939
R21297 gnd.n7333 gnd.n7332 0.152939
R21298 gnd.n7333 gnd.n354 0.152939
R21299 gnd.n7341 gnd.n354 0.152939
R21300 gnd.n7342 gnd.n7341 0.152939
R21301 gnd.n7343 gnd.n7342 0.152939
R21302 gnd.n7343 gnd.n348 0.152939
R21303 gnd.n7351 gnd.n348 0.152939
R21304 gnd.n7352 gnd.n7351 0.152939
R21305 gnd.n7353 gnd.n7352 0.152939
R21306 gnd.n7353 gnd.n342 0.152939
R21307 gnd.n7361 gnd.n342 0.152939
R21308 gnd.n7362 gnd.n7361 0.152939
R21309 gnd.n7363 gnd.n7362 0.152939
R21310 gnd.n7363 gnd.n336 0.152939
R21311 gnd.n7371 gnd.n336 0.152939
R21312 gnd.n7372 gnd.n7371 0.152939
R21313 gnd.n7373 gnd.n7372 0.152939
R21314 gnd.n7373 gnd.n330 0.152939
R21315 gnd.n7381 gnd.n330 0.152939
R21316 gnd.n7382 gnd.n7381 0.152939
R21317 gnd.n7383 gnd.n7382 0.152939
R21318 gnd.n7383 gnd.n324 0.152939
R21319 gnd.n7392 gnd.n324 0.152939
R21320 gnd.n7393 gnd.n7392 0.152939
R21321 gnd.n7394 gnd.n7393 0.152939
R21322 gnd.n312 gnd.n309 0.152939
R21323 gnd.n313 gnd.n312 0.152939
R21324 gnd.n314 gnd.n313 0.152939
R21325 gnd.n315 gnd.n314 0.152939
R21326 gnd.n318 gnd.n315 0.152939
R21327 gnd.n319 gnd.n318 0.152939
R21328 gnd.n320 gnd.n319 0.152939
R21329 gnd.n321 gnd.n320 0.152939
R21330 gnd.n7519 gnd.n252 0.152939
R21331 gnd.n7520 gnd.n7519 0.152939
R21332 gnd.n7521 gnd.n7520 0.152939
R21333 gnd.n7521 gnd.n236 0.152939
R21334 gnd.n7535 gnd.n236 0.152939
R21335 gnd.n7536 gnd.n7535 0.152939
R21336 gnd.n7537 gnd.n7536 0.152939
R21337 gnd.n7537 gnd.n222 0.152939
R21338 gnd.n7551 gnd.n222 0.152939
R21339 gnd.n7552 gnd.n7551 0.152939
R21340 gnd.n7553 gnd.n7552 0.152939
R21341 gnd.n7553 gnd.n205 0.152939
R21342 gnd.n7567 gnd.n205 0.152939
R21343 gnd.n7568 gnd.n7567 0.152939
R21344 gnd.n7569 gnd.n7568 0.152939
R21345 gnd.n7569 gnd.n190 0.152939
R21346 gnd.n7658 gnd.n190 0.152939
R21347 gnd.n7659 gnd.n7658 0.152939
R21348 gnd.n7660 gnd.n7659 0.152939
R21349 gnd.n7660 gnd.n111 0.152939
R21350 gnd.n7740 gnd.n111 0.152939
R21351 gnd.n7739 gnd.n112 0.152939
R21352 gnd.n114 gnd.n112 0.152939
R21353 gnd.n119 gnd.n114 0.152939
R21354 gnd.n120 gnd.n119 0.152939
R21355 gnd.n121 gnd.n120 0.152939
R21356 gnd.n122 gnd.n121 0.152939
R21357 gnd.n126 gnd.n122 0.152939
R21358 gnd.n127 gnd.n126 0.152939
R21359 gnd.n128 gnd.n127 0.152939
R21360 gnd.n129 gnd.n128 0.152939
R21361 gnd.n133 gnd.n129 0.152939
R21362 gnd.n134 gnd.n133 0.152939
R21363 gnd.n135 gnd.n134 0.152939
R21364 gnd.n136 gnd.n135 0.152939
R21365 gnd.n140 gnd.n136 0.152939
R21366 gnd.n141 gnd.n140 0.152939
R21367 gnd.n142 gnd.n141 0.152939
R21368 gnd.n143 gnd.n142 0.152939
R21369 gnd.n147 gnd.n143 0.152939
R21370 gnd.n148 gnd.n147 0.152939
R21371 gnd.n149 gnd.n148 0.152939
R21372 gnd.n150 gnd.n149 0.152939
R21373 gnd.n154 gnd.n150 0.152939
R21374 gnd.n155 gnd.n154 0.152939
R21375 gnd.n156 gnd.n155 0.152939
R21376 gnd.n157 gnd.n156 0.152939
R21377 gnd.n161 gnd.n157 0.152939
R21378 gnd.n162 gnd.n161 0.152939
R21379 gnd.n163 gnd.n162 0.152939
R21380 gnd.n164 gnd.n163 0.152939
R21381 gnd.n168 gnd.n164 0.152939
R21382 gnd.n169 gnd.n168 0.152939
R21383 gnd.n170 gnd.n169 0.152939
R21384 gnd.n171 gnd.n170 0.152939
R21385 gnd.n175 gnd.n171 0.152939
R21386 gnd.n176 gnd.n175 0.152939
R21387 gnd.n7670 gnd.n176 0.152939
R21388 gnd.n7670 gnd.n7669 0.152939
R21389 gnd.n1982 gnd.n1981 0.152939
R21390 gnd.n1981 gnd.n1639 0.152939
R21391 gnd.n4491 gnd.n1639 0.152939
R21392 gnd.n4492 gnd.n4491 0.152939
R21393 gnd.n4493 gnd.n4492 0.152939
R21394 gnd.n4494 gnd.n4493 0.152939
R21395 gnd.n4495 gnd.n4494 0.152939
R21396 gnd.n4496 gnd.n4495 0.152939
R21397 gnd.n4497 gnd.n4496 0.152939
R21398 gnd.n4498 gnd.n4497 0.152939
R21399 gnd.n4499 gnd.n4498 0.152939
R21400 gnd.n4500 gnd.n4499 0.152939
R21401 gnd.n4501 gnd.n4500 0.152939
R21402 gnd.n4502 gnd.n4501 0.152939
R21403 gnd.n4504 gnd.n4502 0.152939
R21404 gnd.n4504 gnd.n4503 0.152939
R21405 gnd.n4503 gnd.n1559 0.152939
R21406 gnd.n1559 gnd.n1557 0.152939
R21407 gnd.n4618 gnd.n1557 0.152939
R21408 gnd.n4619 gnd.n4618 0.152939
R21409 gnd.n4620 gnd.n4619 0.152939
R21410 gnd.n4621 gnd.n4620 0.152939
R21411 gnd.n4621 gnd.n1549 0.152939
R21412 gnd.n4641 gnd.n1549 0.152939
R21413 gnd.n4642 gnd.n4641 0.152939
R21414 gnd.n4643 gnd.n4642 0.152939
R21415 gnd.n301 gnd.n300 0.152939
R21416 gnd.n302 gnd.n301 0.152939
R21417 gnd.n303 gnd.n302 0.152939
R21418 gnd.n7405 gnd.n303 0.152939
R21419 gnd.n7409 gnd.n7405 0.152939
R21420 gnd.n7410 gnd.n7409 0.152939
R21421 gnd.n7411 gnd.n7410 0.152939
R21422 gnd.n7411 gnd.n7403 0.152939
R21423 gnd.n7420 gnd.n7403 0.152939
R21424 gnd.n7421 gnd.n7420 0.152939
R21425 gnd.n7422 gnd.n7421 0.152939
R21426 gnd.n7423 gnd.n7422 0.152939
R21427 gnd.n7424 gnd.n7423 0.152939
R21428 gnd.n7425 gnd.n7424 0.152939
R21429 gnd.n7426 gnd.n7425 0.152939
R21430 gnd.n7427 gnd.n7426 0.152939
R21431 gnd.n7428 gnd.n7427 0.152939
R21432 gnd.n7429 gnd.n7428 0.152939
R21433 gnd.n7430 gnd.n7429 0.152939
R21434 gnd.n7431 gnd.n7430 0.152939
R21435 gnd.n7432 gnd.n7431 0.152939
R21436 gnd.n7433 gnd.n7432 0.152939
R21437 gnd.n7435 gnd.n7433 0.152939
R21438 gnd.n7435 gnd.n7434 0.152939
R21439 gnd.n7434 gnd.n182 0.152939
R21440 gnd.n7668 gnd.n182 0.152939
R21441 gnd.n1913 gnd.n1907 0.152939
R21442 gnd.n1914 gnd.n1913 0.152939
R21443 gnd.n1915 gnd.n1914 0.152939
R21444 gnd.n1915 gnd.n1902 0.152939
R21445 gnd.n1923 gnd.n1902 0.152939
R21446 gnd.n1924 gnd.n1923 0.152939
R21447 gnd.n1925 gnd.n1924 0.152939
R21448 gnd.n1925 gnd.n1898 0.152939
R21449 gnd.n1933 gnd.n1898 0.152939
R21450 gnd.n1934 gnd.n1933 0.152939
R21451 gnd.n1936 gnd.n1934 0.152939
R21452 gnd.n1936 gnd.n1935 0.152939
R21453 gnd.n1935 gnd.n1891 0.152939
R21454 gnd.n1945 gnd.n1891 0.152939
R21455 gnd.n1946 gnd.n1945 0.152939
R21456 gnd.n1953 gnd.n1950 0.152939
R21457 gnd.n1954 gnd.n1953 0.152939
R21458 gnd.n1955 gnd.n1954 0.152939
R21459 gnd.n1956 gnd.n1955 0.152939
R21460 gnd.n1959 gnd.n1956 0.152939
R21461 gnd.n1960 gnd.n1959 0.152939
R21462 gnd.n1961 gnd.n1960 0.152939
R21463 gnd.n1962 gnd.n1961 0.152939
R21464 gnd.n1965 gnd.n1962 0.152939
R21465 gnd.n1966 gnd.n1965 0.152939
R21466 gnd.n1967 gnd.n1966 0.152939
R21467 gnd.n1968 gnd.n1967 0.152939
R21468 gnd.n1971 gnd.n1968 0.152939
R21469 gnd.n1972 gnd.n1971 0.152939
R21470 gnd.n1973 gnd.n1972 0.152939
R21471 gnd.n1974 gnd.n1973 0.152939
R21472 gnd.n1980 gnd.n1974 0.152939
R21473 gnd.n1990 gnd.n1980 0.152939
R21474 gnd.n1990 gnd.n1989 0.152939
R21475 gnd.n1989 gnd.n1988 0.152939
R21476 gnd.n1906 gnd.n1485 0.152939
R21477 gnd.n1486 gnd.n1485 0.152939
R21478 gnd.n1487 gnd.n1486 0.152939
R21479 gnd.n4522 gnd.n1487 0.152939
R21480 gnd.n4523 gnd.n4522 0.152939
R21481 gnd.n4524 gnd.n4523 0.152939
R21482 gnd.n4524 gnd.n1602 0.152939
R21483 gnd.n4553 gnd.n1602 0.152939
R21484 gnd.n4554 gnd.n4553 0.152939
R21485 gnd.n4555 gnd.n4554 0.152939
R21486 gnd.n4556 gnd.n4555 0.152939
R21487 gnd.n4556 gnd.n1575 0.152939
R21488 gnd.n4592 gnd.n1575 0.152939
R21489 gnd.n4593 gnd.n4592 0.152939
R21490 gnd.n4594 gnd.n4593 0.152939
R21491 gnd.n4595 gnd.n4594 0.152939
R21492 gnd.n4595 gnd.n1523 0.152939
R21493 gnd.n4682 gnd.n1523 0.152939
R21494 gnd.n4683 gnd.n4682 0.152939
R21495 gnd.n4684 gnd.n4683 0.152939
R21496 gnd.n4684 gnd.n267 0.152939
R21497 gnd.n2947 gnd.n2941 0.152939
R21498 gnd.n2950 gnd.n2947 0.152939
R21499 gnd.n2951 gnd.n2950 0.152939
R21500 gnd.n2952 gnd.n2951 0.152939
R21501 gnd.n2953 gnd.n2952 0.152939
R21502 gnd.n2956 gnd.n2953 0.152939
R21503 gnd.n2957 gnd.n2956 0.152939
R21504 gnd.n2958 gnd.n2957 0.152939
R21505 gnd.n2959 gnd.n2958 0.152939
R21506 gnd.n2960 gnd.n2959 0.152939
R21507 gnd.n2960 gnd.n2855 0.152939
R21508 gnd.n3303 gnd.n2855 0.152939
R21509 gnd.n3304 gnd.n3303 0.152939
R21510 gnd.n3305 gnd.n3304 0.152939
R21511 gnd.n3305 gnd.n2851 0.152939
R21512 gnd.n3311 gnd.n2851 0.152939
R21513 gnd.n3312 gnd.n3311 0.152939
R21514 gnd.n3313 gnd.n3312 0.152939
R21515 gnd.n3313 gnd.n2847 0.152939
R21516 gnd.n3319 gnd.n2847 0.152939
R21517 gnd.n3320 gnd.n3319 0.152939
R21518 gnd.n3321 gnd.n3320 0.152939
R21519 gnd.n3321 gnd.n2843 0.152939
R21520 gnd.n3330 gnd.n2843 0.152939
R21521 gnd.n3331 gnd.n3330 0.152939
R21522 gnd.n3332 gnd.n3331 0.152939
R21523 gnd.n3332 gnd.n2705 0.152939
R21524 gnd.n3343 gnd.n2705 0.152939
R21525 gnd.n3344 gnd.n3343 0.152939
R21526 gnd.n3345 gnd.n3344 0.152939
R21527 gnd.n3345 gnd.n2699 0.152939
R21528 gnd.n3359 gnd.n2699 0.152939
R21529 gnd.n3360 gnd.n3359 0.152939
R21530 gnd.n3361 gnd.n3360 0.152939
R21531 gnd.n3361 gnd.n2693 0.152939
R21532 gnd.n3375 gnd.n2693 0.152939
R21533 gnd.n3376 gnd.n3375 0.152939
R21534 gnd.n3377 gnd.n3376 0.152939
R21535 gnd.n3377 gnd.n2687 0.152939
R21536 gnd.n3391 gnd.n2687 0.152939
R21537 gnd.n3392 gnd.n3391 0.152939
R21538 gnd.n3393 gnd.n3392 0.152939
R21539 gnd.n3393 gnd.n2384 0.152939
R21540 gnd.n3567 gnd.n2384 0.152939
R21541 gnd.n3568 gnd.n3567 0.152939
R21542 gnd.n3569 gnd.n3568 0.152939
R21543 gnd.n3569 gnd.n2362 0.152939
R21544 gnd.n3595 gnd.n2362 0.152939
R21545 gnd.n3596 gnd.n3595 0.152939
R21546 gnd.n3597 gnd.n3596 0.152939
R21547 gnd.n3598 gnd.n3597 0.152939
R21548 gnd.n3598 gnd.n2334 0.152939
R21549 gnd.n3669 gnd.n2334 0.152939
R21550 gnd.n3670 gnd.n3669 0.152939
R21551 gnd.n3671 gnd.n3670 0.152939
R21552 gnd.n3671 gnd.n2314 0.152939
R21553 gnd.n3694 gnd.n2314 0.152939
R21554 gnd.n3695 gnd.n3694 0.152939
R21555 gnd.n3696 gnd.n3695 0.152939
R21556 gnd.n3696 gnd.n2294 0.152939
R21557 gnd.n3728 gnd.n2294 0.152939
R21558 gnd.n3729 gnd.n3728 0.152939
R21559 gnd.n3730 gnd.n3729 0.152939
R21560 gnd.n3730 gnd.n2277 0.152939
R21561 gnd.n3773 gnd.n2277 0.152939
R21562 gnd.n3774 gnd.n3773 0.152939
R21563 gnd.n3775 gnd.n3774 0.152939
R21564 gnd.n3776 gnd.n3775 0.152939
R21565 gnd.n3776 gnd.n2249 0.152939
R21566 gnd.n3846 gnd.n2249 0.152939
R21567 gnd.n3847 gnd.n3846 0.152939
R21568 gnd.n3848 gnd.n3847 0.152939
R21569 gnd.n3848 gnd.n2229 0.152939
R21570 gnd.n3872 gnd.n2229 0.152939
R21571 gnd.n3873 gnd.n3872 0.152939
R21572 gnd.n3874 gnd.n3873 0.152939
R21573 gnd.n3874 gnd.n2206 0.152939
R21574 gnd.n3905 gnd.n2206 0.152939
R21575 gnd.n3906 gnd.n3905 0.152939
R21576 gnd.n3907 gnd.n3906 0.152939
R21577 gnd.n3907 gnd.n2189 0.152939
R21578 gnd.n3951 gnd.n2189 0.152939
R21579 gnd.n3952 gnd.n3951 0.152939
R21580 gnd.n3953 gnd.n3952 0.152939
R21581 gnd.n3954 gnd.n3953 0.152939
R21582 gnd.n3954 gnd.n2162 0.152939
R21583 gnd.n4008 gnd.n2162 0.152939
R21584 gnd.n4009 gnd.n4008 0.152939
R21585 gnd.n4010 gnd.n4009 0.152939
R21586 gnd.n4010 gnd.n2141 0.152939
R21587 gnd.n4033 gnd.n2141 0.152939
R21588 gnd.n4034 gnd.n4033 0.152939
R21589 gnd.n4035 gnd.n4034 0.152939
R21590 gnd.n4035 gnd.n2119 0.152939
R21591 gnd.n4093 gnd.n2119 0.152939
R21592 gnd.n4094 gnd.n4093 0.152939
R21593 gnd.n4095 gnd.n4094 0.152939
R21594 gnd.n4095 gnd.n2097 0.152939
R21595 gnd.n4122 gnd.n2097 0.152939
R21596 gnd.n4123 gnd.n4122 0.152939
R21597 gnd.n4124 gnd.n4123 0.152939
R21598 gnd.n4125 gnd.n4124 0.152939
R21599 gnd.n4125 gnd.n2069 0.152939
R21600 gnd.n4172 gnd.n2069 0.152939
R21601 gnd.n4173 gnd.n4172 0.152939
R21602 gnd.n4174 gnd.n4173 0.152939
R21603 gnd.n4174 gnd.n2048 0.152939
R21604 gnd.n4198 gnd.n2048 0.152939
R21605 gnd.n4199 gnd.n4198 0.152939
R21606 gnd.n4200 gnd.n4199 0.152939
R21607 gnd.n4201 gnd.n4200 0.152939
R21608 gnd.n4201 gnd.n1844 0.152939
R21609 gnd.n4383 gnd.n1844 0.152939
R21610 gnd.n4384 gnd.n4383 0.152939
R21611 gnd.n4385 gnd.n4384 0.152939
R21612 gnd.n4385 gnd.n1831 0.152939
R21613 gnd.n4403 gnd.n1831 0.152939
R21614 gnd.n4404 gnd.n4403 0.152939
R21615 gnd.n4405 gnd.n4404 0.152939
R21616 gnd.n4405 gnd.n1818 0.152939
R21617 gnd.n4423 gnd.n1818 0.152939
R21618 gnd.n4424 gnd.n4423 0.152939
R21619 gnd.n4425 gnd.n4424 0.152939
R21620 gnd.n4425 gnd.n1805 0.152939
R21621 gnd.n4446 gnd.n1805 0.152939
R21622 gnd.n4447 gnd.n4446 0.152939
R21623 gnd.n4449 gnd.n4447 0.152939
R21624 gnd.n4449 gnd.n4448 0.152939
R21625 gnd.n4448 gnd.n1462 0.152939
R21626 gnd.n1463 gnd.n1462 0.152939
R21627 gnd.n1464 gnd.n1463 0.152939
R21628 gnd.n1470 gnd.n1464 0.152939
R21629 gnd.n1471 gnd.n1470 0.152939
R21630 gnd.n1472 gnd.n1471 0.152939
R21631 gnd.n1473 gnd.n1472 0.152939
R21632 gnd.n1626 gnd.n1473 0.152939
R21633 gnd.n1629 gnd.n1626 0.152939
R21634 gnd.n1630 gnd.n1629 0.152939
R21635 gnd.n1631 gnd.n1630 0.152939
R21636 gnd.n1631 gnd.n1613 0.152939
R21637 gnd.n4541 gnd.n1613 0.152939
R21638 gnd.n4542 gnd.n4541 0.152939
R21639 gnd.n4543 gnd.n4542 0.152939
R21640 gnd.n4544 gnd.n4543 0.152939
R21641 gnd.n4544 gnd.n1586 0.152939
R21642 gnd.n4574 gnd.n1586 0.152939
R21643 gnd.n4575 gnd.n4574 0.152939
R21644 gnd.n4576 gnd.n4575 0.152939
R21645 gnd.n4577 gnd.n4576 0.152939
R21646 gnd.n4578 gnd.n4577 0.152939
R21647 gnd.n4580 gnd.n4578 0.152939
R21648 gnd.n4580 gnd.n4579 0.152939
R21649 gnd.n4579 gnd.n1533 0.152939
R21650 gnd.n1534 gnd.n1533 0.152939
R21651 gnd.n1535 gnd.n1534 0.152939
R21652 gnd.n1536 gnd.n1535 0.152939
R21653 gnd.n1213 gnd.n1212 0.152939
R21654 gnd.n1230 gnd.n1213 0.152939
R21655 gnd.n1231 gnd.n1230 0.152939
R21656 gnd.n1232 gnd.n1231 0.152939
R21657 gnd.n1233 gnd.n1232 0.152939
R21658 gnd.n1252 gnd.n1233 0.152939
R21659 gnd.n1253 gnd.n1252 0.152939
R21660 gnd.n1254 gnd.n1253 0.152939
R21661 gnd.n1255 gnd.n1254 0.152939
R21662 gnd.n1272 gnd.n1255 0.152939
R21663 gnd.n1273 gnd.n1272 0.152939
R21664 gnd.n1274 gnd.n1273 0.152939
R21665 gnd.n1275 gnd.n1274 0.152939
R21666 gnd.n1294 gnd.n1275 0.152939
R21667 gnd.n1295 gnd.n1294 0.152939
R21668 gnd.n1296 gnd.n1295 0.152939
R21669 gnd.n1297 gnd.n1296 0.152939
R21670 gnd.n1315 gnd.n1297 0.152939
R21671 gnd.n1316 gnd.n1315 0.152939
R21672 gnd.n1317 gnd.n1316 0.152939
R21673 gnd.n1318 gnd.n1317 0.152939
R21674 gnd.n2565 gnd.n2564 0.152939
R21675 gnd.n2566 gnd.n2565 0.152939
R21676 gnd.n2567 gnd.n2566 0.152939
R21677 gnd.n2568 gnd.n2567 0.152939
R21678 gnd.n2569 gnd.n2568 0.152939
R21679 gnd.n2570 gnd.n2569 0.152939
R21680 gnd.n2571 gnd.n2570 0.152939
R21681 gnd.n2572 gnd.n2571 0.152939
R21682 gnd.n2573 gnd.n2572 0.152939
R21683 gnd.n2574 gnd.n2573 0.152939
R21684 gnd.n2575 gnd.n2574 0.152939
R21685 gnd.n2576 gnd.n2575 0.152939
R21686 gnd.n2577 gnd.n2576 0.152939
R21687 gnd.n2578 gnd.n2577 0.152939
R21688 gnd.n2578 gnd.n2548 0.152939
R21689 gnd.n3493 gnd.n3492 0.152939
R21690 gnd.n3492 gnd.n2549 0.152939
R21691 gnd.n2609 gnd.n2549 0.152939
R21692 gnd.n2610 gnd.n2609 0.152939
R21693 gnd.n2611 gnd.n2610 0.152939
R21694 gnd.n2612 gnd.n2611 0.152939
R21695 gnd.n2616 gnd.n2612 0.152939
R21696 gnd.n2617 gnd.n2616 0.152939
R21697 gnd.n2618 gnd.n2617 0.152939
R21698 gnd.n2619 gnd.n2618 0.152939
R21699 gnd.n2623 gnd.n2619 0.152939
R21700 gnd.n2624 gnd.n2623 0.152939
R21701 gnd.n2625 gnd.n2624 0.152939
R21702 gnd.n2626 gnd.n2625 0.152939
R21703 gnd.n2630 gnd.n2626 0.152939
R21704 gnd.n2631 gnd.n2630 0.152939
R21705 gnd.n2632 gnd.n2631 0.152939
R21706 gnd.n2633 gnd.n2632 0.152939
R21707 gnd.n2638 gnd.n2633 0.152939
R21708 gnd.n3455 gnd.n2638 0.152939
R21709 gnd.n3046 gnd.n3044 0.152939
R21710 gnd.n3044 gnd.n3019 0.152939
R21711 gnd.n3019 gnd.n3017 0.152939
R21712 gnd.n3107 gnd.n3017 0.152939
R21713 gnd.n3108 gnd.n3107 0.152939
R21714 gnd.n3109 gnd.n3108 0.152939
R21715 gnd.n3109 gnd.n3015 0.152939
R21716 gnd.n3115 gnd.n3015 0.152939
R21717 gnd.n3116 gnd.n3115 0.152939
R21718 gnd.n3117 gnd.n3116 0.152939
R21719 gnd.n3117 gnd.n3013 0.152939
R21720 gnd.n3144 gnd.n3013 0.152939
R21721 gnd.n3145 gnd.n3144 0.152939
R21722 gnd.n3146 gnd.n3145 0.152939
R21723 gnd.n3146 gnd.n3007 0.152939
R21724 gnd.n3160 gnd.n3007 0.152939
R21725 gnd.n3161 gnd.n3160 0.152939
R21726 gnd.n3162 gnd.n3161 0.152939
R21727 gnd.n3162 gnd.n2909 0.152939
R21728 gnd.n3176 gnd.n2909 0.152939
R21729 gnd.n3177 gnd.n3176 0.152939
R21730 gnd.n3178 gnd.n3177 0.152939
R21731 gnd.n3178 gnd.n2903 0.152939
R21732 gnd.n3192 gnd.n2903 0.152939
R21733 gnd.n3193 gnd.n3192 0.152939
R21734 gnd.n3195 gnd.n3193 0.152939
R21735 gnd.n3085 gnd.n3025 0.152939
R21736 gnd.n3026 gnd.n3025 0.152939
R21737 gnd.n3027 gnd.n3026 0.152939
R21738 gnd.n3028 gnd.n3027 0.152939
R21739 gnd.n3029 gnd.n3028 0.152939
R21740 gnd.n3030 gnd.n3029 0.152939
R21741 gnd.n3031 gnd.n3030 0.152939
R21742 gnd.n3032 gnd.n3031 0.152939
R21743 gnd.n3033 gnd.n3032 0.152939
R21744 gnd.n3034 gnd.n3033 0.152939
R21745 gnd.n3035 gnd.n3034 0.152939
R21746 gnd.n3036 gnd.n3035 0.152939
R21747 gnd.n3037 gnd.n3036 0.152939
R21748 gnd.n3038 gnd.n3037 0.152939
R21749 gnd.n3039 gnd.n3038 0.152939
R21750 gnd.n3050 gnd.n3039 0.152939
R21751 gnd.n3050 gnd.n3049 0.152939
R21752 gnd.n3049 gnd.n3048 0.152939
R21753 gnd.n3091 gnd.n3086 0.152939
R21754 gnd.n3091 gnd.n3090 0.152939
R21755 gnd.n3090 gnd.n3089 0.152939
R21756 gnd.n3089 gnd.n3087 0.152939
R21757 gnd.n3087 gnd.n1081 0.152939
R21758 gnd.n1082 gnd.n1081 0.152939
R21759 gnd.n1083 gnd.n1082 0.152939
R21760 gnd.n1099 gnd.n1083 0.152939
R21761 gnd.n1100 gnd.n1099 0.152939
R21762 gnd.n1101 gnd.n1100 0.152939
R21763 gnd.n1102 gnd.n1101 0.152939
R21764 gnd.n1121 gnd.n1102 0.152939
R21765 gnd.n1122 gnd.n1121 0.152939
R21766 gnd.n1123 gnd.n1122 0.152939
R21767 gnd.n1124 gnd.n1123 0.152939
R21768 gnd.n1142 gnd.n1124 0.152939
R21769 gnd.n1143 gnd.n1142 0.152939
R21770 gnd.n1144 gnd.n1143 0.152939
R21771 gnd.n1145 gnd.n1144 0.152939
R21772 gnd.n1163 gnd.n1145 0.152939
R21773 gnd.n1164 gnd.n1163 0.152939
R21774 gnd.n1165 gnd.n1164 0.152939
R21775 gnd.n1166 gnd.n1165 0.152939
R21776 gnd.n1182 gnd.n1166 0.152939
R21777 gnd.n1183 gnd.n1182 0.152939
R21778 gnd.n1184 gnd.n1183 0.152939
R21779 gnd.n1200 gnd.n1185 0.152939
R21780 gnd.n1201 gnd.n1200 0.152939
R21781 gnd.n1202 gnd.n1201 0.152939
R21782 gnd.n1203 gnd.n1202 0.152939
R21783 gnd.n1220 gnd.n1203 0.152939
R21784 gnd.n1221 gnd.n1220 0.152939
R21785 gnd.n1222 gnd.n1221 0.152939
R21786 gnd.n1223 gnd.n1222 0.152939
R21787 gnd.n1241 gnd.n1223 0.152939
R21788 gnd.n1242 gnd.n1241 0.152939
R21789 gnd.n1243 gnd.n1242 0.152939
R21790 gnd.n1244 gnd.n1243 0.152939
R21791 gnd.n1262 gnd.n1244 0.152939
R21792 gnd.n1263 gnd.n1262 0.152939
R21793 gnd.n1264 gnd.n1263 0.152939
R21794 gnd.n1265 gnd.n1264 0.152939
R21795 gnd.n1283 gnd.n1265 0.152939
R21796 gnd.n1284 gnd.n1283 0.152939
R21797 gnd.n1285 gnd.n1284 0.152939
R21798 gnd.n1286 gnd.n1285 0.152939
R21799 gnd.n1305 gnd.n1286 0.152939
R21800 gnd.n1306 gnd.n1305 0.152939
R21801 gnd.n1307 gnd.n1306 0.152939
R21802 gnd.n1308 gnd.n1307 0.152939
R21803 gnd.n1325 gnd.n1308 0.152939
R21804 gnd.n4897 gnd.n1325 0.152939
R21805 gnd.n5056 gnd.n1056 0.152939
R21806 gnd.n5056 gnd.n5055 0.152939
R21807 gnd.n5055 gnd.n5054 0.152939
R21808 gnd.n5054 gnd.n1059 0.152939
R21809 gnd.n3124 gnd.n1059 0.152939
R21810 gnd.n3128 gnd.n3124 0.152939
R21811 gnd.n3129 gnd.n3128 0.152939
R21812 gnd.n3130 gnd.n3129 0.152939
R21813 gnd.n3130 gnd.n3122 0.152939
R21814 gnd.n3136 gnd.n3122 0.152939
R21815 gnd.n3137 gnd.n3136 0.152939
R21816 gnd.n3138 gnd.n3137 0.152939
R21817 gnd.n3138 gnd.n3010 0.152939
R21818 gnd.n3152 gnd.n3010 0.152939
R21819 gnd.n3153 gnd.n3152 0.152939
R21820 gnd.n3154 gnd.n3153 0.152939
R21821 gnd.n3154 gnd.n2913 0.152939
R21822 gnd.n3168 gnd.n2913 0.152939
R21823 gnd.n3169 gnd.n3168 0.152939
R21824 gnd.n3170 gnd.n3169 0.152939
R21825 gnd.n3170 gnd.n2906 0.152939
R21826 gnd.n3184 gnd.n2906 0.152939
R21827 gnd.n3185 gnd.n3184 0.152939
R21828 gnd.n3186 gnd.n3185 0.152939
R21829 gnd.n3186 gnd.n2899 0.152939
R21830 gnd.n3201 gnd.n2899 0.152939
R21831 gnd.n3204 gnd.n3203 0.152939
R21832 gnd.n3204 gnd.n2891 0.152939
R21833 gnd.n3218 gnd.n2891 0.152939
R21834 gnd.n3219 gnd.n3218 0.152939
R21835 gnd.n3220 gnd.n3219 0.152939
R21836 gnd.n3220 gnd.n2884 0.152939
R21837 gnd.n3234 gnd.n2884 0.152939
R21838 gnd.n3235 gnd.n3234 0.152939
R21839 gnd.n3236 gnd.n3235 0.152939
R21840 gnd.n3236 gnd.n2877 0.152939
R21841 gnd.n3250 gnd.n2877 0.152939
R21842 gnd.n3251 gnd.n3250 0.152939
R21843 gnd.n3253 gnd.n3251 0.152939
R21844 gnd.n3253 gnd.n3252 0.152939
R21845 gnd.n3252 gnd.n2871 0.152939
R21846 gnd.n2871 gnd.n2869 0.152939
R21847 gnd.n3269 gnd.n2869 0.152939
R21848 gnd.n3270 gnd.n3269 0.152939
R21849 gnd.n3271 gnd.n3270 0.152939
R21850 gnd.n3271 gnd.n2867 0.152939
R21851 gnd.n3279 gnd.n2867 0.152939
R21852 gnd.n3280 gnd.n3279 0.152939
R21853 gnd.n3282 gnd.n3280 0.152939
R21854 gnd.n3282 gnd.n3281 0.152939
R21855 gnd.n3281 gnd.n2639 0.152939
R21856 gnd.n3454 gnd.n2639 0.152939
R21857 gnd.n1014 gnd.n1013 0.152939
R21858 gnd.n1015 gnd.n1014 0.152939
R21859 gnd.n1016 gnd.n1015 0.152939
R21860 gnd.n1017 gnd.n1016 0.152939
R21861 gnd.n1018 gnd.n1017 0.152939
R21862 gnd.n1019 gnd.n1018 0.152939
R21863 gnd.n1020 gnd.n1019 0.152939
R21864 gnd.n1021 gnd.n1020 0.152939
R21865 gnd.n1022 gnd.n1021 0.152939
R21866 gnd.n1023 gnd.n1022 0.152939
R21867 gnd.n1024 gnd.n1023 0.152939
R21868 gnd.n1025 gnd.n1024 0.152939
R21869 gnd.n1026 gnd.n1025 0.152939
R21870 gnd.n1027 gnd.n1026 0.152939
R21871 gnd.n1028 gnd.n1027 0.152939
R21872 gnd.n1029 gnd.n1028 0.152939
R21873 gnd.n1030 gnd.n1029 0.152939
R21874 gnd.n1033 gnd.n1030 0.152939
R21875 gnd.n1034 gnd.n1033 0.152939
R21876 gnd.n1035 gnd.n1034 0.152939
R21877 gnd.n1036 gnd.n1035 0.152939
R21878 gnd.n1037 gnd.n1036 0.152939
R21879 gnd.n1038 gnd.n1037 0.152939
R21880 gnd.n1039 gnd.n1038 0.152939
R21881 gnd.n1040 gnd.n1039 0.152939
R21882 gnd.n1041 gnd.n1040 0.152939
R21883 gnd.n1042 gnd.n1041 0.152939
R21884 gnd.n1043 gnd.n1042 0.152939
R21885 gnd.n1044 gnd.n1043 0.152939
R21886 gnd.n1045 gnd.n1044 0.152939
R21887 gnd.n1046 gnd.n1045 0.152939
R21888 gnd.n1047 gnd.n1046 0.152939
R21889 gnd.n1048 gnd.n1047 0.152939
R21890 gnd.n1049 gnd.n1048 0.152939
R21891 gnd.n1050 gnd.n1049 0.152939
R21892 gnd.n5064 gnd.n1050 0.152939
R21893 gnd.n5064 gnd.n5063 0.152939
R21894 gnd.n5063 gnd.n5062 0.152939
R21895 gnd.n3097 gnd.n3095 0.152939
R21896 gnd.n3097 gnd.n3096 0.152939
R21897 gnd.n3096 gnd.n1070 0.152939
R21898 gnd.n1071 gnd.n1070 0.152939
R21899 gnd.n1072 gnd.n1071 0.152939
R21900 gnd.n1090 gnd.n1072 0.152939
R21901 gnd.n1091 gnd.n1090 0.152939
R21902 gnd.n1092 gnd.n1091 0.152939
R21903 gnd.n1093 gnd.n1092 0.152939
R21904 gnd.n1110 gnd.n1093 0.152939
R21905 gnd.n1111 gnd.n1110 0.152939
R21906 gnd.n1112 gnd.n1111 0.152939
R21907 gnd.n1113 gnd.n1112 0.152939
R21908 gnd.n1132 gnd.n1113 0.152939
R21909 gnd.n1133 gnd.n1132 0.152939
R21910 gnd.n1134 gnd.n1133 0.152939
R21911 gnd.n1135 gnd.n1134 0.152939
R21912 gnd.n1152 gnd.n1135 0.152939
R21913 gnd.n1153 gnd.n1152 0.152939
R21914 gnd.n1154 gnd.n1153 0.152939
R21915 gnd.n1155 gnd.n1154 0.152939
R21916 gnd.n2927 gnd.n2926 0.152939
R21917 gnd.n2927 gnd.n2918 0.152939
R21918 gnd.n2933 gnd.n2918 0.152939
R21919 gnd.n2934 gnd.n2933 0.152939
R21920 gnd.n2935 gnd.n2934 0.152939
R21921 gnd.n2936 gnd.n2935 0.152939
R21922 gnd.n2937 gnd.n2936 0.152939
R21923 gnd.n2994 gnd.n2937 0.152939
R21924 gnd.n743 gnd.n742 0.152939
R21925 gnd.n744 gnd.n743 0.152939
R21926 gnd.n749 gnd.n744 0.152939
R21927 gnd.n750 gnd.n749 0.152939
R21928 gnd.n751 gnd.n750 0.152939
R21929 gnd.n752 gnd.n751 0.152939
R21930 gnd.n757 gnd.n752 0.152939
R21931 gnd.n758 gnd.n757 0.152939
R21932 gnd.n759 gnd.n758 0.152939
R21933 gnd.n760 gnd.n759 0.152939
R21934 gnd.n765 gnd.n760 0.152939
R21935 gnd.n766 gnd.n765 0.152939
R21936 gnd.n767 gnd.n766 0.152939
R21937 gnd.n768 gnd.n767 0.152939
R21938 gnd.n773 gnd.n768 0.152939
R21939 gnd.n774 gnd.n773 0.152939
R21940 gnd.n775 gnd.n774 0.152939
R21941 gnd.n776 gnd.n775 0.152939
R21942 gnd.n781 gnd.n776 0.152939
R21943 gnd.n782 gnd.n781 0.152939
R21944 gnd.n783 gnd.n782 0.152939
R21945 gnd.n784 gnd.n783 0.152939
R21946 gnd.n789 gnd.n784 0.152939
R21947 gnd.n790 gnd.n789 0.152939
R21948 gnd.n791 gnd.n790 0.152939
R21949 gnd.n792 gnd.n791 0.152939
R21950 gnd.n797 gnd.n792 0.152939
R21951 gnd.n798 gnd.n797 0.152939
R21952 gnd.n799 gnd.n798 0.152939
R21953 gnd.n800 gnd.n799 0.152939
R21954 gnd.n805 gnd.n800 0.152939
R21955 gnd.n806 gnd.n805 0.152939
R21956 gnd.n807 gnd.n806 0.152939
R21957 gnd.n808 gnd.n807 0.152939
R21958 gnd.n813 gnd.n808 0.152939
R21959 gnd.n814 gnd.n813 0.152939
R21960 gnd.n815 gnd.n814 0.152939
R21961 gnd.n816 gnd.n815 0.152939
R21962 gnd.n821 gnd.n816 0.152939
R21963 gnd.n822 gnd.n821 0.152939
R21964 gnd.n823 gnd.n822 0.152939
R21965 gnd.n824 gnd.n823 0.152939
R21966 gnd.n829 gnd.n824 0.152939
R21967 gnd.n830 gnd.n829 0.152939
R21968 gnd.n831 gnd.n830 0.152939
R21969 gnd.n832 gnd.n831 0.152939
R21970 gnd.n837 gnd.n832 0.152939
R21971 gnd.n838 gnd.n837 0.152939
R21972 gnd.n839 gnd.n838 0.152939
R21973 gnd.n840 gnd.n839 0.152939
R21974 gnd.n845 gnd.n840 0.152939
R21975 gnd.n846 gnd.n845 0.152939
R21976 gnd.n847 gnd.n846 0.152939
R21977 gnd.n848 gnd.n847 0.152939
R21978 gnd.n853 gnd.n848 0.152939
R21979 gnd.n854 gnd.n853 0.152939
R21980 gnd.n855 gnd.n854 0.152939
R21981 gnd.n856 gnd.n855 0.152939
R21982 gnd.n861 gnd.n856 0.152939
R21983 gnd.n862 gnd.n861 0.152939
R21984 gnd.n863 gnd.n862 0.152939
R21985 gnd.n864 gnd.n863 0.152939
R21986 gnd.n869 gnd.n864 0.152939
R21987 gnd.n870 gnd.n869 0.152939
R21988 gnd.n871 gnd.n870 0.152939
R21989 gnd.n872 gnd.n871 0.152939
R21990 gnd.n877 gnd.n872 0.152939
R21991 gnd.n878 gnd.n877 0.152939
R21992 gnd.n879 gnd.n878 0.152939
R21993 gnd.n880 gnd.n879 0.152939
R21994 gnd.n885 gnd.n880 0.152939
R21995 gnd.n886 gnd.n885 0.152939
R21996 gnd.n887 gnd.n886 0.152939
R21997 gnd.n888 gnd.n887 0.152939
R21998 gnd.n893 gnd.n888 0.152939
R21999 gnd.n894 gnd.n893 0.152939
R22000 gnd.n895 gnd.n894 0.152939
R22001 gnd.n896 gnd.n895 0.152939
R22002 gnd.n901 gnd.n896 0.152939
R22003 gnd.n902 gnd.n901 0.152939
R22004 gnd.n903 gnd.n902 0.152939
R22005 gnd.n904 gnd.n903 0.152939
R22006 gnd.n2922 gnd.n904 0.152939
R22007 gnd.n2925 gnd.n2922 0.152939
R22008 gnd.n4471 gnd.n4470 0.152939
R22009 gnd.n4470 gnd.n4469 0.152939
R22010 gnd.n4469 gnd.n1780 0.152939
R22011 gnd.n4465 gnd.n1780 0.152939
R22012 gnd.n4465 gnd.n4464 0.152939
R22013 gnd.n4464 gnd.n4463 0.152939
R22014 gnd.n4463 gnd.n1788 0.152939
R22015 gnd.n4459 gnd.n1788 0.152939
R22016 gnd.n4459 gnd.n4458 0.152939
R22017 gnd.n3427 gnd.n2664 0.152939
R22018 gnd.n3423 gnd.n2664 0.152939
R22019 gnd.n3423 gnd.n3422 0.152939
R22020 gnd.n3422 gnd.n3421 0.152939
R22021 gnd.n3421 gnd.n2669 0.152939
R22022 gnd.n3417 gnd.n2669 0.152939
R22023 gnd.n3417 gnd.n3416 0.152939
R22024 gnd.n3416 gnd.n3415 0.152939
R22025 gnd.n3415 gnd.n2674 0.152939
R22026 gnd.n3411 gnd.n2674 0.152939
R22027 gnd.n3411 gnd.n3410 0.152939
R22028 gnd.n3410 gnd.n3409 0.152939
R22029 gnd.n3409 gnd.n2679 0.152939
R22030 gnd.n3405 gnd.n2679 0.152939
R22031 gnd.n3405 gnd.n3404 0.152939
R22032 gnd.n3404 gnd.n3403 0.152939
R22033 gnd.n3403 gnd.n2377 0.152939
R22034 gnd.n3576 gnd.n2377 0.152939
R22035 gnd.n3577 gnd.n3576 0.152939
R22036 gnd.n3579 gnd.n3577 0.152939
R22037 gnd.n3579 gnd.n3578 0.152939
R22038 gnd.n3578 gnd.n2348 0.152939
R22039 gnd.n3615 gnd.n2348 0.152939
R22040 gnd.n3616 gnd.n3615 0.152939
R22041 gnd.n3654 gnd.n3616 0.152939
R22042 gnd.n3654 gnd.n3653 0.152939
R22043 gnd.n3653 gnd.n3652 0.152939
R22044 gnd.n3652 gnd.n3617 0.152939
R22045 gnd.n3648 gnd.n3617 0.152939
R22046 gnd.n3648 gnd.n3647 0.152939
R22047 gnd.n3647 gnd.n3646 0.152939
R22048 gnd.n3646 gnd.n3622 0.152939
R22049 gnd.n3642 gnd.n3622 0.152939
R22050 gnd.n3642 gnd.n3641 0.152939
R22051 gnd.n3641 gnd.n3640 0.152939
R22052 gnd.n3640 gnd.n3628 0.152939
R22053 gnd.n3636 gnd.n3628 0.152939
R22054 gnd.n3636 gnd.n3635 0.152939
R22055 gnd.n3635 gnd.n2263 0.152939
R22056 gnd.n3793 gnd.n2263 0.152939
R22057 gnd.n3794 gnd.n3793 0.152939
R22058 gnd.n3830 gnd.n3794 0.152939
R22059 gnd.n3830 gnd.n3829 0.152939
R22060 gnd.n3829 gnd.n3828 0.152939
R22061 gnd.n3828 gnd.n3795 0.152939
R22062 gnd.n3824 gnd.n3795 0.152939
R22063 gnd.n3824 gnd.n3823 0.152939
R22064 gnd.n3823 gnd.n3822 0.152939
R22065 gnd.n3822 gnd.n3800 0.152939
R22066 gnd.n3818 gnd.n3800 0.152939
R22067 gnd.n3818 gnd.n3817 0.152939
R22068 gnd.n3817 gnd.n3816 0.152939
R22069 gnd.n3816 gnd.n3804 0.152939
R22070 gnd.n3812 gnd.n3804 0.152939
R22071 gnd.n3812 gnd.n3811 0.152939
R22072 gnd.n3811 gnd.n2176 0.152939
R22073 gnd.n3970 gnd.n2176 0.152939
R22074 gnd.n3971 gnd.n3970 0.152939
R22075 gnd.n3992 gnd.n3971 0.152939
R22076 gnd.n3992 gnd.n3991 0.152939
R22077 gnd.n3991 gnd.n3990 0.152939
R22078 gnd.n3990 gnd.n3972 0.152939
R22079 gnd.n3986 gnd.n3972 0.152939
R22080 gnd.n3986 gnd.n3985 0.152939
R22081 gnd.n3985 gnd.n3984 0.152939
R22082 gnd.n3984 gnd.n3977 0.152939
R22083 gnd.n3980 gnd.n3977 0.152939
R22084 gnd.n3980 gnd.n2111 0.152939
R22085 gnd.n4102 gnd.n2111 0.152939
R22086 gnd.n4103 gnd.n4102 0.152939
R22087 gnd.n4105 gnd.n4103 0.152939
R22088 gnd.n4105 gnd.n4104 0.152939
R22089 gnd.n4104 gnd.n2084 0.152939
R22090 gnd.n4141 gnd.n2084 0.152939
R22091 gnd.n4142 gnd.n4141 0.152939
R22092 gnd.n4157 gnd.n4142 0.152939
R22093 gnd.n4157 gnd.n4156 0.152939
R22094 gnd.n4156 gnd.n4155 0.152939
R22095 gnd.n4155 gnd.n4143 0.152939
R22096 gnd.n4151 gnd.n4143 0.152939
R22097 gnd.n4151 gnd.n4150 0.152939
R22098 gnd.n4150 gnd.n4149 0.152939
R22099 gnd.n4149 gnd.n1849 0.152939
R22100 gnd.n4373 gnd.n1849 0.152939
R22101 gnd.n4374 gnd.n4373 0.152939
R22102 gnd.n4375 gnd.n4374 0.152939
R22103 gnd.n4375 gnd.n1837 0.152939
R22104 gnd.n4393 gnd.n1837 0.152939
R22105 gnd.n4394 gnd.n4393 0.152939
R22106 gnd.n4395 gnd.n4394 0.152939
R22107 gnd.n4395 gnd.n1824 0.152939
R22108 gnd.n4413 gnd.n1824 0.152939
R22109 gnd.n4414 gnd.n4413 0.152939
R22110 gnd.n4415 gnd.n4414 0.152939
R22111 gnd.n4415 gnd.n1811 0.152939
R22112 gnd.n4433 gnd.n1811 0.152939
R22113 gnd.n4434 gnd.n4433 0.152939
R22114 gnd.n4436 gnd.n4434 0.152939
R22115 gnd.n4436 gnd.n4435 0.152939
R22116 gnd.n4435 gnd.n1800 0.152939
R22117 gnd.n4457 gnd.n1800 0.152939
R22118 gnd.n3440 gnd.n2645 0.152939
R22119 gnd.n3440 gnd.n3439 0.152939
R22120 gnd.n3439 gnd.n3438 0.152939
R22121 gnd.n3438 gnd.n2652 0.152939
R22122 gnd.n3434 gnd.n2652 0.152939
R22123 gnd.n3434 gnd.n3433 0.152939
R22124 gnd.n3433 gnd.n2659 0.152939
R22125 gnd.n3429 gnd.n2659 0.152939
R22126 gnd.n3429 gnd.n3428 0.152939
R22127 gnd.n3210 gnd.n2894 0.152939
R22128 gnd.n3211 gnd.n3210 0.152939
R22129 gnd.n3212 gnd.n3211 0.152939
R22130 gnd.n3212 gnd.n2888 0.152939
R22131 gnd.n3226 gnd.n2888 0.152939
R22132 gnd.n3227 gnd.n3226 0.152939
R22133 gnd.n3228 gnd.n3227 0.152939
R22134 gnd.n3228 gnd.n2880 0.152939
R22135 gnd.n3242 gnd.n2880 0.152939
R22136 gnd.n3243 gnd.n3242 0.152939
R22137 gnd.n3244 gnd.n3243 0.152939
R22138 gnd.n3244 gnd.n2874 0.152939
R22139 gnd.n3259 gnd.n2874 0.152939
R22140 gnd.n3260 gnd.n3259 0.152939
R22141 gnd.n3261 gnd.n3260 0.152939
R22142 gnd.n3261 gnd.n2861 0.152939
R22143 gnd.n3296 gnd.n2861 0.152939
R22144 gnd.n3296 gnd.n3295 0.152939
R22145 gnd.n3295 gnd.n3294 0.152939
R22146 gnd.n3294 gnd.n2862 0.152939
R22147 gnd.n3290 gnd.n2862 0.152939
R22148 gnd.n3290 gnd.n3289 0.152939
R22149 gnd.n3289 gnd.n3288 0.152939
R22150 gnd.n3288 gnd.n2644 0.152939
R22151 gnd.n3447 gnd.n2644 0.152939
R22152 gnd.n3447 gnd.n3446 0.152939
R22153 gnd.n4894 gnd.n1328 0.152939
R22154 gnd.n4890 gnd.n1328 0.152939
R22155 gnd.n4890 gnd.n4889 0.152939
R22156 gnd.n4889 gnd.n4888 0.152939
R22157 gnd.n4888 gnd.n1333 0.152939
R22158 gnd.n4884 gnd.n1333 0.152939
R22159 gnd.n4884 gnd.n4883 0.152939
R22160 gnd.n4883 gnd.n4882 0.152939
R22161 gnd.n4882 gnd.n1338 0.152939
R22162 gnd.n4878 gnd.n1338 0.152939
R22163 gnd.n4878 gnd.n4877 0.152939
R22164 gnd.n4877 gnd.n4876 0.152939
R22165 gnd.n4876 gnd.n1343 0.152939
R22166 gnd.n4872 gnd.n1343 0.152939
R22167 gnd.n4872 gnd.n4871 0.152939
R22168 gnd.n4871 gnd.n4870 0.152939
R22169 gnd.n4870 gnd.n1348 0.152939
R22170 gnd.n4866 gnd.n1348 0.152939
R22171 gnd.n4866 gnd.n4865 0.152939
R22172 gnd.n4865 gnd.n4864 0.152939
R22173 gnd.n4864 gnd.n1353 0.152939
R22174 gnd.n4860 gnd.n1353 0.152939
R22175 gnd.n4860 gnd.n4859 0.152939
R22176 gnd.n4859 gnd.n4858 0.152939
R22177 gnd.n4858 gnd.n1358 0.152939
R22178 gnd.n4854 gnd.n1358 0.152939
R22179 gnd.n4854 gnd.n4853 0.152939
R22180 gnd.n4853 gnd.n4852 0.152939
R22181 gnd.n4852 gnd.n1363 0.152939
R22182 gnd.n4848 gnd.n1363 0.152939
R22183 gnd.n4848 gnd.n4847 0.152939
R22184 gnd.n4847 gnd.n4846 0.152939
R22185 gnd.n4846 gnd.n1368 0.152939
R22186 gnd.n4842 gnd.n1368 0.152939
R22187 gnd.n4842 gnd.n4841 0.152939
R22188 gnd.n4841 gnd.n4840 0.152939
R22189 gnd.n4840 gnd.n1373 0.152939
R22190 gnd.n4836 gnd.n1373 0.152939
R22191 gnd.n4836 gnd.n4835 0.152939
R22192 gnd.n4835 gnd.n4834 0.152939
R22193 gnd.n4834 gnd.n1378 0.152939
R22194 gnd.n4830 gnd.n1378 0.152939
R22195 gnd.n4830 gnd.n4829 0.152939
R22196 gnd.n4829 gnd.n4828 0.152939
R22197 gnd.n4828 gnd.n1383 0.152939
R22198 gnd.n4824 gnd.n1383 0.152939
R22199 gnd.n4824 gnd.n4823 0.152939
R22200 gnd.n4823 gnd.n4822 0.152939
R22201 gnd.n4822 gnd.n1388 0.152939
R22202 gnd.n4818 gnd.n1388 0.152939
R22203 gnd.n4818 gnd.n4817 0.152939
R22204 gnd.n4817 gnd.n4816 0.152939
R22205 gnd.n4816 gnd.n1393 0.152939
R22206 gnd.n4812 gnd.n1393 0.152939
R22207 gnd.n4812 gnd.n4811 0.152939
R22208 gnd.n4811 gnd.n4810 0.152939
R22209 gnd.n4810 gnd.n1398 0.152939
R22210 gnd.n4806 gnd.n1398 0.152939
R22211 gnd.n4806 gnd.n4805 0.152939
R22212 gnd.n4805 gnd.n4804 0.152939
R22213 gnd.n4804 gnd.n1403 0.152939
R22214 gnd.n4800 gnd.n1403 0.152939
R22215 gnd.n4800 gnd.n4799 0.152939
R22216 gnd.n4799 gnd.n4798 0.152939
R22217 gnd.n4798 gnd.n1408 0.152939
R22218 gnd.n4794 gnd.n1408 0.152939
R22219 gnd.n4794 gnd.n4793 0.152939
R22220 gnd.n4793 gnd.n4792 0.152939
R22221 gnd.n4792 gnd.n1413 0.152939
R22222 gnd.n4788 gnd.n1413 0.152939
R22223 gnd.n4788 gnd.n4787 0.152939
R22224 gnd.n4787 gnd.n4786 0.152939
R22225 gnd.n4786 gnd.n1418 0.152939
R22226 gnd.n4782 gnd.n1418 0.152939
R22227 gnd.n4782 gnd.n4781 0.152939
R22228 gnd.n4781 gnd.n4780 0.152939
R22229 gnd.n4780 gnd.n1423 0.152939
R22230 gnd.n4776 gnd.n1423 0.152939
R22231 gnd.n4776 gnd.n4775 0.152939
R22232 gnd.n4775 gnd.n4774 0.152939
R22233 gnd.n4774 gnd.n1428 0.152939
R22234 gnd.n4770 gnd.n1428 0.152939
R22235 gnd.n4770 gnd.n4769 0.152939
R22236 gnd.n4769 gnd.n4768 0.152939
R22237 gnd.n4768 gnd.n1433 0.152939
R22238 gnd.n4764 gnd.n1433 0.152939
R22239 gnd.n4764 gnd.n4763 0.152939
R22240 gnd.n4763 gnd.n4762 0.152939
R22241 gnd.n4762 gnd.n1438 0.152939
R22242 gnd.n4758 gnd.n1438 0.152939
R22243 gnd.n4758 gnd.n4757 0.152939
R22244 gnd.n4757 gnd.n4756 0.152939
R22245 gnd.n4756 gnd.n1443 0.152939
R22246 gnd.n4752 gnd.n1443 0.152939
R22247 gnd.n4752 gnd.n4751 0.152939
R22248 gnd.n4751 gnd.n4750 0.152939
R22249 gnd.n4750 gnd.n1448 0.152939
R22250 gnd.n4746 gnd.n1448 0.152939
R22251 gnd.n4746 gnd.n4745 0.152939
R22252 gnd.n4745 gnd.n4744 0.152939
R22253 gnd.n4744 gnd.n1453 0.152939
R22254 gnd.n1691 gnd.n1685 0.152939
R22255 gnd.n1685 gnd.n1498 0.152939
R22256 gnd.n4715 gnd.n1498 0.152939
R22257 gnd.n4715 gnd.n4714 0.152939
R22258 gnd.n4714 gnd.n4713 0.152939
R22259 gnd.n4713 gnd.n1499 0.152939
R22260 gnd.n4709 gnd.n1499 0.152939
R22261 gnd.n4709 gnd.n4708 0.152939
R22262 gnd.n4708 gnd.n4707 0.152939
R22263 gnd.n4707 gnd.n1504 0.152939
R22264 gnd.n4703 gnd.n1504 0.152939
R22265 gnd.n4703 gnd.n4702 0.152939
R22266 gnd.n4702 gnd.n4701 0.152939
R22267 gnd.n4701 gnd.n1509 0.152939
R22268 gnd.n4697 gnd.n1509 0.152939
R22269 gnd.n4697 gnd.n4696 0.152939
R22270 gnd.n4696 gnd.n4695 0.152939
R22271 gnd.n4695 gnd.n1514 0.152939
R22272 gnd.n4691 gnd.n1514 0.152939
R22273 gnd.n4691 gnd.n4690 0.152939
R22274 gnd.n4690 gnd.n285 0.152939
R22275 gnd.n7498 gnd.n285 0.152939
R22276 gnd.n7498 gnd.n7497 0.152939
R22277 gnd.n7497 gnd.n7496 0.152939
R22278 gnd.n7496 gnd.n286 0.152939
R22279 gnd.n7492 gnd.n286 0.152939
R22280 gnd.n7490 gnd.n7489 0.152939
R22281 gnd.n7489 gnd.n292 0.152939
R22282 gnd.n292 gnd.n260 0.152939
R22283 gnd.n7511 gnd.n260 0.152939
R22284 gnd.n7512 gnd.n7511 0.152939
R22285 gnd.n7513 gnd.n7512 0.152939
R22286 gnd.n7513 gnd.n244 0.152939
R22287 gnd.n7527 gnd.n244 0.152939
R22288 gnd.n7528 gnd.n7527 0.152939
R22289 gnd.n7529 gnd.n7528 0.152939
R22290 gnd.n7529 gnd.n229 0.152939
R22291 gnd.n7543 gnd.n229 0.152939
R22292 gnd.n7544 gnd.n7543 0.152939
R22293 gnd.n7545 gnd.n7544 0.152939
R22294 gnd.n7545 gnd.n214 0.152939
R22295 gnd.n7559 gnd.n214 0.152939
R22296 gnd.n7560 gnd.n7559 0.152939
R22297 gnd.n7561 gnd.n7560 0.152939
R22298 gnd.n7561 gnd.n199 0.152939
R22299 gnd.n7575 gnd.n199 0.152939
R22300 gnd.n7576 gnd.n7575 0.152939
R22301 gnd.n7652 gnd.n7576 0.152939
R22302 gnd.n7652 gnd.n7651 0.152939
R22303 gnd.n7651 gnd.n7650 0.152939
R22304 gnd.n7650 gnd.n7577 0.152939
R22305 gnd.n7646 gnd.n7577 0.152939
R22306 gnd.n7645 gnd.n7579 0.152939
R22307 gnd.n7641 gnd.n7579 0.152939
R22308 gnd.n7641 gnd.n7640 0.152939
R22309 gnd.n7640 gnd.n7639 0.152939
R22310 gnd.n7639 gnd.n7585 0.152939
R22311 gnd.n7635 gnd.n7585 0.152939
R22312 gnd.n7635 gnd.n7634 0.152939
R22313 gnd.n7634 gnd.n7633 0.152939
R22314 gnd.n7633 gnd.n7593 0.152939
R22315 gnd.n7629 gnd.n7593 0.152939
R22316 gnd.n7629 gnd.n7628 0.152939
R22317 gnd.n7628 gnd.n7627 0.152939
R22318 gnd.n7627 gnd.n7601 0.152939
R22319 gnd.n7623 gnd.n7601 0.152939
R22320 gnd.n7623 gnd.n7622 0.152939
R22321 gnd.n7622 gnd.n7621 0.152939
R22322 gnd.n7621 gnd.n7609 0.152939
R22323 gnd.n7617 gnd.n7609 0.152939
R22324 gnd.n4482 gnd.n4481 0.152939
R22325 gnd.n4484 gnd.n4482 0.152939
R22326 gnd.n4484 gnd.n4483 0.152939
R22327 gnd.n4483 gnd.n1621 0.152939
R22328 gnd.n4531 gnd.n1621 0.152939
R22329 gnd.n4532 gnd.n4531 0.152939
R22330 gnd.n4534 gnd.n4532 0.152939
R22331 gnd.n4534 gnd.n4533 0.152939
R22332 gnd.n4533 gnd.n1594 0.152939
R22333 gnd.n4563 gnd.n1594 0.152939
R22334 gnd.n4564 gnd.n4563 0.152939
R22335 gnd.n4566 gnd.n4564 0.152939
R22336 gnd.n4566 gnd.n4565 0.152939
R22337 gnd.n4565 gnd.n1565 0.152939
R22338 gnd.n4602 gnd.n1565 0.152939
R22339 gnd.n4603 gnd.n4602 0.152939
R22340 gnd.n4608 gnd.n4603 0.152939
R22341 gnd.n4608 gnd.n4607 0.152939
R22342 gnd.n4607 gnd.n4606 0.152939
R22343 gnd.n4606 gnd.n1554 0.152939
R22344 gnd.n4628 gnd.n1554 0.152939
R22345 gnd.n4629 gnd.n4628 0.152939
R22346 gnd.n4633 gnd.n4629 0.152939
R22347 gnd.n4633 gnd.n4632 0.152939
R22348 gnd.n4632 gnd.n4631 0.152939
R22349 gnd.n4631 gnd.n67 0.152939
R22350 gnd.n7784 gnd.n68 0.152939
R22351 gnd.n7780 gnd.n68 0.152939
R22352 gnd.n7780 gnd.n7779 0.152939
R22353 gnd.n7779 gnd.n7778 0.152939
R22354 gnd.n7778 gnd.n74 0.152939
R22355 gnd.n7774 gnd.n74 0.152939
R22356 gnd.n7774 gnd.n7773 0.152939
R22357 gnd.n7773 gnd.n7772 0.152939
R22358 gnd.n7772 gnd.n79 0.152939
R22359 gnd.n7768 gnd.n79 0.152939
R22360 gnd.n7768 gnd.n7767 0.152939
R22361 gnd.n7767 gnd.n7766 0.152939
R22362 gnd.n7766 gnd.n84 0.152939
R22363 gnd.n7762 gnd.n84 0.152939
R22364 gnd.n7762 gnd.n7761 0.152939
R22365 gnd.n7761 gnd.n7760 0.152939
R22366 gnd.n7760 gnd.n89 0.152939
R22367 gnd.n7756 gnd.n89 0.152939
R22368 gnd.n7756 gnd.n7755 0.152939
R22369 gnd.n7755 gnd.n7754 0.152939
R22370 gnd.n7754 gnd.n94 0.152939
R22371 gnd.n7750 gnd.n94 0.152939
R22372 gnd.n7750 gnd.n7749 0.152939
R22373 gnd.n7749 gnd.n7748 0.152939
R22374 gnd.n7748 gnd.n99 0.152939
R22375 gnd.n102 gnd.n99 0.152939
R22376 gnd.n4471 gnd.n1643 0.151415
R22377 gnd.n3445 gnd.n2645 0.151415
R22378 gnd.n309 gnd.n268 0.0889146
R22379 gnd.n2995 gnd.n2994 0.0889146
R22380 gnd.n5951 gnd.n5343 0.0767195
R22381 gnd.n5867 gnd.n5343 0.0767195
R22382 gnd.n7505 gnd.n252 0.0767195
R22383 gnd.n4643 gnd.n291 0.0767195
R22384 gnd.n300 gnd.n291 0.0767195
R22385 gnd.n7505 gnd.n267 0.0767195
R22386 gnd.n1212 gnd.n1175 0.0767195
R22387 gnd.n2898 gnd.n1184 0.0767195
R22388 gnd.n2898 gnd.n1185 0.0767195
R22389 gnd.n3202 gnd.n3201 0.0767195
R22390 gnd.n3203 gnd.n3202 0.0767195
R22391 gnd.n1175 gnd.n1155 0.0767195
R22392 gnd.n7492 gnd.n7491 0.0767195
R22393 gnd.n7491 gnd.n7490 0.0767195
R22394 gnd.n7785 gnd.n67 0.0767195
R22395 gnd.n7785 gnd.n7784 0.0767195
R22396 gnd.n3195 gnd.n3194 0.0695946
R22397 gnd.n3194 gnd.n2894 0.0695946
R22398 gnd.n2995 gnd.n2941 0.0645244
R22399 gnd.n1536 gnd.n268 0.0645244
R22400 gnd.n4896 gnd.n4895 0.063
R22401 gnd.n1693 gnd.n1692 0.063
R22402 gnd.n6459 gnd.n5163 0.0477147
R22403 gnd.n5617 gnd.n5513 0.0442063
R22404 gnd.n5631 gnd.n5513 0.0442063
R22405 gnd.n5632 gnd.n5631 0.0442063
R22406 gnd.n5633 gnd.n5632 0.0442063
R22407 gnd.n5633 gnd.n5501 0.0442063
R22408 gnd.n5647 gnd.n5501 0.0442063
R22409 gnd.n5648 gnd.n5647 0.0442063
R22410 gnd.n5649 gnd.n5648 0.0442063
R22411 gnd.n5649 gnd.n5488 0.0442063
R22412 gnd.n5745 gnd.n5488 0.0442063
R22413 gnd.n5748 gnd.n5747 0.0344674
R22414 gnd.n4475 gnd.n1649 0.0343753
R22415 gnd.n3444 gnd.n2646 0.0343753
R22416 gnd.n5481 gnd.n5480 0.0269946
R22417 gnd.n5758 gnd.n5478 0.0269946
R22418 gnd.n5757 gnd.n5479 0.0269946
R22419 gnd.n5777 gnd.n5460 0.0269946
R22420 gnd.n5779 gnd.n5778 0.0269946
R22421 gnd.n5780 gnd.n5458 0.0269946
R22422 gnd.n5787 gnd.n5783 0.0269946
R22423 gnd.n5786 gnd.n5785 0.0269946
R22424 gnd.n5784 gnd.n5437 0.0269946
R22425 gnd.n5811 gnd.n5438 0.0269946
R22426 gnd.n5810 gnd.n5439 0.0269946
R22427 gnd.n5843 gnd.n5413 0.0269946
R22428 gnd.n5845 gnd.n5844 0.0269946
R22429 gnd.n5846 gnd.n5405 0.0269946
R22430 gnd.n5409 gnd.n5406 0.0269946
R22431 gnd.n5856 gnd.n5407 0.0269946
R22432 gnd.n5855 gnd.n5408 0.0269946
R22433 gnd.n5901 gnd.n5381 0.0269946
R22434 gnd.n5903 gnd.n5902 0.0269946
R22435 gnd.n5912 gnd.n5374 0.0269946
R22436 gnd.n5914 gnd.n5913 0.0269946
R22437 gnd.n5915 gnd.n5372 0.0269946
R22438 gnd.n5922 gnd.n5918 0.0269946
R22439 gnd.n5921 gnd.n5920 0.0269946
R22440 gnd.n5919 gnd.n5351 0.0269946
R22441 gnd.n5944 gnd.n5352 0.0269946
R22442 gnd.n5943 gnd.n5353 0.0269946
R22443 gnd.n5986 gnd.n5278 0.0269946
R22444 gnd.n5988 gnd.n5987 0.0269946
R22445 gnd.n5997 gnd.n5271 0.0269946
R22446 gnd.n5999 gnd.n5998 0.0269946
R22447 gnd.n6000 gnd.n5269 0.0269946
R22448 gnd.n6006 gnd.n6003 0.0269946
R22449 gnd.n6005 gnd.n6004 0.0269946
R22450 gnd.n6031 gnd.n5248 0.0269946
R22451 gnd.n6030 gnd.n5249 0.0269946
R22452 gnd.n6057 gnd.n5234 0.0269946
R22453 gnd.n6059 gnd.n6058 0.0269946
R22454 gnd.n6060 gnd.n5220 0.0269946
R22455 gnd.n6082 gnd.n5218 0.0269946
R22456 gnd.n6084 gnd.n6083 0.0269946
R22457 gnd.n6086 gnd.n6085 0.0269946
R22458 gnd.n6095 gnd.n5210 0.0269946
R22459 gnd.n6097 gnd.n6096 0.0269946
R22460 gnd.n6098 gnd.n924 0.0269946
R22461 gnd.n5201 gnd.n925 0.0269946
R22462 gnd.n5203 gnd.n926 0.0269946
R22463 gnd.n6125 gnd.n6124 0.0269946
R22464 gnd.n6384 gnd.n949 0.0269946
R22465 gnd.n6386 gnd.n950 0.0269946
R22466 gnd.n6388 gnd.n951 0.0269946
R22467 gnd.n6390 gnd.n6389 0.0269946
R22468 gnd.n1694 gnd.n1693 0.0245515
R22469 gnd.n4895 gnd.n1327 0.0245515
R22470 gnd.n5747 gnd.n5746 0.0202011
R22471 gnd.n1695 gnd.n1694 0.0174377
R22472 gnd.n1703 gnd.n1695 0.0174377
R22473 gnd.n1703 gnd.n1702 0.0174377
R22474 gnd.n1702 gnd.n1696 0.0174377
R22475 gnd.n1696 gnd.n1680 0.0174377
R22476 gnd.n1711 gnd.n1680 0.0174377
R22477 gnd.n1713 gnd.n1711 0.0174377
R22478 gnd.n1713 gnd.n1712 0.0174377
R22479 gnd.n1712 gnd.n1675 0.0174377
R22480 gnd.n1722 gnd.n1675 0.0174377
R22481 gnd.n1722 gnd.n1721 0.0174377
R22482 gnd.n1721 gnd.n1676 0.0174377
R22483 gnd.n1676 gnd.n1671 0.0174377
R22484 gnd.n1730 gnd.n1671 0.0174377
R22485 gnd.n1732 gnd.n1730 0.0174377
R22486 gnd.n1732 gnd.n1731 0.0174377
R22487 gnd.n1731 gnd.n1666 0.0174377
R22488 gnd.n1741 gnd.n1666 0.0174377
R22489 gnd.n1741 gnd.n1740 0.0174377
R22490 gnd.n1740 gnd.n1667 0.0174377
R22491 gnd.n1667 gnd.n1662 0.0174377
R22492 gnd.n1749 gnd.n1662 0.0174377
R22493 gnd.n1751 gnd.n1749 0.0174377
R22494 gnd.n1751 gnd.n1750 0.0174377
R22495 gnd.n1750 gnd.n1657 0.0174377
R22496 gnd.n1760 gnd.n1657 0.0174377
R22497 gnd.n1760 gnd.n1759 0.0174377
R22498 gnd.n1759 gnd.n1658 0.0174377
R22499 gnd.n1658 gnd.n1653 0.0174377
R22500 gnd.n1768 gnd.n1653 0.0174377
R22501 gnd.n1770 gnd.n1768 0.0174377
R22502 gnd.n1770 gnd.n1769 0.0174377
R22503 gnd.n1769 gnd.n1648 0.0174377
R22504 gnd.n4476 gnd.n1648 0.0174377
R22505 gnd.n4476 gnd.n4475 0.0174377
R22506 gnd.n2725 gnd.n1327 0.0174377
R22507 gnd.n2727 gnd.n2725 0.0174377
R22508 gnd.n2835 gnd.n2727 0.0174377
R22509 gnd.n2835 gnd.n2834 0.0174377
R22510 gnd.n2834 gnd.n2728 0.0174377
R22511 gnd.n2831 gnd.n2728 0.0174377
R22512 gnd.n2831 gnd.n2830 0.0174377
R22513 gnd.n2830 gnd.n2738 0.0174377
R22514 gnd.n2827 gnd.n2738 0.0174377
R22515 gnd.n2827 gnd.n2826 0.0174377
R22516 gnd.n2826 gnd.n2743 0.0174377
R22517 gnd.n2823 gnd.n2743 0.0174377
R22518 gnd.n2823 gnd.n2822 0.0174377
R22519 gnd.n2822 gnd.n2749 0.0174377
R22520 gnd.n2819 gnd.n2749 0.0174377
R22521 gnd.n2819 gnd.n2818 0.0174377
R22522 gnd.n2818 gnd.n2753 0.0174377
R22523 gnd.n2815 gnd.n2753 0.0174377
R22524 gnd.n2815 gnd.n2814 0.0174377
R22525 gnd.n2814 gnd.n2760 0.0174377
R22526 gnd.n2811 gnd.n2760 0.0174377
R22527 gnd.n2811 gnd.n2810 0.0174377
R22528 gnd.n2810 gnd.n2766 0.0174377
R22529 gnd.n2807 gnd.n2766 0.0174377
R22530 gnd.n2807 gnd.n2806 0.0174377
R22531 gnd.n2806 gnd.n2772 0.0174377
R22532 gnd.n2803 gnd.n2772 0.0174377
R22533 gnd.n2803 gnd.n2802 0.0174377
R22534 gnd.n2802 gnd.n2776 0.0174377
R22535 gnd.n2799 gnd.n2776 0.0174377
R22536 gnd.n2799 gnd.n2798 0.0174377
R22537 gnd.n2798 gnd.n2785 0.0174377
R22538 gnd.n2795 gnd.n2785 0.0174377
R22539 gnd.n2795 gnd.n2794 0.0174377
R22540 gnd.n2794 gnd.n2646 0.0174377
R22541 gnd.n5746 gnd.n5745 0.0148637
R22542 gnd.n6382 gnd.n6126 0.0144266
R22543 gnd.n6383 gnd.n6382 0.0130679
R22544 gnd.n5748 gnd.n5481 0.00797283
R22545 gnd.n5480 gnd.n5478 0.00797283
R22546 gnd.n5758 gnd.n5757 0.00797283
R22547 gnd.n5479 gnd.n5460 0.00797283
R22548 gnd.n5778 gnd.n5777 0.00797283
R22549 gnd.n5780 gnd.n5779 0.00797283
R22550 gnd.n5783 gnd.n5458 0.00797283
R22551 gnd.n5787 gnd.n5786 0.00797283
R22552 gnd.n5785 gnd.n5784 0.00797283
R22553 gnd.n5438 gnd.n5437 0.00797283
R22554 gnd.n5811 gnd.n5810 0.00797283
R22555 gnd.n5439 gnd.n5413 0.00797283
R22556 gnd.n5844 gnd.n5843 0.00797283
R22557 gnd.n5846 gnd.n5845 0.00797283
R22558 gnd.n5409 gnd.n5405 0.00797283
R22559 gnd.n5407 gnd.n5406 0.00797283
R22560 gnd.n5856 gnd.n5855 0.00797283
R22561 gnd.n5408 gnd.n5381 0.00797283
R22562 gnd.n5903 gnd.n5901 0.00797283
R22563 gnd.n5902 gnd.n5374 0.00797283
R22564 gnd.n5913 gnd.n5912 0.00797283
R22565 gnd.n5915 gnd.n5914 0.00797283
R22566 gnd.n5918 gnd.n5372 0.00797283
R22567 gnd.n5922 gnd.n5921 0.00797283
R22568 gnd.n5920 gnd.n5919 0.00797283
R22569 gnd.n5352 gnd.n5351 0.00797283
R22570 gnd.n5944 gnd.n5943 0.00797283
R22571 gnd.n5353 gnd.n5278 0.00797283
R22572 gnd.n5988 gnd.n5986 0.00797283
R22573 gnd.n5987 gnd.n5271 0.00797283
R22574 gnd.n5998 gnd.n5997 0.00797283
R22575 gnd.n6000 gnd.n5999 0.00797283
R22576 gnd.n6003 gnd.n5269 0.00797283
R22577 gnd.n6006 gnd.n6005 0.00797283
R22578 gnd.n6004 gnd.n5248 0.00797283
R22579 gnd.n6031 gnd.n6030 0.00797283
R22580 gnd.n5249 gnd.n5234 0.00797283
R22581 gnd.n6058 gnd.n6057 0.00797283
R22582 gnd.n6060 gnd.n6059 0.00797283
R22583 gnd.n5220 gnd.n5218 0.00797283
R22584 gnd.n6083 gnd.n6082 0.00797283
R22585 gnd.n6086 gnd.n6084 0.00797283
R22586 gnd.n6085 gnd.n5210 0.00797283
R22587 gnd.n6096 gnd.n6095 0.00797283
R22588 gnd.n6098 gnd.n6097 0.00797283
R22589 gnd.n5201 gnd.n924 0.00797283
R22590 gnd.n5203 gnd.n925 0.00797283
R22591 gnd.n6124 gnd.n926 0.00797283
R22592 gnd.n6126 gnd.n6125 0.00797283
R22593 gnd.n6384 gnd.n6383 0.00797283
R22594 gnd.n6386 gnd.n949 0.00797283
R22595 gnd.n6388 gnd.n950 0.00797283
R22596 gnd.n6390 gnd.n951 0.00797283
R22597 gnd.n6389 gnd.n5163 0.00797283
R22598 gnd.n7491 gnd.n291 0.00507153
R22599 gnd.n3202 gnd.n2898 0.00507153
R22600 gnd.n1649 gnd.n1643 0.000838753
R22601 gnd.n3445 gnd.n3444 0.000838753
R22602 commonsourceibias.n35 commonsourceibias.t16 223.028
R22603 commonsourceibias.n128 commonsourceibias.t85 223.028
R22604 commonsourceibias.n217 commonsourceibias.t75 223.028
R22605 commonsourceibias.n364 commonsourceibias.t54 223.028
R22606 commonsourceibias.n305 commonsourceibias.t91 223.028
R22607 commonsourceibias.n499 commonsourceibias.t78 223.028
R22608 commonsourceibias.n99 commonsourceibias.t60 207.983
R22609 commonsourceibias.n192 commonsourceibias.t92 207.983
R22610 commonsourceibias.n281 commonsourceibias.t81 207.983
R22611 commonsourceibias.n430 commonsourceibias.t8 207.983
R22612 commonsourceibias.n476 commonsourceibias.t110 207.983
R22613 commonsourceibias.n565 commonsourceibias.t97 207.983
R22614 commonsourceibias.n97 commonsourceibias.t14 168.701
R22615 commonsourceibias.n91 commonsourceibias.t38 168.701
R22616 commonsourceibias.n17 commonsourceibias.t4 168.701
R22617 commonsourceibias.n83 commonsourceibias.t28 168.701
R22618 commonsourceibias.n77 commonsourceibias.t62 168.701
R22619 commonsourceibias.n22 commonsourceibias.t18 168.701
R22620 commonsourceibias.n69 commonsourceibias.t26 168.701
R22621 commonsourceibias.n63 commonsourceibias.t6 168.701
R22622 commonsourceibias.n25 commonsourceibias.t32 168.701
R22623 commonsourceibias.n27 commonsourceibias.t42 168.701
R22624 commonsourceibias.n29 commonsourceibias.t20 168.701
R22625 commonsourceibias.n46 commonsourceibias.t30 168.701
R22626 commonsourceibias.n40 commonsourceibias.t56 168.701
R22627 commonsourceibias.n34 commonsourceibias.t12 168.701
R22628 commonsourceibias.n190 commonsourceibias.t106 168.701
R22629 commonsourceibias.n184 commonsourceibias.t119 168.701
R22630 commonsourceibias.n5 commonsourceibias.t84 168.701
R22631 commonsourceibias.n176 commonsourceibias.t100 168.701
R22632 commonsourceibias.n170 commonsourceibias.t114 168.701
R22633 commonsourceibias.n10 commonsourceibias.t80 168.701
R22634 commonsourceibias.n162 commonsourceibias.t76 168.701
R22635 commonsourceibias.n156 commonsourceibias.t105 168.701
R22636 commonsourceibias.n118 commonsourceibias.t121 168.701
R22637 commonsourceibias.n120 commonsourceibias.t71 168.701
R22638 commonsourceibias.n122 commonsourceibias.t99 168.701
R22639 commonsourceibias.n139 commonsourceibias.t95 168.701
R22640 commonsourceibias.n133 commonsourceibias.t109 168.701
R22641 commonsourceibias.n127 commonsourceibias.t89 168.701
R22642 commonsourceibias.n216 commonsourceibias.t77 168.701
R22643 commonsourceibias.n222 commonsourceibias.t96 168.701
R22644 commonsourceibias.n228 commonsourceibias.t82 168.701
R22645 commonsourceibias.n211 commonsourceibias.t86 168.701
R22646 commonsourceibias.n209 commonsourceibias.t127 168.701
R22647 commonsourceibias.n207 commonsourceibias.t108 168.701
R22648 commonsourceibias.n245 commonsourceibias.t93 168.701
R22649 commonsourceibias.n251 commonsourceibias.t67 168.701
R22650 commonsourceibias.n204 commonsourceibias.t70 168.701
R22651 commonsourceibias.n259 commonsourceibias.t101 168.701
R22652 commonsourceibias.n265 commonsourceibias.t87 168.701
R22653 commonsourceibias.n199 commonsourceibias.t74 168.701
R22654 commonsourceibias.n273 commonsourceibias.t107 168.701
R22655 commonsourceibias.n279 commonsourceibias.t94 168.701
R22656 commonsourceibias.n363 commonsourceibias.t52 168.701
R22657 commonsourceibias.n369 commonsourceibias.t2 168.701
R22658 commonsourceibias.n375 commonsourceibias.t48 168.701
R22659 commonsourceibias.n358 commonsourceibias.t40 168.701
R22660 commonsourceibias.n356 commonsourceibias.t58 168.701
R22661 commonsourceibias.n354 commonsourceibias.t50 168.701
R22662 commonsourceibias.n392 commonsourceibias.t24 168.701
R22663 commonsourceibias.n398 commonsourceibias.t44 168.701
R22664 commonsourceibias.n400 commonsourceibias.t36 168.701
R22665 commonsourceibias.n407 commonsourceibias.t10 168.701
R22666 commonsourceibias.n413 commonsourceibias.t46 168.701
R22667 commonsourceibias.n415 commonsourceibias.t22 168.701
R22668 commonsourceibias.n422 commonsourceibias.t0 168.701
R22669 commonsourceibias.n428 commonsourceibias.t34 168.701
R22670 commonsourceibias.n474 commonsourceibias.t123 168.701
R22671 commonsourceibias.n468 commonsourceibias.t68 168.701
R22672 commonsourceibias.n461 commonsourceibias.t102 168.701
R22673 commonsourceibias.n459 commonsourceibias.t117 168.701
R22674 commonsourceibias.n453 commonsourceibias.t64 168.701
R22675 commonsourceibias.n446 commonsourceibias.t72 168.701
R22676 commonsourceibias.n444 commonsourceibias.t90 168.701
R22677 commonsourceibias.n304 commonsourceibias.t83 168.701
R22678 commonsourceibias.n310 commonsourceibias.t126 168.701
R22679 commonsourceibias.n316 commonsourceibias.t113 168.701
R22680 commonsourceibias.n299 commonsourceibias.t116 168.701
R22681 commonsourceibias.n297 commonsourceibias.t66 168.701
R22682 commonsourceibias.n295 commonsourceibias.t69 168.701
R22683 commonsourceibias.n333 commonsourceibias.t122 168.701
R22684 commonsourceibias.n498 commonsourceibias.t73 168.701
R22685 commonsourceibias.n504 commonsourceibias.t115 168.701
R22686 commonsourceibias.n510 commonsourceibias.t98 168.701
R22687 commonsourceibias.n493 commonsourceibias.t103 168.701
R22688 commonsourceibias.n491 commonsourceibias.t120 168.701
R22689 commonsourceibias.n489 commonsourceibias.t125 168.701
R22690 commonsourceibias.n527 commonsourceibias.t111 168.701
R22691 commonsourceibias.n533 commonsourceibias.t79 168.701
R22692 commonsourceibias.n535 commonsourceibias.t65 168.701
R22693 commonsourceibias.n542 commonsourceibias.t118 168.701
R22694 commonsourceibias.n548 commonsourceibias.t104 168.701
R22695 commonsourceibias.n550 commonsourceibias.t88 168.701
R22696 commonsourceibias.n557 commonsourceibias.t124 168.701
R22697 commonsourceibias.n563 commonsourceibias.t112 168.701
R22698 commonsourceibias.n36 commonsourceibias.n33 161.3
R22699 commonsourceibias.n38 commonsourceibias.n37 161.3
R22700 commonsourceibias.n39 commonsourceibias.n32 161.3
R22701 commonsourceibias.n42 commonsourceibias.n41 161.3
R22702 commonsourceibias.n43 commonsourceibias.n31 161.3
R22703 commonsourceibias.n45 commonsourceibias.n44 161.3
R22704 commonsourceibias.n47 commonsourceibias.n30 161.3
R22705 commonsourceibias.n49 commonsourceibias.n48 161.3
R22706 commonsourceibias.n51 commonsourceibias.n50 161.3
R22707 commonsourceibias.n52 commonsourceibias.n28 161.3
R22708 commonsourceibias.n54 commonsourceibias.n53 161.3
R22709 commonsourceibias.n56 commonsourceibias.n55 161.3
R22710 commonsourceibias.n57 commonsourceibias.n26 161.3
R22711 commonsourceibias.n59 commonsourceibias.n58 161.3
R22712 commonsourceibias.n61 commonsourceibias.n60 161.3
R22713 commonsourceibias.n62 commonsourceibias.n24 161.3
R22714 commonsourceibias.n65 commonsourceibias.n64 161.3
R22715 commonsourceibias.n66 commonsourceibias.n23 161.3
R22716 commonsourceibias.n68 commonsourceibias.n67 161.3
R22717 commonsourceibias.n70 commonsourceibias.n21 161.3
R22718 commonsourceibias.n72 commonsourceibias.n71 161.3
R22719 commonsourceibias.n73 commonsourceibias.n20 161.3
R22720 commonsourceibias.n75 commonsourceibias.n74 161.3
R22721 commonsourceibias.n76 commonsourceibias.n19 161.3
R22722 commonsourceibias.n79 commonsourceibias.n78 161.3
R22723 commonsourceibias.n80 commonsourceibias.n18 161.3
R22724 commonsourceibias.n82 commonsourceibias.n81 161.3
R22725 commonsourceibias.n84 commonsourceibias.n16 161.3
R22726 commonsourceibias.n86 commonsourceibias.n85 161.3
R22727 commonsourceibias.n87 commonsourceibias.n15 161.3
R22728 commonsourceibias.n89 commonsourceibias.n88 161.3
R22729 commonsourceibias.n90 commonsourceibias.n14 161.3
R22730 commonsourceibias.n93 commonsourceibias.n92 161.3
R22731 commonsourceibias.n94 commonsourceibias.n13 161.3
R22732 commonsourceibias.n96 commonsourceibias.n95 161.3
R22733 commonsourceibias.n98 commonsourceibias.n12 161.3
R22734 commonsourceibias.n129 commonsourceibias.n126 161.3
R22735 commonsourceibias.n131 commonsourceibias.n130 161.3
R22736 commonsourceibias.n132 commonsourceibias.n125 161.3
R22737 commonsourceibias.n135 commonsourceibias.n134 161.3
R22738 commonsourceibias.n136 commonsourceibias.n124 161.3
R22739 commonsourceibias.n138 commonsourceibias.n137 161.3
R22740 commonsourceibias.n140 commonsourceibias.n123 161.3
R22741 commonsourceibias.n142 commonsourceibias.n141 161.3
R22742 commonsourceibias.n144 commonsourceibias.n143 161.3
R22743 commonsourceibias.n145 commonsourceibias.n121 161.3
R22744 commonsourceibias.n147 commonsourceibias.n146 161.3
R22745 commonsourceibias.n149 commonsourceibias.n148 161.3
R22746 commonsourceibias.n150 commonsourceibias.n119 161.3
R22747 commonsourceibias.n152 commonsourceibias.n151 161.3
R22748 commonsourceibias.n154 commonsourceibias.n153 161.3
R22749 commonsourceibias.n155 commonsourceibias.n117 161.3
R22750 commonsourceibias.n158 commonsourceibias.n157 161.3
R22751 commonsourceibias.n159 commonsourceibias.n11 161.3
R22752 commonsourceibias.n161 commonsourceibias.n160 161.3
R22753 commonsourceibias.n163 commonsourceibias.n9 161.3
R22754 commonsourceibias.n165 commonsourceibias.n164 161.3
R22755 commonsourceibias.n166 commonsourceibias.n8 161.3
R22756 commonsourceibias.n168 commonsourceibias.n167 161.3
R22757 commonsourceibias.n169 commonsourceibias.n7 161.3
R22758 commonsourceibias.n172 commonsourceibias.n171 161.3
R22759 commonsourceibias.n173 commonsourceibias.n6 161.3
R22760 commonsourceibias.n175 commonsourceibias.n174 161.3
R22761 commonsourceibias.n177 commonsourceibias.n4 161.3
R22762 commonsourceibias.n179 commonsourceibias.n178 161.3
R22763 commonsourceibias.n180 commonsourceibias.n3 161.3
R22764 commonsourceibias.n182 commonsourceibias.n181 161.3
R22765 commonsourceibias.n183 commonsourceibias.n2 161.3
R22766 commonsourceibias.n186 commonsourceibias.n185 161.3
R22767 commonsourceibias.n187 commonsourceibias.n1 161.3
R22768 commonsourceibias.n189 commonsourceibias.n188 161.3
R22769 commonsourceibias.n191 commonsourceibias.n0 161.3
R22770 commonsourceibias.n280 commonsourceibias.n194 161.3
R22771 commonsourceibias.n278 commonsourceibias.n277 161.3
R22772 commonsourceibias.n276 commonsourceibias.n195 161.3
R22773 commonsourceibias.n275 commonsourceibias.n274 161.3
R22774 commonsourceibias.n272 commonsourceibias.n196 161.3
R22775 commonsourceibias.n271 commonsourceibias.n270 161.3
R22776 commonsourceibias.n269 commonsourceibias.n197 161.3
R22777 commonsourceibias.n268 commonsourceibias.n267 161.3
R22778 commonsourceibias.n266 commonsourceibias.n198 161.3
R22779 commonsourceibias.n264 commonsourceibias.n263 161.3
R22780 commonsourceibias.n262 commonsourceibias.n200 161.3
R22781 commonsourceibias.n261 commonsourceibias.n260 161.3
R22782 commonsourceibias.n258 commonsourceibias.n201 161.3
R22783 commonsourceibias.n257 commonsourceibias.n256 161.3
R22784 commonsourceibias.n255 commonsourceibias.n202 161.3
R22785 commonsourceibias.n254 commonsourceibias.n253 161.3
R22786 commonsourceibias.n252 commonsourceibias.n203 161.3
R22787 commonsourceibias.n250 commonsourceibias.n249 161.3
R22788 commonsourceibias.n248 commonsourceibias.n205 161.3
R22789 commonsourceibias.n247 commonsourceibias.n246 161.3
R22790 commonsourceibias.n244 commonsourceibias.n206 161.3
R22791 commonsourceibias.n243 commonsourceibias.n242 161.3
R22792 commonsourceibias.n241 commonsourceibias.n240 161.3
R22793 commonsourceibias.n239 commonsourceibias.n208 161.3
R22794 commonsourceibias.n238 commonsourceibias.n237 161.3
R22795 commonsourceibias.n236 commonsourceibias.n235 161.3
R22796 commonsourceibias.n234 commonsourceibias.n210 161.3
R22797 commonsourceibias.n233 commonsourceibias.n232 161.3
R22798 commonsourceibias.n231 commonsourceibias.n230 161.3
R22799 commonsourceibias.n229 commonsourceibias.n212 161.3
R22800 commonsourceibias.n227 commonsourceibias.n226 161.3
R22801 commonsourceibias.n225 commonsourceibias.n213 161.3
R22802 commonsourceibias.n224 commonsourceibias.n223 161.3
R22803 commonsourceibias.n221 commonsourceibias.n214 161.3
R22804 commonsourceibias.n220 commonsourceibias.n219 161.3
R22805 commonsourceibias.n218 commonsourceibias.n215 161.3
R22806 commonsourceibias.n429 commonsourceibias.n343 161.3
R22807 commonsourceibias.n427 commonsourceibias.n426 161.3
R22808 commonsourceibias.n425 commonsourceibias.n344 161.3
R22809 commonsourceibias.n424 commonsourceibias.n423 161.3
R22810 commonsourceibias.n421 commonsourceibias.n345 161.3
R22811 commonsourceibias.n420 commonsourceibias.n419 161.3
R22812 commonsourceibias.n418 commonsourceibias.n346 161.3
R22813 commonsourceibias.n417 commonsourceibias.n416 161.3
R22814 commonsourceibias.n414 commonsourceibias.n347 161.3
R22815 commonsourceibias.n412 commonsourceibias.n411 161.3
R22816 commonsourceibias.n410 commonsourceibias.n348 161.3
R22817 commonsourceibias.n409 commonsourceibias.n408 161.3
R22818 commonsourceibias.n406 commonsourceibias.n349 161.3
R22819 commonsourceibias.n405 commonsourceibias.n404 161.3
R22820 commonsourceibias.n403 commonsourceibias.n350 161.3
R22821 commonsourceibias.n402 commonsourceibias.n401 161.3
R22822 commonsourceibias.n399 commonsourceibias.n351 161.3
R22823 commonsourceibias.n397 commonsourceibias.n396 161.3
R22824 commonsourceibias.n395 commonsourceibias.n352 161.3
R22825 commonsourceibias.n394 commonsourceibias.n393 161.3
R22826 commonsourceibias.n391 commonsourceibias.n353 161.3
R22827 commonsourceibias.n390 commonsourceibias.n389 161.3
R22828 commonsourceibias.n388 commonsourceibias.n387 161.3
R22829 commonsourceibias.n386 commonsourceibias.n355 161.3
R22830 commonsourceibias.n385 commonsourceibias.n384 161.3
R22831 commonsourceibias.n383 commonsourceibias.n382 161.3
R22832 commonsourceibias.n381 commonsourceibias.n357 161.3
R22833 commonsourceibias.n380 commonsourceibias.n379 161.3
R22834 commonsourceibias.n378 commonsourceibias.n377 161.3
R22835 commonsourceibias.n376 commonsourceibias.n359 161.3
R22836 commonsourceibias.n374 commonsourceibias.n373 161.3
R22837 commonsourceibias.n372 commonsourceibias.n360 161.3
R22838 commonsourceibias.n371 commonsourceibias.n370 161.3
R22839 commonsourceibias.n368 commonsourceibias.n361 161.3
R22840 commonsourceibias.n367 commonsourceibias.n366 161.3
R22841 commonsourceibias.n365 commonsourceibias.n362 161.3
R22842 commonsourceibias.n335 commonsourceibias.n334 161.3
R22843 commonsourceibias.n332 commonsourceibias.n294 161.3
R22844 commonsourceibias.n331 commonsourceibias.n330 161.3
R22845 commonsourceibias.n329 commonsourceibias.n328 161.3
R22846 commonsourceibias.n327 commonsourceibias.n296 161.3
R22847 commonsourceibias.n326 commonsourceibias.n325 161.3
R22848 commonsourceibias.n324 commonsourceibias.n323 161.3
R22849 commonsourceibias.n322 commonsourceibias.n298 161.3
R22850 commonsourceibias.n321 commonsourceibias.n320 161.3
R22851 commonsourceibias.n319 commonsourceibias.n318 161.3
R22852 commonsourceibias.n317 commonsourceibias.n300 161.3
R22853 commonsourceibias.n315 commonsourceibias.n314 161.3
R22854 commonsourceibias.n313 commonsourceibias.n301 161.3
R22855 commonsourceibias.n312 commonsourceibias.n311 161.3
R22856 commonsourceibias.n309 commonsourceibias.n302 161.3
R22857 commonsourceibias.n308 commonsourceibias.n307 161.3
R22858 commonsourceibias.n306 commonsourceibias.n303 161.3
R22859 commonsourceibias.n441 commonsourceibias.n293 161.3
R22860 commonsourceibias.n475 commonsourceibias.n284 161.3
R22861 commonsourceibias.n473 commonsourceibias.n472 161.3
R22862 commonsourceibias.n471 commonsourceibias.n285 161.3
R22863 commonsourceibias.n470 commonsourceibias.n469 161.3
R22864 commonsourceibias.n467 commonsourceibias.n286 161.3
R22865 commonsourceibias.n466 commonsourceibias.n465 161.3
R22866 commonsourceibias.n464 commonsourceibias.n287 161.3
R22867 commonsourceibias.n463 commonsourceibias.n462 161.3
R22868 commonsourceibias.n460 commonsourceibias.n288 161.3
R22869 commonsourceibias.n458 commonsourceibias.n457 161.3
R22870 commonsourceibias.n456 commonsourceibias.n289 161.3
R22871 commonsourceibias.n455 commonsourceibias.n454 161.3
R22872 commonsourceibias.n452 commonsourceibias.n290 161.3
R22873 commonsourceibias.n451 commonsourceibias.n450 161.3
R22874 commonsourceibias.n449 commonsourceibias.n291 161.3
R22875 commonsourceibias.n448 commonsourceibias.n447 161.3
R22876 commonsourceibias.n445 commonsourceibias.n292 161.3
R22877 commonsourceibias.n443 commonsourceibias.n442 161.3
R22878 commonsourceibias.n564 commonsourceibias.n478 161.3
R22879 commonsourceibias.n562 commonsourceibias.n561 161.3
R22880 commonsourceibias.n560 commonsourceibias.n479 161.3
R22881 commonsourceibias.n559 commonsourceibias.n558 161.3
R22882 commonsourceibias.n556 commonsourceibias.n480 161.3
R22883 commonsourceibias.n555 commonsourceibias.n554 161.3
R22884 commonsourceibias.n553 commonsourceibias.n481 161.3
R22885 commonsourceibias.n552 commonsourceibias.n551 161.3
R22886 commonsourceibias.n549 commonsourceibias.n482 161.3
R22887 commonsourceibias.n547 commonsourceibias.n546 161.3
R22888 commonsourceibias.n545 commonsourceibias.n483 161.3
R22889 commonsourceibias.n544 commonsourceibias.n543 161.3
R22890 commonsourceibias.n541 commonsourceibias.n484 161.3
R22891 commonsourceibias.n540 commonsourceibias.n539 161.3
R22892 commonsourceibias.n538 commonsourceibias.n485 161.3
R22893 commonsourceibias.n537 commonsourceibias.n536 161.3
R22894 commonsourceibias.n534 commonsourceibias.n486 161.3
R22895 commonsourceibias.n532 commonsourceibias.n531 161.3
R22896 commonsourceibias.n530 commonsourceibias.n487 161.3
R22897 commonsourceibias.n529 commonsourceibias.n528 161.3
R22898 commonsourceibias.n526 commonsourceibias.n488 161.3
R22899 commonsourceibias.n525 commonsourceibias.n524 161.3
R22900 commonsourceibias.n523 commonsourceibias.n522 161.3
R22901 commonsourceibias.n521 commonsourceibias.n490 161.3
R22902 commonsourceibias.n520 commonsourceibias.n519 161.3
R22903 commonsourceibias.n518 commonsourceibias.n517 161.3
R22904 commonsourceibias.n516 commonsourceibias.n492 161.3
R22905 commonsourceibias.n515 commonsourceibias.n514 161.3
R22906 commonsourceibias.n513 commonsourceibias.n512 161.3
R22907 commonsourceibias.n511 commonsourceibias.n494 161.3
R22908 commonsourceibias.n509 commonsourceibias.n508 161.3
R22909 commonsourceibias.n507 commonsourceibias.n495 161.3
R22910 commonsourceibias.n506 commonsourceibias.n505 161.3
R22911 commonsourceibias.n503 commonsourceibias.n496 161.3
R22912 commonsourceibias.n502 commonsourceibias.n501 161.3
R22913 commonsourceibias.n500 commonsourceibias.n497 161.3
R22914 commonsourceibias.n111 commonsourceibias.n109 81.5057
R22915 commonsourceibias.n338 commonsourceibias.n336 81.5057
R22916 commonsourceibias.n111 commonsourceibias.n110 80.9324
R22917 commonsourceibias.n113 commonsourceibias.n112 80.9324
R22918 commonsourceibias.n115 commonsourceibias.n114 80.9324
R22919 commonsourceibias.n108 commonsourceibias.n107 80.9324
R22920 commonsourceibias.n106 commonsourceibias.n105 80.9324
R22921 commonsourceibias.n104 commonsourceibias.n103 80.9324
R22922 commonsourceibias.n102 commonsourceibias.n101 80.9324
R22923 commonsourceibias.n433 commonsourceibias.n432 80.9324
R22924 commonsourceibias.n435 commonsourceibias.n434 80.9324
R22925 commonsourceibias.n437 commonsourceibias.n436 80.9324
R22926 commonsourceibias.n439 commonsourceibias.n438 80.9324
R22927 commonsourceibias.n342 commonsourceibias.n341 80.9324
R22928 commonsourceibias.n340 commonsourceibias.n339 80.9324
R22929 commonsourceibias.n338 commonsourceibias.n337 80.9324
R22930 commonsourceibias.n100 commonsourceibias.n99 80.6037
R22931 commonsourceibias.n193 commonsourceibias.n192 80.6037
R22932 commonsourceibias.n282 commonsourceibias.n281 80.6037
R22933 commonsourceibias.n431 commonsourceibias.n430 80.6037
R22934 commonsourceibias.n477 commonsourceibias.n476 80.6037
R22935 commonsourceibias.n566 commonsourceibias.n565 80.6037
R22936 commonsourceibias.n85 commonsourceibias.n84 56.5617
R22937 commonsourceibias.n71 commonsourceibias.n70 56.5617
R22938 commonsourceibias.n62 commonsourceibias.n61 56.5617
R22939 commonsourceibias.n48 commonsourceibias.n47 56.5617
R22940 commonsourceibias.n178 commonsourceibias.n177 56.5617
R22941 commonsourceibias.n164 commonsourceibias.n163 56.5617
R22942 commonsourceibias.n155 commonsourceibias.n154 56.5617
R22943 commonsourceibias.n141 commonsourceibias.n140 56.5617
R22944 commonsourceibias.n230 commonsourceibias.n229 56.5617
R22945 commonsourceibias.n244 commonsourceibias.n243 56.5617
R22946 commonsourceibias.n253 commonsourceibias.n252 56.5617
R22947 commonsourceibias.n267 commonsourceibias.n266 56.5617
R22948 commonsourceibias.n377 commonsourceibias.n376 56.5617
R22949 commonsourceibias.n391 commonsourceibias.n390 56.5617
R22950 commonsourceibias.n401 commonsourceibias.n399 56.5617
R22951 commonsourceibias.n416 commonsourceibias.n414 56.5617
R22952 commonsourceibias.n462 commonsourceibias.n460 56.5617
R22953 commonsourceibias.n447 commonsourceibias.n445 56.5617
R22954 commonsourceibias.n318 commonsourceibias.n317 56.5617
R22955 commonsourceibias.n332 commonsourceibias.n331 56.5617
R22956 commonsourceibias.n512 commonsourceibias.n511 56.5617
R22957 commonsourceibias.n526 commonsourceibias.n525 56.5617
R22958 commonsourceibias.n536 commonsourceibias.n534 56.5617
R22959 commonsourceibias.n551 commonsourceibias.n549 56.5617
R22960 commonsourceibias.n76 commonsourceibias.n75 56.0773
R22961 commonsourceibias.n57 commonsourceibias.n56 56.0773
R22962 commonsourceibias.n169 commonsourceibias.n168 56.0773
R22963 commonsourceibias.n150 commonsourceibias.n149 56.0773
R22964 commonsourceibias.n239 commonsourceibias.n238 56.0773
R22965 commonsourceibias.n258 commonsourceibias.n257 56.0773
R22966 commonsourceibias.n386 commonsourceibias.n385 56.0773
R22967 commonsourceibias.n406 commonsourceibias.n405 56.0773
R22968 commonsourceibias.n452 commonsourceibias.n451 56.0773
R22969 commonsourceibias.n327 commonsourceibias.n326 56.0773
R22970 commonsourceibias.n521 commonsourceibias.n520 56.0773
R22971 commonsourceibias.n541 commonsourceibias.n540 56.0773
R22972 commonsourceibias.n99 commonsourceibias.n98 55.3321
R22973 commonsourceibias.n192 commonsourceibias.n191 55.3321
R22974 commonsourceibias.n281 commonsourceibias.n280 55.3321
R22975 commonsourceibias.n430 commonsourceibias.n429 55.3321
R22976 commonsourceibias.n476 commonsourceibias.n475 55.3321
R22977 commonsourceibias.n565 commonsourceibias.n564 55.3321
R22978 commonsourceibias.n90 commonsourceibias.n89 55.1086
R22979 commonsourceibias.n41 commonsourceibias.n31 55.1086
R22980 commonsourceibias.n183 commonsourceibias.n182 55.1086
R22981 commonsourceibias.n134 commonsourceibias.n124 55.1086
R22982 commonsourceibias.n223 commonsourceibias.n213 55.1086
R22983 commonsourceibias.n272 commonsourceibias.n271 55.1086
R22984 commonsourceibias.n370 commonsourceibias.n360 55.1086
R22985 commonsourceibias.n421 commonsourceibias.n420 55.1086
R22986 commonsourceibias.n467 commonsourceibias.n466 55.1086
R22987 commonsourceibias.n311 commonsourceibias.n301 55.1086
R22988 commonsourceibias.n505 commonsourceibias.n495 55.1086
R22989 commonsourceibias.n556 commonsourceibias.n555 55.1086
R22990 commonsourceibias.n35 commonsourceibias.n34 47.4592
R22991 commonsourceibias.n128 commonsourceibias.n127 47.4592
R22992 commonsourceibias.n217 commonsourceibias.n216 47.4592
R22993 commonsourceibias.n364 commonsourceibias.n363 47.4592
R22994 commonsourceibias.n305 commonsourceibias.n304 47.4592
R22995 commonsourceibias.n499 commonsourceibias.n498 47.4592
R22996 commonsourceibias.n218 commonsourceibias.n217 44.0436
R22997 commonsourceibias.n365 commonsourceibias.n364 44.0436
R22998 commonsourceibias.n306 commonsourceibias.n305 44.0436
R22999 commonsourceibias.n500 commonsourceibias.n499 44.0436
R23000 commonsourceibias.n36 commonsourceibias.n35 44.0436
R23001 commonsourceibias.n129 commonsourceibias.n128 44.0436
R23002 commonsourceibias.n92 commonsourceibias.n13 42.5146
R23003 commonsourceibias.n39 commonsourceibias.n38 42.5146
R23004 commonsourceibias.n185 commonsourceibias.n1 42.5146
R23005 commonsourceibias.n132 commonsourceibias.n131 42.5146
R23006 commonsourceibias.n221 commonsourceibias.n220 42.5146
R23007 commonsourceibias.n274 commonsourceibias.n195 42.5146
R23008 commonsourceibias.n368 commonsourceibias.n367 42.5146
R23009 commonsourceibias.n423 commonsourceibias.n344 42.5146
R23010 commonsourceibias.n469 commonsourceibias.n285 42.5146
R23011 commonsourceibias.n309 commonsourceibias.n308 42.5146
R23012 commonsourceibias.n503 commonsourceibias.n502 42.5146
R23013 commonsourceibias.n558 commonsourceibias.n479 42.5146
R23014 commonsourceibias.n78 commonsourceibias.n18 41.5458
R23015 commonsourceibias.n53 commonsourceibias.n52 41.5458
R23016 commonsourceibias.n171 commonsourceibias.n6 41.5458
R23017 commonsourceibias.n146 commonsourceibias.n145 41.5458
R23018 commonsourceibias.n235 commonsourceibias.n234 41.5458
R23019 commonsourceibias.n260 commonsourceibias.n200 41.5458
R23020 commonsourceibias.n382 commonsourceibias.n381 41.5458
R23021 commonsourceibias.n408 commonsourceibias.n348 41.5458
R23022 commonsourceibias.n454 commonsourceibias.n289 41.5458
R23023 commonsourceibias.n323 commonsourceibias.n322 41.5458
R23024 commonsourceibias.n517 commonsourceibias.n516 41.5458
R23025 commonsourceibias.n543 commonsourceibias.n483 41.5458
R23026 commonsourceibias.n68 commonsourceibias.n23 40.577
R23027 commonsourceibias.n64 commonsourceibias.n23 40.577
R23028 commonsourceibias.n161 commonsourceibias.n11 40.577
R23029 commonsourceibias.n157 commonsourceibias.n11 40.577
R23030 commonsourceibias.n246 commonsourceibias.n205 40.577
R23031 commonsourceibias.n250 commonsourceibias.n205 40.577
R23032 commonsourceibias.n393 commonsourceibias.n352 40.577
R23033 commonsourceibias.n397 commonsourceibias.n352 40.577
R23034 commonsourceibias.n443 commonsourceibias.n293 40.577
R23035 commonsourceibias.n334 commonsourceibias.n293 40.577
R23036 commonsourceibias.n528 commonsourceibias.n487 40.577
R23037 commonsourceibias.n532 commonsourceibias.n487 40.577
R23038 commonsourceibias.n82 commonsourceibias.n18 39.6083
R23039 commonsourceibias.n52 commonsourceibias.n51 39.6083
R23040 commonsourceibias.n175 commonsourceibias.n6 39.6083
R23041 commonsourceibias.n145 commonsourceibias.n144 39.6083
R23042 commonsourceibias.n234 commonsourceibias.n233 39.6083
R23043 commonsourceibias.n264 commonsourceibias.n200 39.6083
R23044 commonsourceibias.n381 commonsourceibias.n380 39.6083
R23045 commonsourceibias.n412 commonsourceibias.n348 39.6083
R23046 commonsourceibias.n458 commonsourceibias.n289 39.6083
R23047 commonsourceibias.n322 commonsourceibias.n321 39.6083
R23048 commonsourceibias.n516 commonsourceibias.n515 39.6083
R23049 commonsourceibias.n547 commonsourceibias.n483 39.6083
R23050 commonsourceibias.n96 commonsourceibias.n13 38.6395
R23051 commonsourceibias.n38 commonsourceibias.n33 38.6395
R23052 commonsourceibias.n189 commonsourceibias.n1 38.6395
R23053 commonsourceibias.n131 commonsourceibias.n126 38.6395
R23054 commonsourceibias.n220 commonsourceibias.n215 38.6395
R23055 commonsourceibias.n278 commonsourceibias.n195 38.6395
R23056 commonsourceibias.n367 commonsourceibias.n362 38.6395
R23057 commonsourceibias.n427 commonsourceibias.n344 38.6395
R23058 commonsourceibias.n473 commonsourceibias.n285 38.6395
R23059 commonsourceibias.n308 commonsourceibias.n303 38.6395
R23060 commonsourceibias.n502 commonsourceibias.n497 38.6395
R23061 commonsourceibias.n562 commonsourceibias.n479 38.6395
R23062 commonsourceibias.n89 commonsourceibias.n15 26.0455
R23063 commonsourceibias.n45 commonsourceibias.n31 26.0455
R23064 commonsourceibias.n182 commonsourceibias.n3 26.0455
R23065 commonsourceibias.n138 commonsourceibias.n124 26.0455
R23066 commonsourceibias.n227 commonsourceibias.n213 26.0455
R23067 commonsourceibias.n271 commonsourceibias.n197 26.0455
R23068 commonsourceibias.n374 commonsourceibias.n360 26.0455
R23069 commonsourceibias.n420 commonsourceibias.n346 26.0455
R23070 commonsourceibias.n466 commonsourceibias.n287 26.0455
R23071 commonsourceibias.n315 commonsourceibias.n301 26.0455
R23072 commonsourceibias.n509 commonsourceibias.n495 26.0455
R23073 commonsourceibias.n555 commonsourceibias.n481 26.0455
R23074 commonsourceibias.n75 commonsourceibias.n20 25.0767
R23075 commonsourceibias.n58 commonsourceibias.n57 25.0767
R23076 commonsourceibias.n168 commonsourceibias.n8 25.0767
R23077 commonsourceibias.n151 commonsourceibias.n150 25.0767
R23078 commonsourceibias.n240 commonsourceibias.n239 25.0767
R23079 commonsourceibias.n257 commonsourceibias.n202 25.0767
R23080 commonsourceibias.n387 commonsourceibias.n386 25.0767
R23081 commonsourceibias.n405 commonsourceibias.n350 25.0767
R23082 commonsourceibias.n451 commonsourceibias.n291 25.0767
R23083 commonsourceibias.n328 commonsourceibias.n327 25.0767
R23084 commonsourceibias.n522 commonsourceibias.n521 25.0767
R23085 commonsourceibias.n540 commonsourceibias.n485 25.0767
R23086 commonsourceibias.n71 commonsourceibias.n22 24.3464
R23087 commonsourceibias.n61 commonsourceibias.n25 24.3464
R23088 commonsourceibias.n164 commonsourceibias.n10 24.3464
R23089 commonsourceibias.n154 commonsourceibias.n118 24.3464
R23090 commonsourceibias.n243 commonsourceibias.n207 24.3464
R23091 commonsourceibias.n253 commonsourceibias.n204 24.3464
R23092 commonsourceibias.n390 commonsourceibias.n354 24.3464
R23093 commonsourceibias.n401 commonsourceibias.n400 24.3464
R23094 commonsourceibias.n447 commonsourceibias.n446 24.3464
R23095 commonsourceibias.n331 commonsourceibias.n295 24.3464
R23096 commonsourceibias.n525 commonsourceibias.n489 24.3464
R23097 commonsourceibias.n536 commonsourceibias.n535 24.3464
R23098 commonsourceibias.n85 commonsourceibias.n17 23.8546
R23099 commonsourceibias.n47 commonsourceibias.n46 23.8546
R23100 commonsourceibias.n178 commonsourceibias.n5 23.8546
R23101 commonsourceibias.n140 commonsourceibias.n139 23.8546
R23102 commonsourceibias.n229 commonsourceibias.n228 23.8546
R23103 commonsourceibias.n267 commonsourceibias.n199 23.8546
R23104 commonsourceibias.n376 commonsourceibias.n375 23.8546
R23105 commonsourceibias.n416 commonsourceibias.n415 23.8546
R23106 commonsourceibias.n462 commonsourceibias.n461 23.8546
R23107 commonsourceibias.n317 commonsourceibias.n316 23.8546
R23108 commonsourceibias.n511 commonsourceibias.n510 23.8546
R23109 commonsourceibias.n551 commonsourceibias.n550 23.8546
R23110 commonsourceibias.n98 commonsourceibias.n97 17.4607
R23111 commonsourceibias.n191 commonsourceibias.n190 17.4607
R23112 commonsourceibias.n280 commonsourceibias.n279 17.4607
R23113 commonsourceibias.n429 commonsourceibias.n428 17.4607
R23114 commonsourceibias.n475 commonsourceibias.n474 17.4607
R23115 commonsourceibias.n564 commonsourceibias.n563 17.4607
R23116 commonsourceibias.n84 commonsourceibias.n83 16.9689
R23117 commonsourceibias.n48 commonsourceibias.n29 16.9689
R23118 commonsourceibias.n177 commonsourceibias.n176 16.9689
R23119 commonsourceibias.n141 commonsourceibias.n122 16.9689
R23120 commonsourceibias.n230 commonsourceibias.n211 16.9689
R23121 commonsourceibias.n266 commonsourceibias.n265 16.9689
R23122 commonsourceibias.n377 commonsourceibias.n358 16.9689
R23123 commonsourceibias.n414 commonsourceibias.n413 16.9689
R23124 commonsourceibias.n460 commonsourceibias.n459 16.9689
R23125 commonsourceibias.n318 commonsourceibias.n299 16.9689
R23126 commonsourceibias.n512 commonsourceibias.n493 16.9689
R23127 commonsourceibias.n549 commonsourceibias.n548 16.9689
R23128 commonsourceibias.n70 commonsourceibias.n69 16.477
R23129 commonsourceibias.n63 commonsourceibias.n62 16.477
R23130 commonsourceibias.n163 commonsourceibias.n162 16.477
R23131 commonsourceibias.n156 commonsourceibias.n155 16.477
R23132 commonsourceibias.n245 commonsourceibias.n244 16.477
R23133 commonsourceibias.n252 commonsourceibias.n251 16.477
R23134 commonsourceibias.n392 commonsourceibias.n391 16.477
R23135 commonsourceibias.n399 commonsourceibias.n398 16.477
R23136 commonsourceibias.n445 commonsourceibias.n444 16.477
R23137 commonsourceibias.n333 commonsourceibias.n332 16.477
R23138 commonsourceibias.n527 commonsourceibias.n526 16.477
R23139 commonsourceibias.n534 commonsourceibias.n533 16.477
R23140 commonsourceibias.n77 commonsourceibias.n76 15.9852
R23141 commonsourceibias.n56 commonsourceibias.n27 15.9852
R23142 commonsourceibias.n170 commonsourceibias.n169 15.9852
R23143 commonsourceibias.n149 commonsourceibias.n120 15.9852
R23144 commonsourceibias.n238 commonsourceibias.n209 15.9852
R23145 commonsourceibias.n259 commonsourceibias.n258 15.9852
R23146 commonsourceibias.n385 commonsourceibias.n356 15.9852
R23147 commonsourceibias.n407 commonsourceibias.n406 15.9852
R23148 commonsourceibias.n453 commonsourceibias.n452 15.9852
R23149 commonsourceibias.n326 commonsourceibias.n297 15.9852
R23150 commonsourceibias.n520 commonsourceibias.n491 15.9852
R23151 commonsourceibias.n542 commonsourceibias.n541 15.9852
R23152 commonsourceibias.n91 commonsourceibias.n90 15.4934
R23153 commonsourceibias.n41 commonsourceibias.n40 15.4934
R23154 commonsourceibias.n184 commonsourceibias.n183 15.4934
R23155 commonsourceibias.n134 commonsourceibias.n133 15.4934
R23156 commonsourceibias.n223 commonsourceibias.n222 15.4934
R23157 commonsourceibias.n273 commonsourceibias.n272 15.4934
R23158 commonsourceibias.n370 commonsourceibias.n369 15.4934
R23159 commonsourceibias.n422 commonsourceibias.n421 15.4934
R23160 commonsourceibias.n468 commonsourceibias.n467 15.4934
R23161 commonsourceibias.n311 commonsourceibias.n310 15.4934
R23162 commonsourceibias.n505 commonsourceibias.n504 15.4934
R23163 commonsourceibias.n557 commonsourceibias.n556 15.4934
R23164 commonsourceibias.n102 commonsourceibias.n100 13.2663
R23165 commonsourceibias.n433 commonsourceibias.n431 13.2663
R23166 commonsourceibias.n568 commonsourceibias.n283 12.2777
R23167 commonsourceibias.n568 commonsourceibias.n567 10.3347
R23168 commonsourceibias.n159 commonsourceibias.n116 9.50363
R23169 commonsourceibias.n441 commonsourceibias.n440 9.50363
R23170 commonsourceibias.n92 commonsourceibias.n91 9.09948
R23171 commonsourceibias.n40 commonsourceibias.n39 9.09948
R23172 commonsourceibias.n185 commonsourceibias.n184 9.09948
R23173 commonsourceibias.n133 commonsourceibias.n132 9.09948
R23174 commonsourceibias.n222 commonsourceibias.n221 9.09948
R23175 commonsourceibias.n274 commonsourceibias.n273 9.09948
R23176 commonsourceibias.n369 commonsourceibias.n368 9.09948
R23177 commonsourceibias.n423 commonsourceibias.n422 9.09948
R23178 commonsourceibias.n469 commonsourceibias.n468 9.09948
R23179 commonsourceibias.n310 commonsourceibias.n309 9.09948
R23180 commonsourceibias.n504 commonsourceibias.n503 9.09948
R23181 commonsourceibias.n558 commonsourceibias.n557 9.09948
R23182 commonsourceibias.n283 commonsourceibias.n193 8.79261
R23183 commonsourceibias.n567 commonsourceibias.n477 8.79261
R23184 commonsourceibias.n78 commonsourceibias.n77 8.60764
R23185 commonsourceibias.n53 commonsourceibias.n27 8.60764
R23186 commonsourceibias.n171 commonsourceibias.n170 8.60764
R23187 commonsourceibias.n146 commonsourceibias.n120 8.60764
R23188 commonsourceibias.n235 commonsourceibias.n209 8.60764
R23189 commonsourceibias.n260 commonsourceibias.n259 8.60764
R23190 commonsourceibias.n382 commonsourceibias.n356 8.60764
R23191 commonsourceibias.n408 commonsourceibias.n407 8.60764
R23192 commonsourceibias.n454 commonsourceibias.n453 8.60764
R23193 commonsourceibias.n323 commonsourceibias.n297 8.60764
R23194 commonsourceibias.n517 commonsourceibias.n491 8.60764
R23195 commonsourceibias.n543 commonsourceibias.n542 8.60764
R23196 commonsourceibias.n69 commonsourceibias.n68 8.11581
R23197 commonsourceibias.n64 commonsourceibias.n63 8.11581
R23198 commonsourceibias.n162 commonsourceibias.n161 8.11581
R23199 commonsourceibias.n157 commonsourceibias.n156 8.11581
R23200 commonsourceibias.n246 commonsourceibias.n245 8.11581
R23201 commonsourceibias.n251 commonsourceibias.n250 8.11581
R23202 commonsourceibias.n393 commonsourceibias.n392 8.11581
R23203 commonsourceibias.n398 commonsourceibias.n397 8.11581
R23204 commonsourceibias.n444 commonsourceibias.n443 8.11581
R23205 commonsourceibias.n334 commonsourceibias.n333 8.11581
R23206 commonsourceibias.n528 commonsourceibias.n527 8.11581
R23207 commonsourceibias.n533 commonsourceibias.n532 8.11581
R23208 commonsourceibias.n83 commonsourceibias.n82 7.62397
R23209 commonsourceibias.n51 commonsourceibias.n29 7.62397
R23210 commonsourceibias.n176 commonsourceibias.n175 7.62397
R23211 commonsourceibias.n144 commonsourceibias.n122 7.62397
R23212 commonsourceibias.n233 commonsourceibias.n211 7.62397
R23213 commonsourceibias.n265 commonsourceibias.n264 7.62397
R23214 commonsourceibias.n380 commonsourceibias.n358 7.62397
R23215 commonsourceibias.n413 commonsourceibias.n412 7.62397
R23216 commonsourceibias.n459 commonsourceibias.n458 7.62397
R23217 commonsourceibias.n321 commonsourceibias.n299 7.62397
R23218 commonsourceibias.n515 commonsourceibias.n493 7.62397
R23219 commonsourceibias.n548 commonsourceibias.n547 7.62397
R23220 commonsourceibias.n97 commonsourceibias.n96 7.13213
R23221 commonsourceibias.n34 commonsourceibias.n33 7.13213
R23222 commonsourceibias.n190 commonsourceibias.n189 7.13213
R23223 commonsourceibias.n127 commonsourceibias.n126 7.13213
R23224 commonsourceibias.n216 commonsourceibias.n215 7.13213
R23225 commonsourceibias.n279 commonsourceibias.n278 7.13213
R23226 commonsourceibias.n363 commonsourceibias.n362 7.13213
R23227 commonsourceibias.n428 commonsourceibias.n427 7.13213
R23228 commonsourceibias.n474 commonsourceibias.n473 7.13213
R23229 commonsourceibias.n304 commonsourceibias.n303 7.13213
R23230 commonsourceibias.n498 commonsourceibias.n497 7.13213
R23231 commonsourceibias.n563 commonsourceibias.n562 7.13213
R23232 commonsourceibias.n283 commonsourceibias.n282 5.06534
R23233 commonsourceibias.n567 commonsourceibias.n566 5.06534
R23234 commonsourceibias commonsourceibias.n568 4.04308
R23235 commonsourceibias.n109 commonsourceibias.t13 2.82907
R23236 commonsourceibias.n109 commonsourceibias.t17 2.82907
R23237 commonsourceibias.n110 commonsourceibias.t31 2.82907
R23238 commonsourceibias.n110 commonsourceibias.t57 2.82907
R23239 commonsourceibias.n112 commonsourceibias.t43 2.82907
R23240 commonsourceibias.n112 commonsourceibias.t21 2.82907
R23241 commonsourceibias.n114 commonsourceibias.t7 2.82907
R23242 commonsourceibias.n114 commonsourceibias.t33 2.82907
R23243 commonsourceibias.n107 commonsourceibias.t19 2.82907
R23244 commonsourceibias.n107 commonsourceibias.t27 2.82907
R23245 commonsourceibias.n105 commonsourceibias.t29 2.82907
R23246 commonsourceibias.n105 commonsourceibias.t63 2.82907
R23247 commonsourceibias.n103 commonsourceibias.t39 2.82907
R23248 commonsourceibias.n103 commonsourceibias.t5 2.82907
R23249 commonsourceibias.n101 commonsourceibias.t61 2.82907
R23250 commonsourceibias.n101 commonsourceibias.t15 2.82907
R23251 commonsourceibias.n432 commonsourceibias.t35 2.82907
R23252 commonsourceibias.n432 commonsourceibias.t9 2.82907
R23253 commonsourceibias.n434 commonsourceibias.t23 2.82907
R23254 commonsourceibias.n434 commonsourceibias.t1 2.82907
R23255 commonsourceibias.n436 commonsourceibias.t11 2.82907
R23256 commonsourceibias.n436 commonsourceibias.t47 2.82907
R23257 commonsourceibias.n438 commonsourceibias.t45 2.82907
R23258 commonsourceibias.n438 commonsourceibias.t37 2.82907
R23259 commonsourceibias.n341 commonsourceibias.t51 2.82907
R23260 commonsourceibias.n341 commonsourceibias.t25 2.82907
R23261 commonsourceibias.n339 commonsourceibias.t41 2.82907
R23262 commonsourceibias.n339 commonsourceibias.t59 2.82907
R23263 commonsourceibias.n337 commonsourceibias.t3 2.82907
R23264 commonsourceibias.n337 commonsourceibias.t49 2.82907
R23265 commonsourceibias.n336 commonsourceibias.t55 2.82907
R23266 commonsourceibias.n336 commonsourceibias.t53 2.82907
R23267 commonsourceibias.n17 commonsourceibias.n15 0.738255
R23268 commonsourceibias.n46 commonsourceibias.n45 0.738255
R23269 commonsourceibias.n5 commonsourceibias.n3 0.738255
R23270 commonsourceibias.n139 commonsourceibias.n138 0.738255
R23271 commonsourceibias.n228 commonsourceibias.n227 0.738255
R23272 commonsourceibias.n199 commonsourceibias.n197 0.738255
R23273 commonsourceibias.n375 commonsourceibias.n374 0.738255
R23274 commonsourceibias.n415 commonsourceibias.n346 0.738255
R23275 commonsourceibias.n461 commonsourceibias.n287 0.738255
R23276 commonsourceibias.n316 commonsourceibias.n315 0.738255
R23277 commonsourceibias.n510 commonsourceibias.n509 0.738255
R23278 commonsourceibias.n550 commonsourceibias.n481 0.738255
R23279 commonsourceibias.n104 commonsourceibias.n102 0.573776
R23280 commonsourceibias.n106 commonsourceibias.n104 0.573776
R23281 commonsourceibias.n108 commonsourceibias.n106 0.573776
R23282 commonsourceibias.n115 commonsourceibias.n113 0.573776
R23283 commonsourceibias.n113 commonsourceibias.n111 0.573776
R23284 commonsourceibias.n340 commonsourceibias.n338 0.573776
R23285 commonsourceibias.n342 commonsourceibias.n340 0.573776
R23286 commonsourceibias.n439 commonsourceibias.n437 0.573776
R23287 commonsourceibias.n437 commonsourceibias.n435 0.573776
R23288 commonsourceibias.n435 commonsourceibias.n433 0.573776
R23289 commonsourceibias.n116 commonsourceibias.n108 0.287138
R23290 commonsourceibias.n116 commonsourceibias.n115 0.287138
R23291 commonsourceibias.n440 commonsourceibias.n342 0.287138
R23292 commonsourceibias.n440 commonsourceibias.n439 0.287138
R23293 commonsourceibias.n100 commonsourceibias.n12 0.285035
R23294 commonsourceibias.n193 commonsourceibias.n0 0.285035
R23295 commonsourceibias.n282 commonsourceibias.n194 0.285035
R23296 commonsourceibias.n431 commonsourceibias.n343 0.285035
R23297 commonsourceibias.n477 commonsourceibias.n284 0.285035
R23298 commonsourceibias.n566 commonsourceibias.n478 0.285035
R23299 commonsourceibias.n22 commonsourceibias.n20 0.246418
R23300 commonsourceibias.n58 commonsourceibias.n25 0.246418
R23301 commonsourceibias.n10 commonsourceibias.n8 0.246418
R23302 commonsourceibias.n151 commonsourceibias.n118 0.246418
R23303 commonsourceibias.n240 commonsourceibias.n207 0.246418
R23304 commonsourceibias.n204 commonsourceibias.n202 0.246418
R23305 commonsourceibias.n387 commonsourceibias.n354 0.246418
R23306 commonsourceibias.n400 commonsourceibias.n350 0.246418
R23307 commonsourceibias.n446 commonsourceibias.n291 0.246418
R23308 commonsourceibias.n328 commonsourceibias.n295 0.246418
R23309 commonsourceibias.n522 commonsourceibias.n489 0.246418
R23310 commonsourceibias.n535 commonsourceibias.n485 0.246418
R23311 commonsourceibias.n95 commonsourceibias.n12 0.189894
R23312 commonsourceibias.n95 commonsourceibias.n94 0.189894
R23313 commonsourceibias.n94 commonsourceibias.n93 0.189894
R23314 commonsourceibias.n93 commonsourceibias.n14 0.189894
R23315 commonsourceibias.n88 commonsourceibias.n14 0.189894
R23316 commonsourceibias.n88 commonsourceibias.n87 0.189894
R23317 commonsourceibias.n87 commonsourceibias.n86 0.189894
R23318 commonsourceibias.n86 commonsourceibias.n16 0.189894
R23319 commonsourceibias.n81 commonsourceibias.n16 0.189894
R23320 commonsourceibias.n81 commonsourceibias.n80 0.189894
R23321 commonsourceibias.n80 commonsourceibias.n79 0.189894
R23322 commonsourceibias.n79 commonsourceibias.n19 0.189894
R23323 commonsourceibias.n74 commonsourceibias.n19 0.189894
R23324 commonsourceibias.n74 commonsourceibias.n73 0.189894
R23325 commonsourceibias.n73 commonsourceibias.n72 0.189894
R23326 commonsourceibias.n72 commonsourceibias.n21 0.189894
R23327 commonsourceibias.n67 commonsourceibias.n21 0.189894
R23328 commonsourceibias.n67 commonsourceibias.n66 0.189894
R23329 commonsourceibias.n66 commonsourceibias.n65 0.189894
R23330 commonsourceibias.n65 commonsourceibias.n24 0.189894
R23331 commonsourceibias.n60 commonsourceibias.n24 0.189894
R23332 commonsourceibias.n60 commonsourceibias.n59 0.189894
R23333 commonsourceibias.n59 commonsourceibias.n26 0.189894
R23334 commonsourceibias.n55 commonsourceibias.n26 0.189894
R23335 commonsourceibias.n55 commonsourceibias.n54 0.189894
R23336 commonsourceibias.n54 commonsourceibias.n28 0.189894
R23337 commonsourceibias.n50 commonsourceibias.n28 0.189894
R23338 commonsourceibias.n50 commonsourceibias.n49 0.189894
R23339 commonsourceibias.n49 commonsourceibias.n30 0.189894
R23340 commonsourceibias.n44 commonsourceibias.n30 0.189894
R23341 commonsourceibias.n44 commonsourceibias.n43 0.189894
R23342 commonsourceibias.n43 commonsourceibias.n42 0.189894
R23343 commonsourceibias.n42 commonsourceibias.n32 0.189894
R23344 commonsourceibias.n37 commonsourceibias.n32 0.189894
R23345 commonsourceibias.n37 commonsourceibias.n36 0.189894
R23346 commonsourceibias.n158 commonsourceibias.n117 0.189894
R23347 commonsourceibias.n153 commonsourceibias.n117 0.189894
R23348 commonsourceibias.n153 commonsourceibias.n152 0.189894
R23349 commonsourceibias.n152 commonsourceibias.n119 0.189894
R23350 commonsourceibias.n148 commonsourceibias.n119 0.189894
R23351 commonsourceibias.n148 commonsourceibias.n147 0.189894
R23352 commonsourceibias.n147 commonsourceibias.n121 0.189894
R23353 commonsourceibias.n143 commonsourceibias.n121 0.189894
R23354 commonsourceibias.n143 commonsourceibias.n142 0.189894
R23355 commonsourceibias.n142 commonsourceibias.n123 0.189894
R23356 commonsourceibias.n137 commonsourceibias.n123 0.189894
R23357 commonsourceibias.n137 commonsourceibias.n136 0.189894
R23358 commonsourceibias.n136 commonsourceibias.n135 0.189894
R23359 commonsourceibias.n135 commonsourceibias.n125 0.189894
R23360 commonsourceibias.n130 commonsourceibias.n125 0.189894
R23361 commonsourceibias.n130 commonsourceibias.n129 0.189894
R23362 commonsourceibias.n188 commonsourceibias.n0 0.189894
R23363 commonsourceibias.n188 commonsourceibias.n187 0.189894
R23364 commonsourceibias.n187 commonsourceibias.n186 0.189894
R23365 commonsourceibias.n186 commonsourceibias.n2 0.189894
R23366 commonsourceibias.n181 commonsourceibias.n2 0.189894
R23367 commonsourceibias.n181 commonsourceibias.n180 0.189894
R23368 commonsourceibias.n180 commonsourceibias.n179 0.189894
R23369 commonsourceibias.n179 commonsourceibias.n4 0.189894
R23370 commonsourceibias.n174 commonsourceibias.n4 0.189894
R23371 commonsourceibias.n174 commonsourceibias.n173 0.189894
R23372 commonsourceibias.n173 commonsourceibias.n172 0.189894
R23373 commonsourceibias.n172 commonsourceibias.n7 0.189894
R23374 commonsourceibias.n167 commonsourceibias.n7 0.189894
R23375 commonsourceibias.n167 commonsourceibias.n166 0.189894
R23376 commonsourceibias.n166 commonsourceibias.n165 0.189894
R23377 commonsourceibias.n165 commonsourceibias.n9 0.189894
R23378 commonsourceibias.n160 commonsourceibias.n9 0.189894
R23379 commonsourceibias.n277 commonsourceibias.n194 0.189894
R23380 commonsourceibias.n277 commonsourceibias.n276 0.189894
R23381 commonsourceibias.n276 commonsourceibias.n275 0.189894
R23382 commonsourceibias.n275 commonsourceibias.n196 0.189894
R23383 commonsourceibias.n270 commonsourceibias.n196 0.189894
R23384 commonsourceibias.n270 commonsourceibias.n269 0.189894
R23385 commonsourceibias.n269 commonsourceibias.n268 0.189894
R23386 commonsourceibias.n268 commonsourceibias.n198 0.189894
R23387 commonsourceibias.n263 commonsourceibias.n198 0.189894
R23388 commonsourceibias.n263 commonsourceibias.n262 0.189894
R23389 commonsourceibias.n262 commonsourceibias.n261 0.189894
R23390 commonsourceibias.n261 commonsourceibias.n201 0.189894
R23391 commonsourceibias.n256 commonsourceibias.n201 0.189894
R23392 commonsourceibias.n256 commonsourceibias.n255 0.189894
R23393 commonsourceibias.n255 commonsourceibias.n254 0.189894
R23394 commonsourceibias.n254 commonsourceibias.n203 0.189894
R23395 commonsourceibias.n249 commonsourceibias.n203 0.189894
R23396 commonsourceibias.n249 commonsourceibias.n248 0.189894
R23397 commonsourceibias.n248 commonsourceibias.n247 0.189894
R23398 commonsourceibias.n247 commonsourceibias.n206 0.189894
R23399 commonsourceibias.n242 commonsourceibias.n206 0.189894
R23400 commonsourceibias.n242 commonsourceibias.n241 0.189894
R23401 commonsourceibias.n241 commonsourceibias.n208 0.189894
R23402 commonsourceibias.n237 commonsourceibias.n208 0.189894
R23403 commonsourceibias.n237 commonsourceibias.n236 0.189894
R23404 commonsourceibias.n236 commonsourceibias.n210 0.189894
R23405 commonsourceibias.n232 commonsourceibias.n210 0.189894
R23406 commonsourceibias.n232 commonsourceibias.n231 0.189894
R23407 commonsourceibias.n231 commonsourceibias.n212 0.189894
R23408 commonsourceibias.n226 commonsourceibias.n212 0.189894
R23409 commonsourceibias.n226 commonsourceibias.n225 0.189894
R23410 commonsourceibias.n225 commonsourceibias.n224 0.189894
R23411 commonsourceibias.n224 commonsourceibias.n214 0.189894
R23412 commonsourceibias.n219 commonsourceibias.n214 0.189894
R23413 commonsourceibias.n219 commonsourceibias.n218 0.189894
R23414 commonsourceibias.n366 commonsourceibias.n365 0.189894
R23415 commonsourceibias.n366 commonsourceibias.n361 0.189894
R23416 commonsourceibias.n371 commonsourceibias.n361 0.189894
R23417 commonsourceibias.n372 commonsourceibias.n371 0.189894
R23418 commonsourceibias.n373 commonsourceibias.n372 0.189894
R23419 commonsourceibias.n373 commonsourceibias.n359 0.189894
R23420 commonsourceibias.n378 commonsourceibias.n359 0.189894
R23421 commonsourceibias.n379 commonsourceibias.n378 0.189894
R23422 commonsourceibias.n379 commonsourceibias.n357 0.189894
R23423 commonsourceibias.n383 commonsourceibias.n357 0.189894
R23424 commonsourceibias.n384 commonsourceibias.n383 0.189894
R23425 commonsourceibias.n384 commonsourceibias.n355 0.189894
R23426 commonsourceibias.n388 commonsourceibias.n355 0.189894
R23427 commonsourceibias.n389 commonsourceibias.n388 0.189894
R23428 commonsourceibias.n389 commonsourceibias.n353 0.189894
R23429 commonsourceibias.n394 commonsourceibias.n353 0.189894
R23430 commonsourceibias.n395 commonsourceibias.n394 0.189894
R23431 commonsourceibias.n396 commonsourceibias.n395 0.189894
R23432 commonsourceibias.n396 commonsourceibias.n351 0.189894
R23433 commonsourceibias.n402 commonsourceibias.n351 0.189894
R23434 commonsourceibias.n403 commonsourceibias.n402 0.189894
R23435 commonsourceibias.n404 commonsourceibias.n403 0.189894
R23436 commonsourceibias.n404 commonsourceibias.n349 0.189894
R23437 commonsourceibias.n409 commonsourceibias.n349 0.189894
R23438 commonsourceibias.n410 commonsourceibias.n409 0.189894
R23439 commonsourceibias.n411 commonsourceibias.n410 0.189894
R23440 commonsourceibias.n411 commonsourceibias.n347 0.189894
R23441 commonsourceibias.n417 commonsourceibias.n347 0.189894
R23442 commonsourceibias.n418 commonsourceibias.n417 0.189894
R23443 commonsourceibias.n419 commonsourceibias.n418 0.189894
R23444 commonsourceibias.n419 commonsourceibias.n345 0.189894
R23445 commonsourceibias.n424 commonsourceibias.n345 0.189894
R23446 commonsourceibias.n425 commonsourceibias.n424 0.189894
R23447 commonsourceibias.n426 commonsourceibias.n425 0.189894
R23448 commonsourceibias.n426 commonsourceibias.n343 0.189894
R23449 commonsourceibias.n307 commonsourceibias.n306 0.189894
R23450 commonsourceibias.n307 commonsourceibias.n302 0.189894
R23451 commonsourceibias.n312 commonsourceibias.n302 0.189894
R23452 commonsourceibias.n313 commonsourceibias.n312 0.189894
R23453 commonsourceibias.n314 commonsourceibias.n313 0.189894
R23454 commonsourceibias.n314 commonsourceibias.n300 0.189894
R23455 commonsourceibias.n319 commonsourceibias.n300 0.189894
R23456 commonsourceibias.n320 commonsourceibias.n319 0.189894
R23457 commonsourceibias.n320 commonsourceibias.n298 0.189894
R23458 commonsourceibias.n324 commonsourceibias.n298 0.189894
R23459 commonsourceibias.n325 commonsourceibias.n324 0.189894
R23460 commonsourceibias.n325 commonsourceibias.n296 0.189894
R23461 commonsourceibias.n329 commonsourceibias.n296 0.189894
R23462 commonsourceibias.n330 commonsourceibias.n329 0.189894
R23463 commonsourceibias.n330 commonsourceibias.n294 0.189894
R23464 commonsourceibias.n335 commonsourceibias.n294 0.189894
R23465 commonsourceibias.n442 commonsourceibias.n292 0.189894
R23466 commonsourceibias.n448 commonsourceibias.n292 0.189894
R23467 commonsourceibias.n449 commonsourceibias.n448 0.189894
R23468 commonsourceibias.n450 commonsourceibias.n449 0.189894
R23469 commonsourceibias.n450 commonsourceibias.n290 0.189894
R23470 commonsourceibias.n455 commonsourceibias.n290 0.189894
R23471 commonsourceibias.n456 commonsourceibias.n455 0.189894
R23472 commonsourceibias.n457 commonsourceibias.n456 0.189894
R23473 commonsourceibias.n457 commonsourceibias.n288 0.189894
R23474 commonsourceibias.n463 commonsourceibias.n288 0.189894
R23475 commonsourceibias.n464 commonsourceibias.n463 0.189894
R23476 commonsourceibias.n465 commonsourceibias.n464 0.189894
R23477 commonsourceibias.n465 commonsourceibias.n286 0.189894
R23478 commonsourceibias.n470 commonsourceibias.n286 0.189894
R23479 commonsourceibias.n471 commonsourceibias.n470 0.189894
R23480 commonsourceibias.n472 commonsourceibias.n471 0.189894
R23481 commonsourceibias.n472 commonsourceibias.n284 0.189894
R23482 commonsourceibias.n501 commonsourceibias.n500 0.189894
R23483 commonsourceibias.n501 commonsourceibias.n496 0.189894
R23484 commonsourceibias.n506 commonsourceibias.n496 0.189894
R23485 commonsourceibias.n507 commonsourceibias.n506 0.189894
R23486 commonsourceibias.n508 commonsourceibias.n507 0.189894
R23487 commonsourceibias.n508 commonsourceibias.n494 0.189894
R23488 commonsourceibias.n513 commonsourceibias.n494 0.189894
R23489 commonsourceibias.n514 commonsourceibias.n513 0.189894
R23490 commonsourceibias.n514 commonsourceibias.n492 0.189894
R23491 commonsourceibias.n518 commonsourceibias.n492 0.189894
R23492 commonsourceibias.n519 commonsourceibias.n518 0.189894
R23493 commonsourceibias.n519 commonsourceibias.n490 0.189894
R23494 commonsourceibias.n523 commonsourceibias.n490 0.189894
R23495 commonsourceibias.n524 commonsourceibias.n523 0.189894
R23496 commonsourceibias.n524 commonsourceibias.n488 0.189894
R23497 commonsourceibias.n529 commonsourceibias.n488 0.189894
R23498 commonsourceibias.n530 commonsourceibias.n529 0.189894
R23499 commonsourceibias.n531 commonsourceibias.n530 0.189894
R23500 commonsourceibias.n531 commonsourceibias.n486 0.189894
R23501 commonsourceibias.n537 commonsourceibias.n486 0.189894
R23502 commonsourceibias.n538 commonsourceibias.n537 0.189894
R23503 commonsourceibias.n539 commonsourceibias.n538 0.189894
R23504 commonsourceibias.n539 commonsourceibias.n484 0.189894
R23505 commonsourceibias.n544 commonsourceibias.n484 0.189894
R23506 commonsourceibias.n545 commonsourceibias.n544 0.189894
R23507 commonsourceibias.n546 commonsourceibias.n545 0.189894
R23508 commonsourceibias.n546 commonsourceibias.n482 0.189894
R23509 commonsourceibias.n552 commonsourceibias.n482 0.189894
R23510 commonsourceibias.n553 commonsourceibias.n552 0.189894
R23511 commonsourceibias.n554 commonsourceibias.n553 0.189894
R23512 commonsourceibias.n554 commonsourceibias.n480 0.189894
R23513 commonsourceibias.n559 commonsourceibias.n480 0.189894
R23514 commonsourceibias.n560 commonsourceibias.n559 0.189894
R23515 commonsourceibias.n561 commonsourceibias.n560 0.189894
R23516 commonsourceibias.n561 commonsourceibias.n478 0.189894
R23517 commonsourceibias.n159 commonsourceibias.n158 0.170955
R23518 commonsourceibias.n160 commonsourceibias.n159 0.170955
R23519 commonsourceibias.n441 commonsourceibias.n335 0.170955
R23520 commonsourceibias.n442 commonsourceibias.n441 0.170955
R23521 diffpairibias.n0 diffpairibias.t27 436.822
R23522 diffpairibias.n27 diffpairibias.t24 435.479
R23523 diffpairibias.n26 diffpairibias.t21 435.479
R23524 diffpairibias.n25 diffpairibias.t22 435.479
R23525 diffpairibias.n24 diffpairibias.t26 435.479
R23526 diffpairibias.n23 diffpairibias.t20 435.479
R23527 diffpairibias.n0 diffpairibias.t23 435.479
R23528 diffpairibias.n1 diffpairibias.t28 435.479
R23529 diffpairibias.n2 diffpairibias.t25 435.479
R23530 diffpairibias.n3 diffpairibias.t29 435.479
R23531 diffpairibias.n13 diffpairibias.t14 377.536
R23532 diffpairibias.n13 diffpairibias.t0 376.193
R23533 diffpairibias.n14 diffpairibias.t10 376.193
R23534 diffpairibias.n15 diffpairibias.t12 376.193
R23535 diffpairibias.n16 diffpairibias.t6 376.193
R23536 diffpairibias.n17 diffpairibias.t2 376.193
R23537 diffpairibias.n18 diffpairibias.t16 376.193
R23538 diffpairibias.n19 diffpairibias.t4 376.193
R23539 diffpairibias.n20 diffpairibias.t18 376.193
R23540 diffpairibias.n21 diffpairibias.t8 376.193
R23541 diffpairibias.n4 diffpairibias.t15 113.368
R23542 diffpairibias.n4 diffpairibias.t1 112.698
R23543 diffpairibias.n5 diffpairibias.t11 112.698
R23544 diffpairibias.n6 diffpairibias.t13 112.698
R23545 diffpairibias.n7 diffpairibias.t7 112.698
R23546 diffpairibias.n8 diffpairibias.t3 112.698
R23547 diffpairibias.n9 diffpairibias.t17 112.698
R23548 diffpairibias.n10 diffpairibias.t5 112.698
R23549 diffpairibias.n11 diffpairibias.t19 112.698
R23550 diffpairibias.n12 diffpairibias.t9 112.698
R23551 diffpairibias.n22 diffpairibias.n21 4.77242
R23552 diffpairibias.n22 diffpairibias.n12 4.30807
R23553 diffpairibias.n23 diffpairibias.n22 4.13945
R23554 diffpairibias.n21 diffpairibias.n20 1.34352
R23555 diffpairibias.n20 diffpairibias.n19 1.34352
R23556 diffpairibias.n19 diffpairibias.n18 1.34352
R23557 diffpairibias.n18 diffpairibias.n17 1.34352
R23558 diffpairibias.n17 diffpairibias.n16 1.34352
R23559 diffpairibias.n16 diffpairibias.n15 1.34352
R23560 diffpairibias.n15 diffpairibias.n14 1.34352
R23561 diffpairibias.n14 diffpairibias.n13 1.34352
R23562 diffpairibias.n3 diffpairibias.n2 1.34352
R23563 diffpairibias.n2 diffpairibias.n1 1.34352
R23564 diffpairibias.n1 diffpairibias.n0 1.34352
R23565 diffpairibias.n24 diffpairibias.n23 1.34352
R23566 diffpairibias.n25 diffpairibias.n24 1.34352
R23567 diffpairibias.n26 diffpairibias.n25 1.34352
R23568 diffpairibias.n27 diffpairibias.n26 1.34352
R23569 diffpairibias.n28 diffpairibias.n27 0.862419
R23570 diffpairibias diffpairibias.n28 0.684875
R23571 diffpairibias.n12 diffpairibias.n11 0.672012
R23572 diffpairibias.n11 diffpairibias.n10 0.672012
R23573 diffpairibias.n10 diffpairibias.n9 0.672012
R23574 diffpairibias.n9 diffpairibias.n8 0.672012
R23575 diffpairibias.n8 diffpairibias.n7 0.672012
R23576 diffpairibias.n7 diffpairibias.n6 0.672012
R23577 diffpairibias.n6 diffpairibias.n5 0.672012
R23578 diffpairibias.n5 diffpairibias.n4 0.672012
R23579 diffpairibias.n28 diffpairibias.n3 0.190907
R23580 output.n41 output.n15 289.615
R23581 output.n72 output.n46 289.615
R23582 output.n104 output.n78 289.615
R23583 output.n136 output.n110 289.615
R23584 output.n77 output.n45 197.26
R23585 output.n77 output.n76 196.298
R23586 output.n109 output.n108 196.298
R23587 output.n141 output.n140 196.298
R23588 output.n42 output.n41 185
R23589 output.n40 output.n39 185
R23590 output.n19 output.n18 185
R23591 output.n34 output.n33 185
R23592 output.n32 output.n31 185
R23593 output.n23 output.n22 185
R23594 output.n26 output.n25 185
R23595 output.n73 output.n72 185
R23596 output.n71 output.n70 185
R23597 output.n50 output.n49 185
R23598 output.n65 output.n64 185
R23599 output.n63 output.n62 185
R23600 output.n54 output.n53 185
R23601 output.n57 output.n56 185
R23602 output.n105 output.n104 185
R23603 output.n103 output.n102 185
R23604 output.n82 output.n81 185
R23605 output.n97 output.n96 185
R23606 output.n95 output.n94 185
R23607 output.n86 output.n85 185
R23608 output.n89 output.n88 185
R23609 output.n137 output.n136 185
R23610 output.n135 output.n134 185
R23611 output.n114 output.n113 185
R23612 output.n129 output.n128 185
R23613 output.n127 output.n126 185
R23614 output.n118 output.n117 185
R23615 output.n121 output.n120 185
R23616 output.t19 output.n24 147.661
R23617 output.t18 output.n55 147.661
R23618 output.t1 output.n87 147.661
R23619 output.t0 output.n119 147.661
R23620 output.n41 output.n40 104.615
R23621 output.n40 output.n18 104.615
R23622 output.n33 output.n18 104.615
R23623 output.n33 output.n32 104.615
R23624 output.n32 output.n22 104.615
R23625 output.n25 output.n22 104.615
R23626 output.n72 output.n71 104.615
R23627 output.n71 output.n49 104.615
R23628 output.n64 output.n49 104.615
R23629 output.n64 output.n63 104.615
R23630 output.n63 output.n53 104.615
R23631 output.n56 output.n53 104.615
R23632 output.n104 output.n103 104.615
R23633 output.n103 output.n81 104.615
R23634 output.n96 output.n81 104.615
R23635 output.n96 output.n95 104.615
R23636 output.n95 output.n85 104.615
R23637 output.n88 output.n85 104.615
R23638 output.n136 output.n135 104.615
R23639 output.n135 output.n113 104.615
R23640 output.n128 output.n113 104.615
R23641 output.n128 output.n127 104.615
R23642 output.n127 output.n117 104.615
R23643 output.n120 output.n117 104.615
R23644 output.n1 output.t14 77.056
R23645 output.n14 output.t15 76.6694
R23646 output.n1 output.n0 72.7095
R23647 output.n3 output.n2 72.7095
R23648 output.n5 output.n4 72.7095
R23649 output.n7 output.n6 72.7095
R23650 output.n9 output.n8 72.7095
R23651 output.n11 output.n10 72.7095
R23652 output.n13 output.n12 72.7095
R23653 output.n25 output.t19 52.3082
R23654 output.n56 output.t18 52.3082
R23655 output.n88 output.t1 52.3082
R23656 output.n120 output.t0 52.3082
R23657 output.n26 output.n24 15.6674
R23658 output.n57 output.n55 15.6674
R23659 output.n89 output.n87 15.6674
R23660 output.n121 output.n119 15.6674
R23661 output.n27 output.n23 12.8005
R23662 output.n58 output.n54 12.8005
R23663 output.n90 output.n86 12.8005
R23664 output.n122 output.n118 12.8005
R23665 output.n31 output.n30 12.0247
R23666 output.n62 output.n61 12.0247
R23667 output.n94 output.n93 12.0247
R23668 output.n126 output.n125 12.0247
R23669 output.n34 output.n21 11.249
R23670 output.n65 output.n52 11.249
R23671 output.n97 output.n84 11.249
R23672 output.n129 output.n116 11.249
R23673 output.n35 output.n19 10.4732
R23674 output.n66 output.n50 10.4732
R23675 output.n98 output.n82 10.4732
R23676 output.n130 output.n114 10.4732
R23677 output.n39 output.n38 9.69747
R23678 output.n70 output.n69 9.69747
R23679 output.n102 output.n101 9.69747
R23680 output.n134 output.n133 9.69747
R23681 output.n45 output.n44 9.45567
R23682 output.n76 output.n75 9.45567
R23683 output.n108 output.n107 9.45567
R23684 output.n140 output.n139 9.45567
R23685 output.n44 output.n43 9.3005
R23686 output.n17 output.n16 9.3005
R23687 output.n38 output.n37 9.3005
R23688 output.n36 output.n35 9.3005
R23689 output.n21 output.n20 9.3005
R23690 output.n30 output.n29 9.3005
R23691 output.n28 output.n27 9.3005
R23692 output.n75 output.n74 9.3005
R23693 output.n48 output.n47 9.3005
R23694 output.n69 output.n68 9.3005
R23695 output.n67 output.n66 9.3005
R23696 output.n52 output.n51 9.3005
R23697 output.n61 output.n60 9.3005
R23698 output.n59 output.n58 9.3005
R23699 output.n107 output.n106 9.3005
R23700 output.n80 output.n79 9.3005
R23701 output.n101 output.n100 9.3005
R23702 output.n99 output.n98 9.3005
R23703 output.n84 output.n83 9.3005
R23704 output.n93 output.n92 9.3005
R23705 output.n91 output.n90 9.3005
R23706 output.n139 output.n138 9.3005
R23707 output.n112 output.n111 9.3005
R23708 output.n133 output.n132 9.3005
R23709 output.n131 output.n130 9.3005
R23710 output.n116 output.n115 9.3005
R23711 output.n125 output.n124 9.3005
R23712 output.n123 output.n122 9.3005
R23713 output.n42 output.n17 8.92171
R23714 output.n73 output.n48 8.92171
R23715 output.n105 output.n80 8.92171
R23716 output.n137 output.n112 8.92171
R23717 output output.n141 8.15037
R23718 output.n43 output.n15 8.14595
R23719 output.n74 output.n46 8.14595
R23720 output.n106 output.n78 8.14595
R23721 output.n138 output.n110 8.14595
R23722 output.n45 output.n15 5.81868
R23723 output.n76 output.n46 5.81868
R23724 output.n108 output.n78 5.81868
R23725 output.n140 output.n110 5.81868
R23726 output.n43 output.n42 5.04292
R23727 output.n74 output.n73 5.04292
R23728 output.n106 output.n105 5.04292
R23729 output.n138 output.n137 5.04292
R23730 output.n28 output.n24 4.38594
R23731 output.n59 output.n55 4.38594
R23732 output.n91 output.n87 4.38594
R23733 output.n123 output.n119 4.38594
R23734 output.n39 output.n17 4.26717
R23735 output.n70 output.n48 4.26717
R23736 output.n102 output.n80 4.26717
R23737 output.n134 output.n112 4.26717
R23738 output.n0 output.t4 3.9605
R23739 output.n0 output.t8 3.9605
R23740 output.n2 output.t11 3.9605
R23741 output.n2 output.t16 3.9605
R23742 output.n4 output.t17 3.9605
R23743 output.n4 output.t6 3.9605
R23744 output.n6 output.t10 3.9605
R23745 output.n6 output.t2 3.9605
R23746 output.n8 output.t5 3.9605
R23747 output.n8 output.t3 3.9605
R23748 output.n10 output.t9 3.9605
R23749 output.n10 output.t12 3.9605
R23750 output.n12 output.t13 3.9605
R23751 output.n12 output.t7 3.9605
R23752 output.n38 output.n19 3.49141
R23753 output.n69 output.n50 3.49141
R23754 output.n101 output.n82 3.49141
R23755 output.n133 output.n114 3.49141
R23756 output.n35 output.n34 2.71565
R23757 output.n66 output.n65 2.71565
R23758 output.n98 output.n97 2.71565
R23759 output.n130 output.n129 2.71565
R23760 output.n31 output.n21 1.93989
R23761 output.n62 output.n52 1.93989
R23762 output.n94 output.n84 1.93989
R23763 output.n126 output.n116 1.93989
R23764 output.n30 output.n23 1.16414
R23765 output.n61 output.n54 1.16414
R23766 output.n93 output.n86 1.16414
R23767 output.n125 output.n118 1.16414
R23768 output.n141 output.n109 0.962709
R23769 output.n109 output.n77 0.962709
R23770 output.n27 output.n26 0.388379
R23771 output.n58 output.n57 0.388379
R23772 output.n90 output.n89 0.388379
R23773 output.n122 output.n121 0.388379
R23774 output.n14 output.n13 0.387128
R23775 output.n13 output.n11 0.387128
R23776 output.n11 output.n9 0.387128
R23777 output.n9 output.n7 0.387128
R23778 output.n7 output.n5 0.387128
R23779 output.n5 output.n3 0.387128
R23780 output.n3 output.n1 0.387128
R23781 output.n44 output.n16 0.155672
R23782 output.n37 output.n16 0.155672
R23783 output.n37 output.n36 0.155672
R23784 output.n36 output.n20 0.155672
R23785 output.n29 output.n20 0.155672
R23786 output.n29 output.n28 0.155672
R23787 output.n75 output.n47 0.155672
R23788 output.n68 output.n47 0.155672
R23789 output.n68 output.n67 0.155672
R23790 output.n67 output.n51 0.155672
R23791 output.n60 output.n51 0.155672
R23792 output.n60 output.n59 0.155672
R23793 output.n107 output.n79 0.155672
R23794 output.n100 output.n79 0.155672
R23795 output.n100 output.n99 0.155672
R23796 output.n99 output.n83 0.155672
R23797 output.n92 output.n83 0.155672
R23798 output.n92 output.n91 0.155672
R23799 output.n139 output.n111 0.155672
R23800 output.n132 output.n111 0.155672
R23801 output.n132 output.n131 0.155672
R23802 output.n131 output.n115 0.155672
R23803 output.n124 output.n115 0.155672
R23804 output.n124 output.n123 0.155672
R23805 output output.n14 0.126227
R23806 a_n2650_8322.n10 a_n2650_8322.t3 74.6477
R23807 a_n2650_8322.n1 a_n2650_8322.t23 74.6477
R23808 a_n2650_8322.n24 a_n2650_8322.t25 74.6474
R23809 a_n2650_8322.n18 a_n2650_8322.t22 74.2899
R23810 a_n2650_8322.n11 a_n2650_8322.t1 74.2899
R23811 a_n2650_8322.n12 a_n2650_8322.t4 74.2899
R23812 a_n2650_8322.n15 a_n2650_8322.t5 74.2899
R23813 a_n2650_8322.n8 a_n2650_8322.t8 74.2899
R23814 a_n2650_8322.n24 a_n2650_8322.n23 70.6783
R23815 a_n2650_8322.n22 a_n2650_8322.n21 70.6783
R23816 a_n2650_8322.n20 a_n2650_8322.n19 70.6783
R23817 a_n2650_8322.n10 a_n2650_8322.n9 70.6783
R23818 a_n2650_8322.n14 a_n2650_8322.n13 70.6783
R23819 a_n2650_8322.n1 a_n2650_8322.n0 70.6783
R23820 a_n2650_8322.n3 a_n2650_8322.n2 70.6783
R23821 a_n2650_8322.n5 a_n2650_8322.n4 70.6783
R23822 a_n2650_8322.n7 a_n2650_8322.n6 70.6783
R23823 a_n2650_8322.n26 a_n2650_8322.n25 70.6782
R23824 a_n2650_8322.n16 a_n2650_8322.n8 24.1867
R23825 a_n2650_8322.n17 a_n2650_8322.t28 9.90091
R23826 a_n2650_8322.n16 a_n2650_8322.n15 7.67184
R23827 a_n2650_8322.n18 a_n2650_8322.n17 6.55222
R23828 a_n2650_8322.n17 a_n2650_8322.n16 5.3452
R23829 a_n2650_8322.n23 a_n2650_8322.t20 3.61217
R23830 a_n2650_8322.n23 a_n2650_8322.t16 3.61217
R23831 a_n2650_8322.n21 a_n2650_8322.t24 3.61217
R23832 a_n2650_8322.n21 a_n2650_8322.t14 3.61217
R23833 a_n2650_8322.n19 a_n2650_8322.t12 3.61217
R23834 a_n2650_8322.n19 a_n2650_8322.t11 3.61217
R23835 a_n2650_8322.n9 a_n2650_8322.t7 3.61217
R23836 a_n2650_8322.n9 a_n2650_8322.t6 3.61217
R23837 a_n2650_8322.n13 a_n2650_8322.t2 3.61217
R23838 a_n2650_8322.n13 a_n2650_8322.t0 3.61217
R23839 a_n2650_8322.n0 a_n2650_8322.t26 3.61217
R23840 a_n2650_8322.n0 a_n2650_8322.t18 3.61217
R23841 a_n2650_8322.n2 a_n2650_8322.t10 3.61217
R23842 a_n2650_8322.n2 a_n2650_8322.t9 3.61217
R23843 a_n2650_8322.n4 a_n2650_8322.t21 3.61217
R23844 a_n2650_8322.n4 a_n2650_8322.t15 3.61217
R23845 a_n2650_8322.n6 a_n2650_8322.t19 3.61217
R23846 a_n2650_8322.n6 a_n2650_8322.t17 3.61217
R23847 a_n2650_8322.n26 a_n2650_8322.t13 3.61217
R23848 a_n2650_8322.t27 a_n2650_8322.n26 3.61217
R23849 a_n2650_8322.n15 a_n2650_8322.n14 0.358259
R23850 a_n2650_8322.n14 a_n2650_8322.n12 0.358259
R23851 a_n2650_8322.n11 a_n2650_8322.n10 0.358259
R23852 a_n2650_8322.n8 a_n2650_8322.n7 0.358259
R23853 a_n2650_8322.n7 a_n2650_8322.n5 0.358259
R23854 a_n2650_8322.n5 a_n2650_8322.n3 0.358259
R23855 a_n2650_8322.n3 a_n2650_8322.n1 0.358259
R23856 a_n2650_8322.n20 a_n2650_8322.n18 0.358259
R23857 a_n2650_8322.n22 a_n2650_8322.n20 0.358259
R23858 a_n2650_8322.n25 a_n2650_8322.n22 0.358259
R23859 a_n2650_8322.n25 a_n2650_8322.n24 0.358259
R23860 a_n2650_8322.n12 a_n2650_8322.n11 0.101793
R23861 a_n2650_8322.t30 a_n2650_8322.t33 0.0788333
R23862 a_n2650_8322.t29 a_n2650_8322.t31 0.0788333
R23863 a_n2650_8322.t28 a_n2650_8322.t32 0.0788333
R23864 a_n2650_8322.t29 a_n2650_8322.t30 0.0318333
R23865 a_n2650_8322.t28 a_n2650_8322.t31 0.0318333
R23866 a_n2650_8322.t33 a_n2650_8322.t31 0.0318333
R23867 a_n2650_8322.t32 a_n2650_8322.t29 0.0318333
R23868 minus.n61 minus.t24 251.488
R23869 minus.n12 minus.t16 251.488
R23870 minus.n102 minus.t4 243.255
R23871 minus.n96 minus.t14 231.093
R23872 minus.n47 minus.t9 231.093
R23873 minus.n101 minus.n99 224.169
R23874 minus.n101 minus.n100 223.454
R23875 minus.n50 minus.t21 187.445
R23876 minus.n89 minus.t18 187.445
R23877 minus.n83 minus.t15 187.445
R23878 minus.n54 minus.t7 187.445
R23879 minus.n56 minus.t6 187.445
R23880 minus.n71 minus.t12 187.445
R23881 minus.n65 minus.t11 187.445
R23882 minus.n60 minus.t19 187.445
R23883 minus.n11 minus.t10 187.445
R23884 minus.n16 minus.t8 187.445
R23885 minus.n22 minus.t5 187.445
R23886 minus.n7 minus.t22 187.445
R23887 minus.n5 minus.t23 187.445
R23888 minus.n34 minus.t17 187.445
R23889 minus.n40 minus.t20 187.445
R23890 minus.n1 minus.t13 187.445
R23891 minus.n63 minus.n62 161.3
R23892 minus.n64 minus.n59 161.3
R23893 minus.n67 minus.n66 161.3
R23894 minus.n68 minus.n58 161.3
R23895 minus.n70 minus.n69 161.3
R23896 minus.n72 minus.n57 161.3
R23897 minus.n74 minus.n73 161.3
R23898 minus.n76 minus.n75 161.3
R23899 minus.n77 minus.n55 161.3
R23900 minus.n79 minus.n78 161.3
R23901 minus.n81 minus.n80 161.3
R23902 minus.n82 minus.n53 161.3
R23903 minus.n85 minus.n84 161.3
R23904 minus.n86 minus.n52 161.3
R23905 minus.n88 minus.n87 161.3
R23906 minus.n90 minus.n51 161.3
R23907 minus.n92 minus.n91 161.3
R23908 minus.n94 minus.n93 161.3
R23909 minus.n95 minus.n49 161.3
R23910 minus.n97 minus.n96 161.3
R23911 minus.n48 minus.n47 161.3
R23912 minus.n46 minus.n0 161.3
R23913 minus.n45 minus.n44 161.3
R23914 minus.n43 minus.n42 161.3
R23915 minus.n41 minus.n2 161.3
R23916 minus.n39 minus.n38 161.3
R23917 minus.n37 minus.n3 161.3
R23918 minus.n36 minus.n35 161.3
R23919 minus.n33 minus.n4 161.3
R23920 minus.n32 minus.n31 161.3
R23921 minus.n30 minus.n29 161.3
R23922 minus.n28 minus.n6 161.3
R23923 minus.n27 minus.n26 161.3
R23924 minus.n25 minus.n24 161.3
R23925 minus.n23 minus.n8 161.3
R23926 minus.n21 minus.n20 161.3
R23927 minus.n19 minus.n9 161.3
R23928 minus.n18 minus.n17 161.3
R23929 minus.n15 minus.n10 161.3
R23930 minus.n14 minus.n13 161.3
R23931 minus.n91 minus.n90 56.5617
R23932 minus.n64 minus.n63 56.5617
R23933 minus.n15 minus.n14 56.5617
R23934 minus.n42 minus.n41 56.5617
R23935 minus.n82 minus.n81 56.5617
R23936 minus.n73 minus.n72 56.5617
R23937 minus.n24 minus.n23 56.5617
R23938 minus.n33 minus.n32 56.5617
R23939 minus.n95 minus.n94 48.3272
R23940 minus.n46 minus.n45 48.3272
R23941 minus.n84 minus.n52 44.4521
R23942 minus.n70 minus.n58 44.4521
R23943 minus.n21 minus.n9 44.4521
R23944 minus.n35 minus.n3 44.4521
R23945 minus.n13 minus.n12 43.0014
R23946 minus.n62 minus.n61 43.0014
R23947 minus.n78 minus.n77 40.577
R23948 minus.n77 minus.n76 40.577
R23949 minus.n28 minus.n27 40.577
R23950 minus.n29 minus.n28 40.577
R23951 minus.n61 minus.n60 39.4345
R23952 minus.n12 minus.n11 39.4345
R23953 minus.n88 minus.n52 36.702
R23954 minus.n66 minus.n58 36.702
R23955 minus.n17 minus.n9 36.702
R23956 minus.n39 minus.n3 36.702
R23957 minus.n98 minus.n97 33.563
R23958 minus.n90 minus.n89 20.9036
R23959 minus.n65 minus.n64 20.9036
R23960 minus.n16 minus.n15 20.9036
R23961 minus.n41 minus.n40 20.9036
R23962 minus.n100 minus.t3 19.8005
R23963 minus.n100 minus.t0 19.8005
R23964 minus.n99 minus.t2 19.8005
R23965 minus.n99 minus.t1 19.8005
R23966 minus.n81 minus.n54 18.9362
R23967 minus.n73 minus.n56 18.9362
R23968 minus.n24 minus.n7 18.9362
R23969 minus.n32 minus.n5 18.9362
R23970 minus.n83 minus.n82 16.9689
R23971 minus.n72 minus.n71 16.9689
R23972 minus.n23 minus.n22 16.9689
R23973 minus.n34 minus.n33 16.9689
R23974 minus.n91 minus.n50 15.0015
R23975 minus.n63 minus.n60 15.0015
R23976 minus.n14 minus.n11 15.0015
R23977 minus.n42 minus.n1 15.0015
R23978 minus.n96 minus.n95 12.4157
R23979 minus.n47 minus.n46 12.4157
R23980 minus.n98 minus.n48 12.1577
R23981 minus minus.n103 11.6918
R23982 minus.n94 minus.n50 9.59132
R23983 minus.n45 minus.n1 9.59132
R23984 minus.n84 minus.n83 7.62397
R23985 minus.n71 minus.n70 7.62397
R23986 minus.n22 minus.n21 7.62397
R23987 minus.n35 minus.n34 7.62397
R23988 minus.n78 minus.n54 5.65662
R23989 minus.n76 minus.n56 5.65662
R23990 minus.n27 minus.n7 5.65662
R23991 minus.n29 minus.n5 5.65662
R23992 minus.n103 minus.n102 4.80222
R23993 minus.n89 minus.n88 3.68928
R23994 minus.n66 minus.n65 3.68928
R23995 minus.n17 minus.n16 3.68928
R23996 minus.n40 minus.n39 3.68928
R23997 minus.n103 minus.n98 0.972091
R23998 minus.n102 minus.n101 0.716017
R23999 minus.n97 minus.n49 0.189894
R24000 minus.n93 minus.n49 0.189894
R24001 minus.n93 minus.n92 0.189894
R24002 minus.n92 minus.n51 0.189894
R24003 minus.n87 minus.n51 0.189894
R24004 minus.n87 minus.n86 0.189894
R24005 minus.n86 minus.n85 0.189894
R24006 minus.n85 minus.n53 0.189894
R24007 minus.n80 minus.n53 0.189894
R24008 minus.n80 minus.n79 0.189894
R24009 minus.n79 minus.n55 0.189894
R24010 minus.n75 minus.n55 0.189894
R24011 minus.n75 minus.n74 0.189894
R24012 minus.n74 minus.n57 0.189894
R24013 minus.n69 minus.n57 0.189894
R24014 minus.n69 minus.n68 0.189894
R24015 minus.n68 minus.n67 0.189894
R24016 minus.n67 minus.n59 0.189894
R24017 minus.n62 minus.n59 0.189894
R24018 minus.n13 minus.n10 0.189894
R24019 minus.n18 minus.n10 0.189894
R24020 minus.n19 minus.n18 0.189894
R24021 minus.n20 minus.n19 0.189894
R24022 minus.n20 minus.n8 0.189894
R24023 minus.n25 minus.n8 0.189894
R24024 minus.n26 minus.n25 0.189894
R24025 minus.n26 minus.n6 0.189894
R24026 minus.n30 minus.n6 0.189894
R24027 minus.n31 minus.n30 0.189894
R24028 minus.n31 minus.n4 0.189894
R24029 minus.n36 minus.n4 0.189894
R24030 minus.n37 minus.n36 0.189894
R24031 minus.n38 minus.n37 0.189894
R24032 minus.n38 minus.n2 0.189894
R24033 minus.n43 minus.n2 0.189894
R24034 minus.n44 minus.n43 0.189894
R24035 minus.n44 minus.n0 0.189894
R24036 minus.n48 minus.n0 0.189894
R24037 outputibias.n27 outputibias.n1 289.615
R24038 outputibias.n58 outputibias.n32 289.615
R24039 outputibias.n90 outputibias.n64 289.615
R24040 outputibias.n122 outputibias.n96 289.615
R24041 outputibias.n28 outputibias.n27 185
R24042 outputibias.n26 outputibias.n25 185
R24043 outputibias.n5 outputibias.n4 185
R24044 outputibias.n20 outputibias.n19 185
R24045 outputibias.n18 outputibias.n17 185
R24046 outputibias.n9 outputibias.n8 185
R24047 outputibias.n12 outputibias.n11 185
R24048 outputibias.n59 outputibias.n58 185
R24049 outputibias.n57 outputibias.n56 185
R24050 outputibias.n36 outputibias.n35 185
R24051 outputibias.n51 outputibias.n50 185
R24052 outputibias.n49 outputibias.n48 185
R24053 outputibias.n40 outputibias.n39 185
R24054 outputibias.n43 outputibias.n42 185
R24055 outputibias.n91 outputibias.n90 185
R24056 outputibias.n89 outputibias.n88 185
R24057 outputibias.n68 outputibias.n67 185
R24058 outputibias.n83 outputibias.n82 185
R24059 outputibias.n81 outputibias.n80 185
R24060 outputibias.n72 outputibias.n71 185
R24061 outputibias.n75 outputibias.n74 185
R24062 outputibias.n123 outputibias.n122 185
R24063 outputibias.n121 outputibias.n120 185
R24064 outputibias.n100 outputibias.n99 185
R24065 outputibias.n115 outputibias.n114 185
R24066 outputibias.n113 outputibias.n112 185
R24067 outputibias.n104 outputibias.n103 185
R24068 outputibias.n107 outputibias.n106 185
R24069 outputibias.n0 outputibias.t8 178.945
R24070 outputibias.n133 outputibias.t11 177.018
R24071 outputibias.n132 outputibias.t9 177.018
R24072 outputibias.n0 outputibias.t10 177.018
R24073 outputibias.t5 outputibias.n10 147.661
R24074 outputibias.t7 outputibias.n41 147.661
R24075 outputibias.t1 outputibias.n73 147.661
R24076 outputibias.t3 outputibias.n105 147.661
R24077 outputibias.n128 outputibias.t4 132.363
R24078 outputibias.n128 outputibias.t6 130.436
R24079 outputibias.n129 outputibias.t0 130.436
R24080 outputibias.n130 outputibias.t2 130.436
R24081 outputibias.n27 outputibias.n26 104.615
R24082 outputibias.n26 outputibias.n4 104.615
R24083 outputibias.n19 outputibias.n4 104.615
R24084 outputibias.n19 outputibias.n18 104.615
R24085 outputibias.n18 outputibias.n8 104.615
R24086 outputibias.n11 outputibias.n8 104.615
R24087 outputibias.n58 outputibias.n57 104.615
R24088 outputibias.n57 outputibias.n35 104.615
R24089 outputibias.n50 outputibias.n35 104.615
R24090 outputibias.n50 outputibias.n49 104.615
R24091 outputibias.n49 outputibias.n39 104.615
R24092 outputibias.n42 outputibias.n39 104.615
R24093 outputibias.n90 outputibias.n89 104.615
R24094 outputibias.n89 outputibias.n67 104.615
R24095 outputibias.n82 outputibias.n67 104.615
R24096 outputibias.n82 outputibias.n81 104.615
R24097 outputibias.n81 outputibias.n71 104.615
R24098 outputibias.n74 outputibias.n71 104.615
R24099 outputibias.n122 outputibias.n121 104.615
R24100 outputibias.n121 outputibias.n99 104.615
R24101 outputibias.n114 outputibias.n99 104.615
R24102 outputibias.n114 outputibias.n113 104.615
R24103 outputibias.n113 outputibias.n103 104.615
R24104 outputibias.n106 outputibias.n103 104.615
R24105 outputibias.n63 outputibias.n31 95.6354
R24106 outputibias.n63 outputibias.n62 94.6732
R24107 outputibias.n95 outputibias.n94 94.6732
R24108 outputibias.n127 outputibias.n126 94.6732
R24109 outputibias.n11 outputibias.t5 52.3082
R24110 outputibias.n42 outputibias.t7 52.3082
R24111 outputibias.n74 outputibias.t1 52.3082
R24112 outputibias.n106 outputibias.t3 52.3082
R24113 outputibias.n12 outputibias.n10 15.6674
R24114 outputibias.n43 outputibias.n41 15.6674
R24115 outputibias.n75 outputibias.n73 15.6674
R24116 outputibias.n107 outputibias.n105 15.6674
R24117 outputibias.n13 outputibias.n9 12.8005
R24118 outputibias.n44 outputibias.n40 12.8005
R24119 outputibias.n76 outputibias.n72 12.8005
R24120 outputibias.n108 outputibias.n104 12.8005
R24121 outputibias.n17 outputibias.n16 12.0247
R24122 outputibias.n48 outputibias.n47 12.0247
R24123 outputibias.n80 outputibias.n79 12.0247
R24124 outputibias.n112 outputibias.n111 12.0247
R24125 outputibias.n20 outputibias.n7 11.249
R24126 outputibias.n51 outputibias.n38 11.249
R24127 outputibias.n83 outputibias.n70 11.249
R24128 outputibias.n115 outputibias.n102 11.249
R24129 outputibias.n21 outputibias.n5 10.4732
R24130 outputibias.n52 outputibias.n36 10.4732
R24131 outputibias.n84 outputibias.n68 10.4732
R24132 outputibias.n116 outputibias.n100 10.4732
R24133 outputibias.n25 outputibias.n24 9.69747
R24134 outputibias.n56 outputibias.n55 9.69747
R24135 outputibias.n88 outputibias.n87 9.69747
R24136 outputibias.n120 outputibias.n119 9.69747
R24137 outputibias.n31 outputibias.n30 9.45567
R24138 outputibias.n62 outputibias.n61 9.45567
R24139 outputibias.n94 outputibias.n93 9.45567
R24140 outputibias.n126 outputibias.n125 9.45567
R24141 outputibias.n30 outputibias.n29 9.3005
R24142 outputibias.n3 outputibias.n2 9.3005
R24143 outputibias.n24 outputibias.n23 9.3005
R24144 outputibias.n22 outputibias.n21 9.3005
R24145 outputibias.n7 outputibias.n6 9.3005
R24146 outputibias.n16 outputibias.n15 9.3005
R24147 outputibias.n14 outputibias.n13 9.3005
R24148 outputibias.n61 outputibias.n60 9.3005
R24149 outputibias.n34 outputibias.n33 9.3005
R24150 outputibias.n55 outputibias.n54 9.3005
R24151 outputibias.n53 outputibias.n52 9.3005
R24152 outputibias.n38 outputibias.n37 9.3005
R24153 outputibias.n47 outputibias.n46 9.3005
R24154 outputibias.n45 outputibias.n44 9.3005
R24155 outputibias.n93 outputibias.n92 9.3005
R24156 outputibias.n66 outputibias.n65 9.3005
R24157 outputibias.n87 outputibias.n86 9.3005
R24158 outputibias.n85 outputibias.n84 9.3005
R24159 outputibias.n70 outputibias.n69 9.3005
R24160 outputibias.n79 outputibias.n78 9.3005
R24161 outputibias.n77 outputibias.n76 9.3005
R24162 outputibias.n125 outputibias.n124 9.3005
R24163 outputibias.n98 outputibias.n97 9.3005
R24164 outputibias.n119 outputibias.n118 9.3005
R24165 outputibias.n117 outputibias.n116 9.3005
R24166 outputibias.n102 outputibias.n101 9.3005
R24167 outputibias.n111 outputibias.n110 9.3005
R24168 outputibias.n109 outputibias.n108 9.3005
R24169 outputibias.n28 outputibias.n3 8.92171
R24170 outputibias.n59 outputibias.n34 8.92171
R24171 outputibias.n91 outputibias.n66 8.92171
R24172 outputibias.n123 outputibias.n98 8.92171
R24173 outputibias.n29 outputibias.n1 8.14595
R24174 outputibias.n60 outputibias.n32 8.14595
R24175 outputibias.n92 outputibias.n64 8.14595
R24176 outputibias.n124 outputibias.n96 8.14595
R24177 outputibias.n31 outputibias.n1 5.81868
R24178 outputibias.n62 outputibias.n32 5.81868
R24179 outputibias.n94 outputibias.n64 5.81868
R24180 outputibias.n126 outputibias.n96 5.81868
R24181 outputibias.n131 outputibias.n130 5.20947
R24182 outputibias.n29 outputibias.n28 5.04292
R24183 outputibias.n60 outputibias.n59 5.04292
R24184 outputibias.n92 outputibias.n91 5.04292
R24185 outputibias.n124 outputibias.n123 5.04292
R24186 outputibias.n131 outputibias.n127 4.42209
R24187 outputibias.n14 outputibias.n10 4.38594
R24188 outputibias.n45 outputibias.n41 4.38594
R24189 outputibias.n77 outputibias.n73 4.38594
R24190 outputibias.n109 outputibias.n105 4.38594
R24191 outputibias.n132 outputibias.n131 4.28454
R24192 outputibias.n25 outputibias.n3 4.26717
R24193 outputibias.n56 outputibias.n34 4.26717
R24194 outputibias.n88 outputibias.n66 4.26717
R24195 outputibias.n120 outputibias.n98 4.26717
R24196 outputibias.n24 outputibias.n5 3.49141
R24197 outputibias.n55 outputibias.n36 3.49141
R24198 outputibias.n87 outputibias.n68 3.49141
R24199 outputibias.n119 outputibias.n100 3.49141
R24200 outputibias.n21 outputibias.n20 2.71565
R24201 outputibias.n52 outputibias.n51 2.71565
R24202 outputibias.n84 outputibias.n83 2.71565
R24203 outputibias.n116 outputibias.n115 2.71565
R24204 outputibias.n17 outputibias.n7 1.93989
R24205 outputibias.n48 outputibias.n38 1.93989
R24206 outputibias.n80 outputibias.n70 1.93989
R24207 outputibias.n112 outputibias.n102 1.93989
R24208 outputibias.n130 outputibias.n129 1.9266
R24209 outputibias.n129 outputibias.n128 1.9266
R24210 outputibias.n133 outputibias.n132 1.92658
R24211 outputibias.n134 outputibias.n133 1.29913
R24212 outputibias.n16 outputibias.n9 1.16414
R24213 outputibias.n47 outputibias.n40 1.16414
R24214 outputibias.n79 outputibias.n72 1.16414
R24215 outputibias.n111 outputibias.n104 1.16414
R24216 outputibias.n127 outputibias.n95 0.962709
R24217 outputibias.n95 outputibias.n63 0.962709
R24218 outputibias.n13 outputibias.n12 0.388379
R24219 outputibias.n44 outputibias.n43 0.388379
R24220 outputibias.n76 outputibias.n75 0.388379
R24221 outputibias.n108 outputibias.n107 0.388379
R24222 outputibias.n134 outputibias.n0 0.337251
R24223 outputibias outputibias.n134 0.302375
R24224 outputibias.n30 outputibias.n2 0.155672
R24225 outputibias.n23 outputibias.n2 0.155672
R24226 outputibias.n23 outputibias.n22 0.155672
R24227 outputibias.n22 outputibias.n6 0.155672
R24228 outputibias.n15 outputibias.n6 0.155672
R24229 outputibias.n15 outputibias.n14 0.155672
R24230 outputibias.n61 outputibias.n33 0.155672
R24231 outputibias.n54 outputibias.n33 0.155672
R24232 outputibias.n54 outputibias.n53 0.155672
R24233 outputibias.n53 outputibias.n37 0.155672
R24234 outputibias.n46 outputibias.n37 0.155672
R24235 outputibias.n46 outputibias.n45 0.155672
R24236 outputibias.n93 outputibias.n65 0.155672
R24237 outputibias.n86 outputibias.n65 0.155672
R24238 outputibias.n86 outputibias.n85 0.155672
R24239 outputibias.n85 outputibias.n69 0.155672
R24240 outputibias.n78 outputibias.n69 0.155672
R24241 outputibias.n78 outputibias.n77 0.155672
R24242 outputibias.n125 outputibias.n97 0.155672
R24243 outputibias.n118 outputibias.n97 0.155672
R24244 outputibias.n118 outputibias.n117 0.155672
R24245 outputibias.n117 outputibias.n101 0.155672
R24246 outputibias.n110 outputibias.n101 0.155672
R24247 outputibias.n110 outputibias.n109 0.155672
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.141215p
C5 commonsourceibias output 0.006808f
C6 minus diffpairibias 5.12e-19
C7 CSoutput minus 2.88948f
C8 vdd plus 0.099732f
C9 plus diffpairibias 4.13e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.893164f
C13 commonsourceibias diffpairibias 0.052527f
C14 CSoutput commonsourceibias 37.4715f
C15 minus plus 9.943621f
C16 minus commonsourceibias 0.337885f
C17 plus commonsourceibias 0.284038f
C18 diffpairibias gnd 59.99123f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.150736p
C22 plus gnd 36.4707f
C23 minus gnd 29.65454f
C24 CSoutput gnd 0.102137p
C25 vdd gnd 0.508888p
C26 outputibias.t10 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t5 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t7 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t1 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t3 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t2 gnd 0.108319f
C161 outputibias.t0 gnd 0.108319f
C162 outputibias.t6 gnd 0.108319f
C163 outputibias.t4 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t9 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t11 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 minus.n0 gnd 0.030108f
C174 minus.t13 gnd 0.506264f
C175 minus.n1 gnd 0.204756f
C176 minus.n2 gnd 0.030108f
C177 minus.t20 gnd 0.506264f
C178 minus.n3 gnd 0.024937f
C179 minus.n4 gnd 0.030108f
C180 minus.t17 gnd 0.506264f
C181 minus.t23 gnd 0.506264f
C182 minus.n5 gnd 0.204756f
C183 minus.n6 gnd 0.030108f
C184 minus.t22 gnd 0.506264f
C185 minus.n7 gnd 0.204756f
C186 minus.n8 gnd 0.030108f
C187 minus.t5 gnd 0.506264f
C188 minus.n9 gnd 0.024937f
C189 minus.n10 gnd 0.030108f
C190 minus.t8 gnd 0.506264f
C191 minus.t10 gnd 0.506264f
C192 minus.n11 gnd 0.235461f
C193 minus.t16 gnd 0.567388f
C194 minus.n12 gnd 0.238474f
C195 minus.n13 gnd 0.128509f
C196 minus.n14 gnd 0.038015f
C197 minus.n15 gnd 0.034634f
C198 minus.n16 gnd 0.204756f
C199 minus.n17 gnd 0.036951f
C200 minus.n18 gnd 0.030108f
C201 minus.n19 gnd 0.030108f
C202 minus.n20 gnd 0.030108f
C203 minus.n21 gnd 0.039031f
C204 minus.n22 gnd 0.204756f
C205 minus.n23 gnd 0.036888f
C206 minus.n24 gnd 0.035761f
C207 minus.n25 gnd 0.030108f
C208 minus.n26 gnd 0.030108f
C209 minus.n27 gnd 0.038301f
C210 minus.n28 gnd 0.024317f
C211 minus.n29 gnd 0.038301f
C212 minus.n30 gnd 0.030108f
C213 minus.n31 gnd 0.030108f
C214 minus.n32 gnd 0.035761f
C215 minus.n33 gnd 0.036888f
C216 minus.n34 gnd 0.204756f
C217 minus.n35 gnd 0.039031f
C218 minus.n36 gnd 0.030108f
C219 minus.n37 gnd 0.030108f
C220 minus.n38 gnd 0.030108f
C221 minus.n39 gnd 0.036951f
C222 minus.n40 gnd 0.204756f
C223 minus.n41 gnd 0.034634f
C224 minus.n42 gnd 0.038015f
C225 minus.n43 gnd 0.030108f
C226 minus.n44 gnd 0.030108f
C227 minus.n45 gnd 0.03929f
C228 minus.n46 gnd 0.011661f
C229 minus.t9 gnd 0.547525f
C230 minus.n47 gnd 0.237444f
C231 minus.n48 gnd 0.353241f
C232 minus.n49 gnd 0.030108f
C233 minus.t14 gnd 0.547525f
C234 minus.t21 gnd 0.506264f
C235 minus.n50 gnd 0.204756f
C236 minus.n51 gnd 0.030108f
C237 minus.t18 gnd 0.506264f
C238 minus.n52 gnd 0.024937f
C239 minus.n53 gnd 0.030108f
C240 minus.t15 gnd 0.506264f
C241 minus.t7 gnd 0.506264f
C242 minus.n54 gnd 0.204756f
C243 minus.n55 gnd 0.030108f
C244 minus.t6 gnd 0.506264f
C245 minus.n56 gnd 0.204756f
C246 minus.n57 gnd 0.030108f
C247 minus.t12 gnd 0.506264f
C248 minus.n58 gnd 0.024937f
C249 minus.n59 gnd 0.030108f
C250 minus.t11 gnd 0.506264f
C251 minus.t19 gnd 0.506264f
C252 minus.n60 gnd 0.235461f
C253 minus.t24 gnd 0.567388f
C254 minus.n61 gnd 0.238474f
C255 minus.n62 gnd 0.128509f
C256 minus.n63 gnd 0.038015f
C257 minus.n64 gnd 0.034634f
C258 minus.n65 gnd 0.204756f
C259 minus.n66 gnd 0.036951f
C260 minus.n67 gnd 0.030108f
C261 minus.n68 gnd 0.030108f
C262 minus.n69 gnd 0.030108f
C263 minus.n70 gnd 0.039031f
C264 minus.n71 gnd 0.204756f
C265 minus.n72 gnd 0.036888f
C266 minus.n73 gnd 0.035761f
C267 minus.n74 gnd 0.030108f
C268 minus.n75 gnd 0.030108f
C269 minus.n76 gnd 0.038301f
C270 minus.n77 gnd 0.024317f
C271 minus.n78 gnd 0.038301f
C272 minus.n79 gnd 0.030108f
C273 minus.n80 gnd 0.030108f
C274 minus.n81 gnd 0.035761f
C275 minus.n82 gnd 0.036888f
C276 minus.n83 gnd 0.204756f
C277 minus.n84 gnd 0.039031f
C278 minus.n85 gnd 0.030108f
C279 minus.n86 gnd 0.030108f
C280 minus.n87 gnd 0.030108f
C281 minus.n88 gnd 0.036951f
C282 minus.n89 gnd 0.204756f
C283 minus.n90 gnd 0.034634f
C284 minus.n91 gnd 0.038015f
C285 minus.n92 gnd 0.030108f
C286 minus.n93 gnd 0.030108f
C287 minus.n94 gnd 0.03929f
C288 minus.n95 gnd 0.011661f
C289 minus.n96 gnd 0.237444f
C290 minus.n97 gnd 1.01764f
C291 minus.n98 gnd 1.51235f
C292 minus.t2 gnd 0.009282f
C293 minus.t1 gnd 0.009282f
C294 minus.n99 gnd 0.03052f
C295 minus.t3 gnd 0.009282f
C296 minus.t0 gnd 0.009282f
C297 minus.n100 gnd 0.030101f
C298 minus.n101 gnd 0.256902f
C299 minus.t4 gnd 0.05166f
C300 minus.n102 gnd 0.140189f
C301 minus.n103 gnd 1.99138f
C302 a_n2650_8322.t13 gnd 0.097992f
C303 a_n2650_8322.t31 gnd 20.329401f
C304 a_n2650_8322.t33 gnd 20.186901f
C305 a_n2650_8322.t30 gnd 20.186901f
C306 a_n2650_8322.t29 gnd 20.329401f
C307 a_n2650_8322.t32 gnd 20.186901f
C308 a_n2650_8322.t28 gnd 29.294302f
C309 a_n2650_8322.t23 gnd 0.917551f
C310 a_n2650_8322.t26 gnd 0.097992f
C311 a_n2650_8322.t18 gnd 0.097992f
C312 a_n2650_8322.n0 gnd 0.690258f
C313 a_n2650_8322.n1 gnd 0.771262f
C314 a_n2650_8322.t10 gnd 0.097992f
C315 a_n2650_8322.t9 gnd 0.097992f
C316 a_n2650_8322.n2 gnd 0.690258f
C317 a_n2650_8322.n3 gnd 0.391868f
C318 a_n2650_8322.t21 gnd 0.097992f
C319 a_n2650_8322.t15 gnd 0.097992f
C320 a_n2650_8322.n4 gnd 0.690258f
C321 a_n2650_8322.n5 gnd 0.391868f
C322 a_n2650_8322.t19 gnd 0.097992f
C323 a_n2650_8322.t17 gnd 0.097992f
C324 a_n2650_8322.n6 gnd 0.690258f
C325 a_n2650_8322.n7 gnd 0.391868f
C326 a_n2650_8322.t8 gnd 0.915724f
C327 a_n2650_8322.n8 gnd 1.70884f
C328 a_n2650_8322.t3 gnd 0.917551f
C329 a_n2650_8322.t7 gnd 0.097992f
C330 a_n2650_8322.t6 gnd 0.097992f
C331 a_n2650_8322.n9 gnd 0.690258f
C332 a_n2650_8322.n10 gnd 0.771262f
C333 a_n2650_8322.t1 gnd 0.915724f
C334 a_n2650_8322.n11 gnd 0.38811f
C335 a_n2650_8322.t4 gnd 0.915724f
C336 a_n2650_8322.n12 gnd 0.38811f
C337 a_n2650_8322.t2 gnd 0.097992f
C338 a_n2650_8322.t0 gnd 0.097992f
C339 a_n2650_8322.n13 gnd 0.690258f
C340 a_n2650_8322.n14 gnd 0.391868f
C341 a_n2650_8322.t5 gnd 0.915724f
C342 a_n2650_8322.n15 gnd 1.27333f
C343 a_n2650_8322.n16 gnd 2.0805f
C344 a_n2650_8322.n17 gnd 3.60069f
C345 a_n2650_8322.t22 gnd 0.915724f
C346 a_n2650_8322.n18 gnd 0.996043f
C347 a_n2650_8322.t12 gnd 0.097992f
C348 a_n2650_8322.t11 gnd 0.097992f
C349 a_n2650_8322.n19 gnd 0.690258f
C350 a_n2650_8322.n20 gnd 0.391868f
C351 a_n2650_8322.t24 gnd 0.097992f
C352 a_n2650_8322.t14 gnd 0.097992f
C353 a_n2650_8322.n21 gnd 0.690258f
C354 a_n2650_8322.n22 gnd 0.391868f
C355 a_n2650_8322.t25 gnd 0.917548f
C356 a_n2650_8322.t20 gnd 0.097992f
C357 a_n2650_8322.t16 gnd 0.097992f
C358 a_n2650_8322.n23 gnd 0.690258f
C359 a_n2650_8322.n24 gnd 0.771264f
C360 a_n2650_8322.n25 gnd 0.391867f
C361 a_n2650_8322.n26 gnd 0.69026f
C362 a_n2650_8322.t27 gnd 0.097992f
C363 output.t14 gnd 0.464308f
C364 output.t4 gnd 0.044422f
C365 output.t8 gnd 0.044422f
C366 output.n0 gnd 0.364624f
C367 output.n1 gnd 0.614102f
C368 output.t11 gnd 0.044422f
C369 output.t16 gnd 0.044422f
C370 output.n2 gnd 0.364624f
C371 output.n3 gnd 0.350265f
C372 output.t17 gnd 0.044422f
C373 output.t6 gnd 0.044422f
C374 output.n4 gnd 0.364624f
C375 output.n5 gnd 0.350265f
C376 output.t10 gnd 0.044422f
C377 output.t2 gnd 0.044422f
C378 output.n6 gnd 0.364624f
C379 output.n7 gnd 0.350265f
C380 output.t5 gnd 0.044422f
C381 output.t3 gnd 0.044422f
C382 output.n8 gnd 0.364624f
C383 output.n9 gnd 0.350265f
C384 output.t9 gnd 0.044422f
C385 output.t12 gnd 0.044422f
C386 output.n10 gnd 0.364624f
C387 output.n11 gnd 0.350265f
C388 output.t13 gnd 0.044422f
C389 output.t7 gnd 0.044422f
C390 output.n12 gnd 0.364624f
C391 output.n13 gnd 0.350265f
C392 output.t15 gnd 0.462979f
C393 output.n14 gnd 0.28994f
C394 output.n15 gnd 0.015803f
C395 output.n16 gnd 0.011243f
C396 output.n17 gnd 0.006041f
C397 output.n18 gnd 0.01428f
C398 output.n19 gnd 0.006397f
C399 output.n20 gnd 0.011243f
C400 output.n21 gnd 0.006041f
C401 output.n22 gnd 0.01428f
C402 output.n23 gnd 0.006397f
C403 output.n24 gnd 0.048111f
C404 output.t19 gnd 0.023274f
C405 output.n25 gnd 0.01071f
C406 output.n26 gnd 0.008435f
C407 output.n27 gnd 0.006041f
C408 output.n28 gnd 0.267512f
C409 output.n29 gnd 0.011243f
C410 output.n30 gnd 0.006041f
C411 output.n31 gnd 0.006397f
C412 output.n32 gnd 0.01428f
C413 output.n33 gnd 0.01428f
C414 output.n34 gnd 0.006397f
C415 output.n35 gnd 0.006041f
C416 output.n36 gnd 0.011243f
C417 output.n37 gnd 0.011243f
C418 output.n38 gnd 0.006041f
C419 output.n39 gnd 0.006397f
C420 output.n40 gnd 0.01428f
C421 output.n41 gnd 0.030913f
C422 output.n42 gnd 0.006397f
C423 output.n43 gnd 0.006041f
C424 output.n44 gnd 0.025987f
C425 output.n45 gnd 0.097665f
C426 output.n46 gnd 0.015803f
C427 output.n47 gnd 0.011243f
C428 output.n48 gnd 0.006041f
C429 output.n49 gnd 0.01428f
C430 output.n50 gnd 0.006397f
C431 output.n51 gnd 0.011243f
C432 output.n52 gnd 0.006041f
C433 output.n53 gnd 0.01428f
C434 output.n54 gnd 0.006397f
C435 output.n55 gnd 0.048111f
C436 output.t18 gnd 0.023274f
C437 output.n56 gnd 0.01071f
C438 output.n57 gnd 0.008435f
C439 output.n58 gnd 0.006041f
C440 output.n59 gnd 0.267512f
C441 output.n60 gnd 0.011243f
C442 output.n61 gnd 0.006041f
C443 output.n62 gnd 0.006397f
C444 output.n63 gnd 0.01428f
C445 output.n64 gnd 0.01428f
C446 output.n65 gnd 0.006397f
C447 output.n66 gnd 0.006041f
C448 output.n67 gnd 0.011243f
C449 output.n68 gnd 0.011243f
C450 output.n69 gnd 0.006041f
C451 output.n70 gnd 0.006397f
C452 output.n71 gnd 0.01428f
C453 output.n72 gnd 0.030913f
C454 output.n73 gnd 0.006397f
C455 output.n74 gnd 0.006041f
C456 output.n75 gnd 0.025987f
C457 output.n76 gnd 0.09306f
C458 output.n77 gnd 1.65264f
C459 output.n78 gnd 0.015803f
C460 output.n79 gnd 0.011243f
C461 output.n80 gnd 0.006041f
C462 output.n81 gnd 0.01428f
C463 output.n82 gnd 0.006397f
C464 output.n83 gnd 0.011243f
C465 output.n84 gnd 0.006041f
C466 output.n85 gnd 0.01428f
C467 output.n86 gnd 0.006397f
C468 output.n87 gnd 0.048111f
C469 output.t1 gnd 0.023274f
C470 output.n88 gnd 0.01071f
C471 output.n89 gnd 0.008435f
C472 output.n90 gnd 0.006041f
C473 output.n91 gnd 0.267512f
C474 output.n92 gnd 0.011243f
C475 output.n93 gnd 0.006041f
C476 output.n94 gnd 0.006397f
C477 output.n95 gnd 0.01428f
C478 output.n96 gnd 0.01428f
C479 output.n97 gnd 0.006397f
C480 output.n98 gnd 0.006041f
C481 output.n99 gnd 0.011243f
C482 output.n100 gnd 0.011243f
C483 output.n101 gnd 0.006041f
C484 output.n102 gnd 0.006397f
C485 output.n103 gnd 0.01428f
C486 output.n104 gnd 0.030913f
C487 output.n105 gnd 0.006397f
C488 output.n106 gnd 0.006041f
C489 output.n107 gnd 0.025987f
C490 output.n108 gnd 0.09306f
C491 output.n109 gnd 0.713089f
C492 output.n110 gnd 0.015803f
C493 output.n111 gnd 0.011243f
C494 output.n112 gnd 0.006041f
C495 output.n113 gnd 0.01428f
C496 output.n114 gnd 0.006397f
C497 output.n115 gnd 0.011243f
C498 output.n116 gnd 0.006041f
C499 output.n117 gnd 0.01428f
C500 output.n118 gnd 0.006397f
C501 output.n119 gnd 0.048111f
C502 output.t0 gnd 0.023274f
C503 output.n120 gnd 0.01071f
C504 output.n121 gnd 0.008435f
C505 output.n122 gnd 0.006041f
C506 output.n123 gnd 0.267512f
C507 output.n124 gnd 0.011243f
C508 output.n125 gnd 0.006041f
C509 output.n126 gnd 0.006397f
C510 output.n127 gnd 0.01428f
C511 output.n128 gnd 0.01428f
C512 output.n129 gnd 0.006397f
C513 output.n130 gnd 0.006041f
C514 output.n131 gnd 0.011243f
C515 output.n132 gnd 0.011243f
C516 output.n133 gnd 0.006041f
C517 output.n134 gnd 0.006397f
C518 output.n135 gnd 0.01428f
C519 output.n136 gnd 0.030913f
C520 output.n137 gnd 0.006397f
C521 output.n138 gnd 0.006041f
C522 output.n139 gnd 0.025987f
C523 output.n140 gnd 0.09306f
C524 output.n141 gnd 1.67353f
C525 diffpairibias.t27 gnd 0.090128f
C526 diffpairibias.t23 gnd 0.08996f
C527 diffpairibias.n0 gnd 0.105991f
C528 diffpairibias.t28 gnd 0.08996f
C529 diffpairibias.n1 gnd 0.051736f
C530 diffpairibias.t25 gnd 0.08996f
C531 diffpairibias.n2 gnd 0.051736f
C532 diffpairibias.t29 gnd 0.08996f
C533 diffpairibias.n3 gnd 0.041084f
C534 diffpairibias.t15 gnd 0.086371f
C535 diffpairibias.t1 gnd 0.085993f
C536 diffpairibias.n4 gnd 0.13579f
C537 diffpairibias.t11 gnd 0.085993f
C538 diffpairibias.n5 gnd 0.072463f
C539 diffpairibias.t13 gnd 0.085993f
C540 diffpairibias.n6 gnd 0.072463f
C541 diffpairibias.t7 gnd 0.085993f
C542 diffpairibias.n7 gnd 0.072463f
C543 diffpairibias.t3 gnd 0.085993f
C544 diffpairibias.n8 gnd 0.072463f
C545 diffpairibias.t17 gnd 0.085993f
C546 diffpairibias.n9 gnd 0.072463f
C547 diffpairibias.t5 gnd 0.085993f
C548 diffpairibias.n10 gnd 0.072463f
C549 diffpairibias.t19 gnd 0.085993f
C550 diffpairibias.n11 gnd 0.072463f
C551 diffpairibias.t9 gnd 0.085993f
C552 diffpairibias.n12 gnd 0.102883f
C553 diffpairibias.t14 gnd 0.086899f
C554 diffpairibias.t0 gnd 0.086748f
C555 diffpairibias.n13 gnd 0.094648f
C556 diffpairibias.t10 gnd 0.086748f
C557 diffpairibias.n14 gnd 0.052262f
C558 diffpairibias.t12 gnd 0.086748f
C559 diffpairibias.n15 gnd 0.052262f
C560 diffpairibias.t6 gnd 0.086748f
C561 diffpairibias.n16 gnd 0.052262f
C562 diffpairibias.t2 gnd 0.086748f
C563 diffpairibias.n17 gnd 0.052262f
C564 diffpairibias.t16 gnd 0.086748f
C565 diffpairibias.n18 gnd 0.052262f
C566 diffpairibias.t4 gnd 0.086748f
C567 diffpairibias.n19 gnd 0.052262f
C568 diffpairibias.t18 gnd 0.086748f
C569 diffpairibias.n20 gnd 0.052262f
C570 diffpairibias.t8 gnd 0.086748f
C571 diffpairibias.n21 gnd 0.061849f
C572 diffpairibias.n22 gnd 0.233513f
C573 diffpairibias.t20 gnd 0.08996f
C574 diffpairibias.n23 gnd 0.051747f
C575 diffpairibias.t26 gnd 0.08996f
C576 diffpairibias.n24 gnd 0.051736f
C577 diffpairibias.t22 gnd 0.08996f
C578 diffpairibias.n25 gnd 0.051736f
C579 diffpairibias.t21 gnd 0.08996f
C580 diffpairibias.n26 gnd 0.051736f
C581 diffpairibias.t24 gnd 0.08996f
C582 diffpairibias.n27 gnd 0.04729f
C583 diffpairibias.n28 gnd 0.047711f
C584 commonsourceibias.n0 gnd 0.010571f
C585 commonsourceibias.t92 gnd 0.160069f
C586 commonsourceibias.t106 gnd 0.148006f
C587 commonsourceibias.n1 gnd 0.006439f
C588 commonsourceibias.n2 gnd 0.007922f
C589 commonsourceibias.t119 gnd 0.148006f
C590 commonsourceibias.n3 gnd 0.008036f
C591 commonsourceibias.n4 gnd 0.007922f
C592 commonsourceibias.t84 gnd 0.148006f
C593 commonsourceibias.n5 gnd 0.059054f
C594 commonsourceibias.t100 gnd 0.148006f
C595 commonsourceibias.n6 gnd 0.006408f
C596 commonsourceibias.n7 gnd 0.007922f
C597 commonsourceibias.t114 gnd 0.148006f
C598 commonsourceibias.n8 gnd 0.007648f
C599 commonsourceibias.n9 gnd 0.007922f
C600 commonsourceibias.t80 gnd 0.148006f
C601 commonsourceibias.n10 gnd 0.059054f
C602 commonsourceibias.t76 gnd 0.148006f
C603 commonsourceibias.n11 gnd 0.006398f
C604 commonsourceibias.n12 gnd 0.010571f
C605 commonsourceibias.t60 gnd 0.160069f
C606 commonsourceibias.t14 gnd 0.148006f
C607 commonsourceibias.n13 gnd 0.006439f
C608 commonsourceibias.n14 gnd 0.007922f
C609 commonsourceibias.t38 gnd 0.148006f
C610 commonsourceibias.n15 gnd 0.008036f
C611 commonsourceibias.n16 gnd 0.007922f
C612 commonsourceibias.t4 gnd 0.148006f
C613 commonsourceibias.n17 gnd 0.059054f
C614 commonsourceibias.t28 gnd 0.148006f
C615 commonsourceibias.n18 gnd 0.006408f
C616 commonsourceibias.n19 gnd 0.007922f
C617 commonsourceibias.t62 gnd 0.148006f
C618 commonsourceibias.n20 gnd 0.007648f
C619 commonsourceibias.n21 gnd 0.007922f
C620 commonsourceibias.t18 gnd 0.148006f
C621 commonsourceibias.n22 gnd 0.059054f
C622 commonsourceibias.t26 gnd 0.148006f
C623 commonsourceibias.n23 gnd 0.006398f
C624 commonsourceibias.n24 gnd 0.007922f
C625 commonsourceibias.t6 gnd 0.148006f
C626 commonsourceibias.t32 gnd 0.148006f
C627 commonsourceibias.n25 gnd 0.059054f
C628 commonsourceibias.n26 gnd 0.007922f
C629 commonsourceibias.t42 gnd 0.148006f
C630 commonsourceibias.n27 gnd 0.059054f
C631 commonsourceibias.n28 gnd 0.007922f
C632 commonsourceibias.t20 gnd 0.148006f
C633 commonsourceibias.n29 gnd 0.059054f
C634 commonsourceibias.n30 gnd 0.007922f
C635 commonsourceibias.t30 gnd 0.148006f
C636 commonsourceibias.n31 gnd 0.009005f
C637 commonsourceibias.n32 gnd 0.007922f
C638 commonsourceibias.t56 gnd 0.148006f
C639 commonsourceibias.n33 gnd 0.010649f
C640 commonsourceibias.t16 gnd 0.164876f
C641 commonsourceibias.t12 gnd 0.148006f
C642 commonsourceibias.n34 gnd 0.065802f
C643 commonsourceibias.n35 gnd 0.070497f
C644 commonsourceibias.n36 gnd 0.03372f
C645 commonsourceibias.n37 gnd 0.007922f
C646 commonsourceibias.n38 gnd 0.006439f
C647 commonsourceibias.n39 gnd 0.010916f
C648 commonsourceibias.n40 gnd 0.059054f
C649 commonsourceibias.n41 gnd 0.010963f
C650 commonsourceibias.n42 gnd 0.007922f
C651 commonsourceibias.n43 gnd 0.007922f
C652 commonsourceibias.n44 gnd 0.007922f
C653 commonsourceibias.n45 gnd 0.008036f
C654 commonsourceibias.n46 gnd 0.059054f
C655 commonsourceibias.n47 gnd 0.009764f
C656 commonsourceibias.n48 gnd 0.010802f
C657 commonsourceibias.n49 gnd 0.007922f
C658 commonsourceibias.n50 gnd 0.007922f
C659 commonsourceibias.n51 gnd 0.010731f
C660 commonsourceibias.n52 gnd 0.006408f
C661 commonsourceibias.n53 gnd 0.010864f
C662 commonsourceibias.n54 gnd 0.007922f
C663 commonsourceibias.n55 gnd 0.007922f
C664 commonsourceibias.n56 gnd 0.010931f
C665 commonsourceibias.n57 gnd 0.009425f
C666 commonsourceibias.n58 gnd 0.007648f
C667 commonsourceibias.n59 gnd 0.007922f
C668 commonsourceibias.n60 gnd 0.007922f
C669 commonsourceibias.n61 gnd 0.00969f
C670 commonsourceibias.n62 gnd 0.010876f
C671 commonsourceibias.n63 gnd 0.059054f
C672 commonsourceibias.n64 gnd 0.010803f
C673 commonsourceibias.n65 gnd 0.007922f
C674 commonsourceibias.n66 gnd 0.007922f
C675 commonsourceibias.n67 gnd 0.007922f
C676 commonsourceibias.n68 gnd 0.010803f
C677 commonsourceibias.n69 gnd 0.059054f
C678 commonsourceibias.n70 gnd 0.010876f
C679 commonsourceibias.n71 gnd 0.00969f
C680 commonsourceibias.n72 gnd 0.007922f
C681 commonsourceibias.n73 gnd 0.007922f
C682 commonsourceibias.n74 gnd 0.007922f
C683 commonsourceibias.n75 gnd 0.009425f
C684 commonsourceibias.n76 gnd 0.010931f
C685 commonsourceibias.n77 gnd 0.059054f
C686 commonsourceibias.n78 gnd 0.010864f
C687 commonsourceibias.n79 gnd 0.007922f
C688 commonsourceibias.n80 gnd 0.007922f
C689 commonsourceibias.n81 gnd 0.007922f
C690 commonsourceibias.n82 gnd 0.010731f
C691 commonsourceibias.n83 gnd 0.059054f
C692 commonsourceibias.n84 gnd 0.010802f
C693 commonsourceibias.n85 gnd 0.009764f
C694 commonsourceibias.n86 gnd 0.007922f
C695 commonsourceibias.n87 gnd 0.007922f
C696 commonsourceibias.n88 gnd 0.007922f
C697 commonsourceibias.n89 gnd 0.009005f
C698 commonsourceibias.n90 gnd 0.010963f
C699 commonsourceibias.n91 gnd 0.059054f
C700 commonsourceibias.n92 gnd 0.010916f
C701 commonsourceibias.n93 gnd 0.007922f
C702 commonsourceibias.n94 gnd 0.007922f
C703 commonsourceibias.n95 gnd 0.007922f
C704 commonsourceibias.n96 gnd 0.010649f
C705 commonsourceibias.n97 gnd 0.059054f
C706 commonsourceibias.n98 gnd 0.010674f
C707 commonsourceibias.n99 gnd 0.071211f
C708 commonsourceibias.n100 gnd 0.079625f
C709 commonsourceibias.t61 gnd 0.017095f
C710 commonsourceibias.t15 gnd 0.017095f
C711 commonsourceibias.n101 gnd 0.151055f
C712 commonsourceibias.n102 gnd 0.130846f
C713 commonsourceibias.t39 gnd 0.017095f
C714 commonsourceibias.t5 gnd 0.017095f
C715 commonsourceibias.n103 gnd 0.151055f
C716 commonsourceibias.n104 gnd 0.069385f
C717 commonsourceibias.t29 gnd 0.017095f
C718 commonsourceibias.t63 gnd 0.017095f
C719 commonsourceibias.n105 gnd 0.151055f
C720 commonsourceibias.n106 gnd 0.069385f
C721 commonsourceibias.t19 gnd 0.017095f
C722 commonsourceibias.t27 gnd 0.017095f
C723 commonsourceibias.n107 gnd 0.151055f
C724 commonsourceibias.n108 gnd 0.057968f
C725 commonsourceibias.t13 gnd 0.017095f
C726 commonsourceibias.t17 gnd 0.017095f
C727 commonsourceibias.n109 gnd 0.15156f
C728 commonsourceibias.t31 gnd 0.017095f
C729 commonsourceibias.t57 gnd 0.017095f
C730 commonsourceibias.n110 gnd 0.151055f
C731 commonsourceibias.n111 gnd 0.140755f
C732 commonsourceibias.t43 gnd 0.017095f
C733 commonsourceibias.t21 gnd 0.017095f
C734 commonsourceibias.n112 gnd 0.151055f
C735 commonsourceibias.n113 gnd 0.069385f
C736 commonsourceibias.t7 gnd 0.017095f
C737 commonsourceibias.t33 gnd 0.017095f
C738 commonsourceibias.n114 gnd 0.151055f
C739 commonsourceibias.n115 gnd 0.057968f
C740 commonsourceibias.n116 gnd 0.070193f
C741 commonsourceibias.n117 gnd 0.007922f
C742 commonsourceibias.t105 gnd 0.148006f
C743 commonsourceibias.t121 gnd 0.148006f
C744 commonsourceibias.n118 gnd 0.059054f
C745 commonsourceibias.n119 gnd 0.007922f
C746 commonsourceibias.t71 gnd 0.148006f
C747 commonsourceibias.n120 gnd 0.059054f
C748 commonsourceibias.n121 gnd 0.007922f
C749 commonsourceibias.t99 gnd 0.148006f
C750 commonsourceibias.n122 gnd 0.059054f
C751 commonsourceibias.n123 gnd 0.007922f
C752 commonsourceibias.t95 gnd 0.148006f
C753 commonsourceibias.n124 gnd 0.009005f
C754 commonsourceibias.n125 gnd 0.007922f
C755 commonsourceibias.t109 gnd 0.148006f
C756 commonsourceibias.n126 gnd 0.010649f
C757 commonsourceibias.t85 gnd 0.164876f
C758 commonsourceibias.t89 gnd 0.148006f
C759 commonsourceibias.n127 gnd 0.065802f
C760 commonsourceibias.n128 gnd 0.070497f
C761 commonsourceibias.n129 gnd 0.03372f
C762 commonsourceibias.n130 gnd 0.007922f
C763 commonsourceibias.n131 gnd 0.006439f
C764 commonsourceibias.n132 gnd 0.010916f
C765 commonsourceibias.n133 gnd 0.059054f
C766 commonsourceibias.n134 gnd 0.010963f
C767 commonsourceibias.n135 gnd 0.007922f
C768 commonsourceibias.n136 gnd 0.007922f
C769 commonsourceibias.n137 gnd 0.007922f
C770 commonsourceibias.n138 gnd 0.008036f
C771 commonsourceibias.n139 gnd 0.059054f
C772 commonsourceibias.n140 gnd 0.009764f
C773 commonsourceibias.n141 gnd 0.010802f
C774 commonsourceibias.n142 gnd 0.007922f
C775 commonsourceibias.n143 gnd 0.007922f
C776 commonsourceibias.n144 gnd 0.010731f
C777 commonsourceibias.n145 gnd 0.006408f
C778 commonsourceibias.n146 gnd 0.010864f
C779 commonsourceibias.n147 gnd 0.007922f
C780 commonsourceibias.n148 gnd 0.007922f
C781 commonsourceibias.n149 gnd 0.010931f
C782 commonsourceibias.n150 gnd 0.009425f
C783 commonsourceibias.n151 gnd 0.007648f
C784 commonsourceibias.n152 gnd 0.007922f
C785 commonsourceibias.n153 gnd 0.007922f
C786 commonsourceibias.n154 gnd 0.00969f
C787 commonsourceibias.n155 gnd 0.010876f
C788 commonsourceibias.n156 gnd 0.059054f
C789 commonsourceibias.n157 gnd 0.010803f
C790 commonsourceibias.n158 gnd 0.007884f
C791 commonsourceibias.n159 gnd 0.057266f
C792 commonsourceibias.n160 gnd 0.007884f
C793 commonsourceibias.n161 gnd 0.010803f
C794 commonsourceibias.n162 gnd 0.059054f
C795 commonsourceibias.n163 gnd 0.010876f
C796 commonsourceibias.n164 gnd 0.00969f
C797 commonsourceibias.n165 gnd 0.007922f
C798 commonsourceibias.n166 gnd 0.007922f
C799 commonsourceibias.n167 gnd 0.007922f
C800 commonsourceibias.n168 gnd 0.009425f
C801 commonsourceibias.n169 gnd 0.010931f
C802 commonsourceibias.n170 gnd 0.059054f
C803 commonsourceibias.n171 gnd 0.010864f
C804 commonsourceibias.n172 gnd 0.007922f
C805 commonsourceibias.n173 gnd 0.007922f
C806 commonsourceibias.n174 gnd 0.007922f
C807 commonsourceibias.n175 gnd 0.010731f
C808 commonsourceibias.n176 gnd 0.059054f
C809 commonsourceibias.n177 gnd 0.010802f
C810 commonsourceibias.n178 gnd 0.009764f
C811 commonsourceibias.n179 gnd 0.007922f
C812 commonsourceibias.n180 gnd 0.007922f
C813 commonsourceibias.n181 gnd 0.007922f
C814 commonsourceibias.n182 gnd 0.009005f
C815 commonsourceibias.n183 gnd 0.010963f
C816 commonsourceibias.n184 gnd 0.059054f
C817 commonsourceibias.n185 gnd 0.010916f
C818 commonsourceibias.n186 gnd 0.007922f
C819 commonsourceibias.n187 gnd 0.007922f
C820 commonsourceibias.n188 gnd 0.007922f
C821 commonsourceibias.n189 gnd 0.010649f
C822 commonsourceibias.n190 gnd 0.059054f
C823 commonsourceibias.n191 gnd 0.010674f
C824 commonsourceibias.n192 gnd 0.071211f
C825 commonsourceibias.n193 gnd 0.047027f
C826 commonsourceibias.n194 gnd 0.010571f
C827 commonsourceibias.t94 gnd 0.148006f
C828 commonsourceibias.n195 gnd 0.006439f
C829 commonsourceibias.n196 gnd 0.007922f
C830 commonsourceibias.t107 gnd 0.148006f
C831 commonsourceibias.n197 gnd 0.008036f
C832 commonsourceibias.n198 gnd 0.007922f
C833 commonsourceibias.t74 gnd 0.148006f
C834 commonsourceibias.n199 gnd 0.059054f
C835 commonsourceibias.t87 gnd 0.148006f
C836 commonsourceibias.n200 gnd 0.006408f
C837 commonsourceibias.n201 gnd 0.007922f
C838 commonsourceibias.t101 gnd 0.148006f
C839 commonsourceibias.n202 gnd 0.007648f
C840 commonsourceibias.n203 gnd 0.007922f
C841 commonsourceibias.t70 gnd 0.148006f
C842 commonsourceibias.n204 gnd 0.059054f
C843 commonsourceibias.t67 gnd 0.148006f
C844 commonsourceibias.n205 gnd 0.006398f
C845 commonsourceibias.n206 gnd 0.007922f
C846 commonsourceibias.t93 gnd 0.148006f
C847 commonsourceibias.t108 gnd 0.148006f
C848 commonsourceibias.n207 gnd 0.059054f
C849 commonsourceibias.n208 gnd 0.007922f
C850 commonsourceibias.t127 gnd 0.148006f
C851 commonsourceibias.n209 gnd 0.059054f
C852 commonsourceibias.n210 gnd 0.007922f
C853 commonsourceibias.t86 gnd 0.148006f
C854 commonsourceibias.n211 gnd 0.059054f
C855 commonsourceibias.n212 gnd 0.007922f
C856 commonsourceibias.t82 gnd 0.148006f
C857 commonsourceibias.n213 gnd 0.009005f
C858 commonsourceibias.n214 gnd 0.007922f
C859 commonsourceibias.t96 gnd 0.148006f
C860 commonsourceibias.n215 gnd 0.010649f
C861 commonsourceibias.t75 gnd 0.164876f
C862 commonsourceibias.t77 gnd 0.148006f
C863 commonsourceibias.n216 gnd 0.065802f
C864 commonsourceibias.n217 gnd 0.070497f
C865 commonsourceibias.n218 gnd 0.03372f
C866 commonsourceibias.n219 gnd 0.007922f
C867 commonsourceibias.n220 gnd 0.006439f
C868 commonsourceibias.n221 gnd 0.010916f
C869 commonsourceibias.n222 gnd 0.059054f
C870 commonsourceibias.n223 gnd 0.010963f
C871 commonsourceibias.n224 gnd 0.007922f
C872 commonsourceibias.n225 gnd 0.007922f
C873 commonsourceibias.n226 gnd 0.007922f
C874 commonsourceibias.n227 gnd 0.008036f
C875 commonsourceibias.n228 gnd 0.059054f
C876 commonsourceibias.n229 gnd 0.009764f
C877 commonsourceibias.n230 gnd 0.010802f
C878 commonsourceibias.n231 gnd 0.007922f
C879 commonsourceibias.n232 gnd 0.007922f
C880 commonsourceibias.n233 gnd 0.010731f
C881 commonsourceibias.n234 gnd 0.006408f
C882 commonsourceibias.n235 gnd 0.010864f
C883 commonsourceibias.n236 gnd 0.007922f
C884 commonsourceibias.n237 gnd 0.007922f
C885 commonsourceibias.n238 gnd 0.010931f
C886 commonsourceibias.n239 gnd 0.009425f
C887 commonsourceibias.n240 gnd 0.007648f
C888 commonsourceibias.n241 gnd 0.007922f
C889 commonsourceibias.n242 gnd 0.007922f
C890 commonsourceibias.n243 gnd 0.00969f
C891 commonsourceibias.n244 gnd 0.010876f
C892 commonsourceibias.n245 gnd 0.059054f
C893 commonsourceibias.n246 gnd 0.010803f
C894 commonsourceibias.n247 gnd 0.007922f
C895 commonsourceibias.n248 gnd 0.007922f
C896 commonsourceibias.n249 gnd 0.007922f
C897 commonsourceibias.n250 gnd 0.010803f
C898 commonsourceibias.n251 gnd 0.059054f
C899 commonsourceibias.n252 gnd 0.010876f
C900 commonsourceibias.n253 gnd 0.00969f
C901 commonsourceibias.n254 gnd 0.007922f
C902 commonsourceibias.n255 gnd 0.007922f
C903 commonsourceibias.n256 gnd 0.007922f
C904 commonsourceibias.n257 gnd 0.009425f
C905 commonsourceibias.n258 gnd 0.010931f
C906 commonsourceibias.n259 gnd 0.059054f
C907 commonsourceibias.n260 gnd 0.010864f
C908 commonsourceibias.n261 gnd 0.007922f
C909 commonsourceibias.n262 gnd 0.007922f
C910 commonsourceibias.n263 gnd 0.007922f
C911 commonsourceibias.n264 gnd 0.010731f
C912 commonsourceibias.n265 gnd 0.059054f
C913 commonsourceibias.n266 gnd 0.010802f
C914 commonsourceibias.n267 gnd 0.009764f
C915 commonsourceibias.n268 gnd 0.007922f
C916 commonsourceibias.n269 gnd 0.007922f
C917 commonsourceibias.n270 gnd 0.007922f
C918 commonsourceibias.n271 gnd 0.009005f
C919 commonsourceibias.n272 gnd 0.010963f
C920 commonsourceibias.n273 gnd 0.059054f
C921 commonsourceibias.n274 gnd 0.010916f
C922 commonsourceibias.n275 gnd 0.007922f
C923 commonsourceibias.n276 gnd 0.007922f
C924 commonsourceibias.n277 gnd 0.007922f
C925 commonsourceibias.n278 gnd 0.010649f
C926 commonsourceibias.n279 gnd 0.059054f
C927 commonsourceibias.n280 gnd 0.010674f
C928 commonsourceibias.t81 gnd 0.160069f
C929 commonsourceibias.n281 gnd 0.071211f
C930 commonsourceibias.n282 gnd 0.025411f
C931 commonsourceibias.n283 gnd 0.458519f
C932 commonsourceibias.n284 gnd 0.010571f
C933 commonsourceibias.t110 gnd 0.160069f
C934 commonsourceibias.t123 gnd 0.148006f
C935 commonsourceibias.n285 gnd 0.006439f
C936 commonsourceibias.n286 gnd 0.007922f
C937 commonsourceibias.t68 gnd 0.148006f
C938 commonsourceibias.n287 gnd 0.008036f
C939 commonsourceibias.n288 gnd 0.007922f
C940 commonsourceibias.t117 gnd 0.148006f
C941 commonsourceibias.n289 gnd 0.006408f
C942 commonsourceibias.n290 gnd 0.007922f
C943 commonsourceibias.t64 gnd 0.148006f
C944 commonsourceibias.n291 gnd 0.007648f
C945 commonsourceibias.n292 gnd 0.007922f
C946 commonsourceibias.t90 gnd 0.148006f
C947 commonsourceibias.n293 gnd 0.006398f
C948 commonsourceibias.n294 gnd 0.007922f
C949 commonsourceibias.t122 gnd 0.148006f
C950 commonsourceibias.t69 gnd 0.148006f
C951 commonsourceibias.n295 gnd 0.059054f
C952 commonsourceibias.n296 gnd 0.007922f
C953 commonsourceibias.t66 gnd 0.148006f
C954 commonsourceibias.n297 gnd 0.059054f
C955 commonsourceibias.n298 gnd 0.007922f
C956 commonsourceibias.t116 gnd 0.148006f
C957 commonsourceibias.n299 gnd 0.059054f
C958 commonsourceibias.n300 gnd 0.007922f
C959 commonsourceibias.t113 gnd 0.148006f
C960 commonsourceibias.n301 gnd 0.009005f
C961 commonsourceibias.n302 gnd 0.007922f
C962 commonsourceibias.t126 gnd 0.148006f
C963 commonsourceibias.n303 gnd 0.010649f
C964 commonsourceibias.t91 gnd 0.164876f
C965 commonsourceibias.t83 gnd 0.148006f
C966 commonsourceibias.n304 gnd 0.065802f
C967 commonsourceibias.n305 gnd 0.070497f
C968 commonsourceibias.n306 gnd 0.03372f
C969 commonsourceibias.n307 gnd 0.007922f
C970 commonsourceibias.n308 gnd 0.006439f
C971 commonsourceibias.n309 gnd 0.010916f
C972 commonsourceibias.n310 gnd 0.059054f
C973 commonsourceibias.n311 gnd 0.010963f
C974 commonsourceibias.n312 gnd 0.007922f
C975 commonsourceibias.n313 gnd 0.007922f
C976 commonsourceibias.n314 gnd 0.007922f
C977 commonsourceibias.n315 gnd 0.008036f
C978 commonsourceibias.n316 gnd 0.059054f
C979 commonsourceibias.n317 gnd 0.009764f
C980 commonsourceibias.n318 gnd 0.010802f
C981 commonsourceibias.n319 gnd 0.007922f
C982 commonsourceibias.n320 gnd 0.007922f
C983 commonsourceibias.n321 gnd 0.010731f
C984 commonsourceibias.n322 gnd 0.006408f
C985 commonsourceibias.n323 gnd 0.010864f
C986 commonsourceibias.n324 gnd 0.007922f
C987 commonsourceibias.n325 gnd 0.007922f
C988 commonsourceibias.n326 gnd 0.010931f
C989 commonsourceibias.n327 gnd 0.009425f
C990 commonsourceibias.n328 gnd 0.007648f
C991 commonsourceibias.n329 gnd 0.007922f
C992 commonsourceibias.n330 gnd 0.007922f
C993 commonsourceibias.n331 gnd 0.00969f
C994 commonsourceibias.n332 gnd 0.010876f
C995 commonsourceibias.n333 gnd 0.059054f
C996 commonsourceibias.n334 gnd 0.010803f
C997 commonsourceibias.n335 gnd 0.007884f
C998 commonsourceibias.t55 gnd 0.017095f
C999 commonsourceibias.t53 gnd 0.017095f
C1000 commonsourceibias.n336 gnd 0.15156f
C1001 commonsourceibias.t3 gnd 0.017095f
C1002 commonsourceibias.t49 gnd 0.017095f
C1003 commonsourceibias.n337 gnd 0.151055f
C1004 commonsourceibias.n338 gnd 0.140755f
C1005 commonsourceibias.t41 gnd 0.017095f
C1006 commonsourceibias.t59 gnd 0.017095f
C1007 commonsourceibias.n339 gnd 0.151055f
C1008 commonsourceibias.n340 gnd 0.069385f
C1009 commonsourceibias.t51 gnd 0.017095f
C1010 commonsourceibias.t25 gnd 0.017095f
C1011 commonsourceibias.n341 gnd 0.151055f
C1012 commonsourceibias.n342 gnd 0.057968f
C1013 commonsourceibias.n343 gnd 0.010571f
C1014 commonsourceibias.t34 gnd 0.148006f
C1015 commonsourceibias.n344 gnd 0.006439f
C1016 commonsourceibias.n345 gnd 0.007922f
C1017 commonsourceibias.t0 gnd 0.148006f
C1018 commonsourceibias.n346 gnd 0.008036f
C1019 commonsourceibias.n347 gnd 0.007922f
C1020 commonsourceibias.t46 gnd 0.148006f
C1021 commonsourceibias.n348 gnd 0.006408f
C1022 commonsourceibias.n349 gnd 0.007922f
C1023 commonsourceibias.t10 gnd 0.148006f
C1024 commonsourceibias.n350 gnd 0.007648f
C1025 commonsourceibias.n351 gnd 0.007922f
C1026 commonsourceibias.t44 gnd 0.148006f
C1027 commonsourceibias.n352 gnd 0.006398f
C1028 commonsourceibias.n353 gnd 0.007922f
C1029 commonsourceibias.t24 gnd 0.148006f
C1030 commonsourceibias.t50 gnd 0.148006f
C1031 commonsourceibias.n354 gnd 0.059054f
C1032 commonsourceibias.n355 gnd 0.007922f
C1033 commonsourceibias.t58 gnd 0.148006f
C1034 commonsourceibias.n356 gnd 0.059054f
C1035 commonsourceibias.n357 gnd 0.007922f
C1036 commonsourceibias.t40 gnd 0.148006f
C1037 commonsourceibias.n358 gnd 0.059054f
C1038 commonsourceibias.n359 gnd 0.007922f
C1039 commonsourceibias.t48 gnd 0.148006f
C1040 commonsourceibias.n360 gnd 0.009005f
C1041 commonsourceibias.n361 gnd 0.007922f
C1042 commonsourceibias.t2 gnd 0.148006f
C1043 commonsourceibias.n362 gnd 0.010649f
C1044 commonsourceibias.t54 gnd 0.164876f
C1045 commonsourceibias.t52 gnd 0.148006f
C1046 commonsourceibias.n363 gnd 0.065802f
C1047 commonsourceibias.n364 gnd 0.070497f
C1048 commonsourceibias.n365 gnd 0.03372f
C1049 commonsourceibias.n366 gnd 0.007922f
C1050 commonsourceibias.n367 gnd 0.006439f
C1051 commonsourceibias.n368 gnd 0.010916f
C1052 commonsourceibias.n369 gnd 0.059054f
C1053 commonsourceibias.n370 gnd 0.010963f
C1054 commonsourceibias.n371 gnd 0.007922f
C1055 commonsourceibias.n372 gnd 0.007922f
C1056 commonsourceibias.n373 gnd 0.007922f
C1057 commonsourceibias.n374 gnd 0.008036f
C1058 commonsourceibias.n375 gnd 0.059054f
C1059 commonsourceibias.n376 gnd 0.009764f
C1060 commonsourceibias.n377 gnd 0.010802f
C1061 commonsourceibias.n378 gnd 0.007922f
C1062 commonsourceibias.n379 gnd 0.007922f
C1063 commonsourceibias.n380 gnd 0.010731f
C1064 commonsourceibias.n381 gnd 0.006408f
C1065 commonsourceibias.n382 gnd 0.010864f
C1066 commonsourceibias.n383 gnd 0.007922f
C1067 commonsourceibias.n384 gnd 0.007922f
C1068 commonsourceibias.n385 gnd 0.010931f
C1069 commonsourceibias.n386 gnd 0.009425f
C1070 commonsourceibias.n387 gnd 0.007648f
C1071 commonsourceibias.n388 gnd 0.007922f
C1072 commonsourceibias.n389 gnd 0.007922f
C1073 commonsourceibias.n390 gnd 0.00969f
C1074 commonsourceibias.n391 gnd 0.010876f
C1075 commonsourceibias.n392 gnd 0.059054f
C1076 commonsourceibias.n393 gnd 0.010803f
C1077 commonsourceibias.n394 gnd 0.007922f
C1078 commonsourceibias.n395 gnd 0.007922f
C1079 commonsourceibias.n396 gnd 0.007922f
C1080 commonsourceibias.n397 gnd 0.010803f
C1081 commonsourceibias.n398 gnd 0.059054f
C1082 commonsourceibias.n399 gnd 0.010876f
C1083 commonsourceibias.t36 gnd 0.148006f
C1084 commonsourceibias.n400 gnd 0.059054f
C1085 commonsourceibias.n401 gnd 0.00969f
C1086 commonsourceibias.n402 gnd 0.007922f
C1087 commonsourceibias.n403 gnd 0.007922f
C1088 commonsourceibias.n404 gnd 0.007922f
C1089 commonsourceibias.n405 gnd 0.009425f
C1090 commonsourceibias.n406 gnd 0.010931f
C1091 commonsourceibias.n407 gnd 0.059054f
C1092 commonsourceibias.n408 gnd 0.010864f
C1093 commonsourceibias.n409 gnd 0.007922f
C1094 commonsourceibias.n410 gnd 0.007922f
C1095 commonsourceibias.n411 gnd 0.007922f
C1096 commonsourceibias.n412 gnd 0.010731f
C1097 commonsourceibias.n413 gnd 0.059054f
C1098 commonsourceibias.n414 gnd 0.010802f
C1099 commonsourceibias.t22 gnd 0.148006f
C1100 commonsourceibias.n415 gnd 0.059054f
C1101 commonsourceibias.n416 gnd 0.009764f
C1102 commonsourceibias.n417 gnd 0.007922f
C1103 commonsourceibias.n418 gnd 0.007922f
C1104 commonsourceibias.n419 gnd 0.007922f
C1105 commonsourceibias.n420 gnd 0.009005f
C1106 commonsourceibias.n421 gnd 0.010963f
C1107 commonsourceibias.n422 gnd 0.059054f
C1108 commonsourceibias.n423 gnd 0.010916f
C1109 commonsourceibias.n424 gnd 0.007922f
C1110 commonsourceibias.n425 gnd 0.007922f
C1111 commonsourceibias.n426 gnd 0.007922f
C1112 commonsourceibias.n427 gnd 0.010649f
C1113 commonsourceibias.n428 gnd 0.059054f
C1114 commonsourceibias.n429 gnd 0.010674f
C1115 commonsourceibias.t8 gnd 0.160069f
C1116 commonsourceibias.n430 gnd 0.071211f
C1117 commonsourceibias.n431 gnd 0.079625f
C1118 commonsourceibias.t35 gnd 0.017095f
C1119 commonsourceibias.t9 gnd 0.017095f
C1120 commonsourceibias.n432 gnd 0.151055f
C1121 commonsourceibias.n433 gnd 0.130846f
C1122 commonsourceibias.t23 gnd 0.017095f
C1123 commonsourceibias.t1 gnd 0.017095f
C1124 commonsourceibias.n434 gnd 0.151055f
C1125 commonsourceibias.n435 gnd 0.069385f
C1126 commonsourceibias.t11 gnd 0.017095f
C1127 commonsourceibias.t47 gnd 0.017095f
C1128 commonsourceibias.n436 gnd 0.151055f
C1129 commonsourceibias.n437 gnd 0.069385f
C1130 commonsourceibias.t45 gnd 0.017095f
C1131 commonsourceibias.t37 gnd 0.017095f
C1132 commonsourceibias.n438 gnd 0.151055f
C1133 commonsourceibias.n439 gnd 0.057968f
C1134 commonsourceibias.n440 gnd 0.070193f
C1135 commonsourceibias.n441 gnd 0.057266f
C1136 commonsourceibias.n442 gnd 0.007884f
C1137 commonsourceibias.n443 gnd 0.010803f
C1138 commonsourceibias.n444 gnd 0.059054f
C1139 commonsourceibias.n445 gnd 0.010876f
C1140 commonsourceibias.t72 gnd 0.148006f
C1141 commonsourceibias.n446 gnd 0.059054f
C1142 commonsourceibias.n447 gnd 0.00969f
C1143 commonsourceibias.n448 gnd 0.007922f
C1144 commonsourceibias.n449 gnd 0.007922f
C1145 commonsourceibias.n450 gnd 0.007922f
C1146 commonsourceibias.n451 gnd 0.009425f
C1147 commonsourceibias.n452 gnd 0.010931f
C1148 commonsourceibias.n453 gnd 0.059054f
C1149 commonsourceibias.n454 gnd 0.010864f
C1150 commonsourceibias.n455 gnd 0.007922f
C1151 commonsourceibias.n456 gnd 0.007922f
C1152 commonsourceibias.n457 gnd 0.007922f
C1153 commonsourceibias.n458 gnd 0.010731f
C1154 commonsourceibias.n459 gnd 0.059054f
C1155 commonsourceibias.n460 gnd 0.010802f
C1156 commonsourceibias.t102 gnd 0.148006f
C1157 commonsourceibias.n461 gnd 0.059054f
C1158 commonsourceibias.n462 gnd 0.009764f
C1159 commonsourceibias.n463 gnd 0.007922f
C1160 commonsourceibias.n464 gnd 0.007922f
C1161 commonsourceibias.n465 gnd 0.007922f
C1162 commonsourceibias.n466 gnd 0.009005f
C1163 commonsourceibias.n467 gnd 0.010963f
C1164 commonsourceibias.n468 gnd 0.059054f
C1165 commonsourceibias.n469 gnd 0.010916f
C1166 commonsourceibias.n470 gnd 0.007922f
C1167 commonsourceibias.n471 gnd 0.007922f
C1168 commonsourceibias.n472 gnd 0.007922f
C1169 commonsourceibias.n473 gnd 0.010649f
C1170 commonsourceibias.n474 gnd 0.059054f
C1171 commonsourceibias.n475 gnd 0.010674f
C1172 commonsourceibias.n476 gnd 0.071211f
C1173 commonsourceibias.n477 gnd 0.047027f
C1174 commonsourceibias.n478 gnd 0.010571f
C1175 commonsourceibias.t112 gnd 0.148006f
C1176 commonsourceibias.n479 gnd 0.006439f
C1177 commonsourceibias.n480 gnd 0.007922f
C1178 commonsourceibias.t124 gnd 0.148006f
C1179 commonsourceibias.n481 gnd 0.008036f
C1180 commonsourceibias.n482 gnd 0.007922f
C1181 commonsourceibias.t104 gnd 0.148006f
C1182 commonsourceibias.n483 gnd 0.006408f
C1183 commonsourceibias.n484 gnd 0.007922f
C1184 commonsourceibias.t118 gnd 0.148006f
C1185 commonsourceibias.n485 gnd 0.007648f
C1186 commonsourceibias.n486 gnd 0.007922f
C1187 commonsourceibias.t79 gnd 0.148006f
C1188 commonsourceibias.n487 gnd 0.006398f
C1189 commonsourceibias.n488 gnd 0.007922f
C1190 commonsourceibias.t111 gnd 0.148006f
C1191 commonsourceibias.t125 gnd 0.148006f
C1192 commonsourceibias.n489 gnd 0.059054f
C1193 commonsourceibias.n490 gnd 0.007922f
C1194 commonsourceibias.t120 gnd 0.148006f
C1195 commonsourceibias.n491 gnd 0.059054f
C1196 commonsourceibias.n492 gnd 0.007922f
C1197 commonsourceibias.t103 gnd 0.148006f
C1198 commonsourceibias.n493 gnd 0.059054f
C1199 commonsourceibias.n494 gnd 0.007922f
C1200 commonsourceibias.t98 gnd 0.148006f
C1201 commonsourceibias.n495 gnd 0.009005f
C1202 commonsourceibias.n496 gnd 0.007922f
C1203 commonsourceibias.t115 gnd 0.148006f
C1204 commonsourceibias.n497 gnd 0.010649f
C1205 commonsourceibias.t78 gnd 0.164876f
C1206 commonsourceibias.t73 gnd 0.148006f
C1207 commonsourceibias.n498 gnd 0.065802f
C1208 commonsourceibias.n499 gnd 0.070497f
C1209 commonsourceibias.n500 gnd 0.03372f
C1210 commonsourceibias.n501 gnd 0.007922f
C1211 commonsourceibias.n502 gnd 0.006439f
C1212 commonsourceibias.n503 gnd 0.010916f
C1213 commonsourceibias.n504 gnd 0.059054f
C1214 commonsourceibias.n505 gnd 0.010963f
C1215 commonsourceibias.n506 gnd 0.007922f
C1216 commonsourceibias.n507 gnd 0.007922f
C1217 commonsourceibias.n508 gnd 0.007922f
C1218 commonsourceibias.n509 gnd 0.008036f
C1219 commonsourceibias.n510 gnd 0.059054f
C1220 commonsourceibias.n511 gnd 0.009764f
C1221 commonsourceibias.n512 gnd 0.010802f
C1222 commonsourceibias.n513 gnd 0.007922f
C1223 commonsourceibias.n514 gnd 0.007922f
C1224 commonsourceibias.n515 gnd 0.010731f
C1225 commonsourceibias.n516 gnd 0.006408f
C1226 commonsourceibias.n517 gnd 0.010864f
C1227 commonsourceibias.n518 gnd 0.007922f
C1228 commonsourceibias.n519 gnd 0.007922f
C1229 commonsourceibias.n520 gnd 0.010931f
C1230 commonsourceibias.n521 gnd 0.009425f
C1231 commonsourceibias.n522 gnd 0.007648f
C1232 commonsourceibias.n523 gnd 0.007922f
C1233 commonsourceibias.n524 gnd 0.007922f
C1234 commonsourceibias.n525 gnd 0.00969f
C1235 commonsourceibias.n526 gnd 0.010876f
C1236 commonsourceibias.n527 gnd 0.059054f
C1237 commonsourceibias.n528 gnd 0.010803f
C1238 commonsourceibias.n529 gnd 0.007922f
C1239 commonsourceibias.n530 gnd 0.007922f
C1240 commonsourceibias.n531 gnd 0.007922f
C1241 commonsourceibias.n532 gnd 0.010803f
C1242 commonsourceibias.n533 gnd 0.059054f
C1243 commonsourceibias.n534 gnd 0.010876f
C1244 commonsourceibias.t65 gnd 0.148006f
C1245 commonsourceibias.n535 gnd 0.059054f
C1246 commonsourceibias.n536 gnd 0.00969f
C1247 commonsourceibias.n537 gnd 0.007922f
C1248 commonsourceibias.n538 gnd 0.007922f
C1249 commonsourceibias.n539 gnd 0.007922f
C1250 commonsourceibias.n540 gnd 0.009425f
C1251 commonsourceibias.n541 gnd 0.010931f
C1252 commonsourceibias.n542 gnd 0.059054f
C1253 commonsourceibias.n543 gnd 0.010864f
C1254 commonsourceibias.n544 gnd 0.007922f
C1255 commonsourceibias.n545 gnd 0.007922f
C1256 commonsourceibias.n546 gnd 0.007922f
C1257 commonsourceibias.n547 gnd 0.010731f
C1258 commonsourceibias.n548 gnd 0.059054f
C1259 commonsourceibias.n549 gnd 0.010802f
C1260 commonsourceibias.t88 gnd 0.148006f
C1261 commonsourceibias.n550 gnd 0.059054f
C1262 commonsourceibias.n551 gnd 0.009764f
C1263 commonsourceibias.n552 gnd 0.007922f
C1264 commonsourceibias.n553 gnd 0.007922f
C1265 commonsourceibias.n554 gnd 0.007922f
C1266 commonsourceibias.n555 gnd 0.009005f
C1267 commonsourceibias.n556 gnd 0.010963f
C1268 commonsourceibias.n557 gnd 0.059054f
C1269 commonsourceibias.n558 gnd 0.010916f
C1270 commonsourceibias.n559 gnd 0.007922f
C1271 commonsourceibias.n560 gnd 0.007922f
C1272 commonsourceibias.n561 gnd 0.007922f
C1273 commonsourceibias.n562 gnd 0.010649f
C1274 commonsourceibias.n563 gnd 0.059054f
C1275 commonsourceibias.n564 gnd 0.010674f
C1276 commonsourceibias.t97 gnd 0.160069f
C1277 commonsourceibias.n565 gnd 0.071211f
C1278 commonsourceibias.n566 gnd 0.025411f
C1279 commonsourceibias.n567 gnd 0.219034f
C1280 commonsourceibias.n568 gnd 4.63083f
C1281 a_n3827_n3924.t23 gnd 0.089565f
C1282 a_n3827_n3924.t33 gnd 0.930867f
C1283 a_n3827_n3924.n0 gnd 0.351909f
C1284 a_n3827_n3924.t15 gnd 1.15846f
C1285 a_n3827_n3924.n1 gnd 1.34803f
C1286 a_n3827_n3924.t2 gnd 0.930867f
C1287 a_n3827_n3924.n2 gnd 0.351909f
C1288 a_n3827_n3924.t6 gnd 0.089565f
C1289 a_n3827_n3924.t5 gnd 0.089565f
C1290 a_n3827_n3924.n3 gnd 0.731494f
C1291 a_n3827_n3924.n4 gnd 0.368632f
C1292 a_n3827_n3924.t0 gnd 0.089565f
C1293 a_n3827_n3924.t19 gnd 0.089565f
C1294 a_n3827_n3924.n5 gnd 0.731494f
C1295 a_n3827_n3924.n6 gnd 0.368632f
C1296 a_n3827_n3924.t1 gnd 0.089565f
C1297 a_n3827_n3924.t4 gnd 0.089565f
C1298 a_n3827_n3924.n7 gnd 0.731494f
C1299 a_n3827_n3924.n8 gnd 0.368632f
C1300 a_n3827_n3924.t49 gnd 0.089565f
C1301 a_n3827_n3924.t47 gnd 0.089565f
C1302 a_n3827_n3924.n9 gnd 0.731494f
C1303 a_n3827_n3924.n10 gnd 0.368632f
C1304 a_n3827_n3924.t44 gnd 0.930867f
C1305 a_n3827_n3924.n11 gnd 0.871363f
C1306 a_n3827_n3924.t17 gnd 1.15823f
C1307 a_n3827_n3924.t7 gnd 1.15658f
C1308 a_n3827_n3924.n12 gnd 1.17173f
C1309 a_n3827_n3924.t12 gnd 1.15658f
C1310 a_n3827_n3924.n13 gnd 0.610864f
C1311 a_n3827_n3924.t10 gnd 1.15658f
C1312 a_n3827_n3924.n14 gnd 0.8146f
C1313 a_n3827_n3924.t42 gnd 1.15658f
C1314 a_n3827_n3924.n15 gnd 0.8146f
C1315 a_n3827_n3924.t14 gnd 1.15658f
C1316 a_n3827_n3924.n16 gnd 0.8146f
C1317 a_n3827_n3924.t48 gnd 1.15658f
C1318 a_n3827_n3924.n17 gnd 0.8146f
C1319 a_n3827_n3924.t9 gnd 1.15658f
C1320 a_n3827_n3924.n18 gnd 0.8146f
C1321 a_n3827_n3924.t8 gnd 1.15658f
C1322 a_n3827_n3924.n19 gnd 0.676219f
C1323 a_n3827_n3924.n20 gnd 0.440278f
C1324 a_n3827_n3924.n21 gnd 0.844371f
C1325 a_n3827_n3924.t38 gnd 0.930864f
C1326 a_n3827_n3924.n22 gnd 0.578206f
C1327 a_n3827_n3924.t32 gnd 0.089565f
C1328 a_n3827_n3924.t36 gnd 0.089565f
C1329 a_n3827_n3924.n23 gnd 0.731493f
C1330 a_n3827_n3924.n24 gnd 0.368633f
C1331 a_n3827_n3924.t37 gnd 0.089565f
C1332 a_n3827_n3924.t25 gnd 0.089565f
C1333 a_n3827_n3924.n25 gnd 0.731493f
C1334 a_n3827_n3924.n26 gnd 0.368633f
C1335 a_n3827_n3924.t26 gnd 0.089565f
C1336 a_n3827_n3924.t20 gnd 0.089565f
C1337 a_n3827_n3924.n27 gnd 0.731493f
C1338 a_n3827_n3924.n28 gnd 0.368633f
C1339 a_n3827_n3924.t22 gnd 0.089565f
C1340 a_n3827_n3924.t35 gnd 0.089565f
C1341 a_n3827_n3924.n29 gnd 0.731493f
C1342 a_n3827_n3924.n30 gnd 0.368633f
C1343 a_n3827_n3924.t30 gnd 0.930864f
C1344 a_n3827_n3924.n31 gnd 0.351913f
C1345 a_n3827_n3924.t13 gnd 0.930864f
C1346 a_n3827_n3924.n32 gnd 0.351913f
C1347 a_n3827_n3924.t46 gnd 0.089565f
C1348 a_n3827_n3924.t11 gnd 0.089565f
C1349 a_n3827_n3924.n33 gnd 0.731493f
C1350 a_n3827_n3924.n34 gnd 0.368633f
C1351 a_n3827_n3924.t16 gnd 0.089565f
C1352 a_n3827_n3924.t40 gnd 0.089565f
C1353 a_n3827_n3924.n35 gnd 0.731493f
C1354 a_n3827_n3924.n36 gnd 0.368633f
C1355 a_n3827_n3924.t3 gnd 0.089565f
C1356 a_n3827_n3924.t45 gnd 0.089565f
C1357 a_n3827_n3924.n37 gnd 0.731493f
C1358 a_n3827_n3924.n38 gnd 0.368633f
C1359 a_n3827_n3924.t41 gnd 0.089565f
C1360 a_n3827_n3924.t18 gnd 0.089565f
C1361 a_n3827_n3924.n39 gnd 0.731493f
C1362 a_n3827_n3924.n40 gnd 0.368633f
C1363 a_n3827_n3924.t43 gnd 0.930864f
C1364 a_n3827_n3924.n41 gnd 0.578206f
C1365 a_n3827_n3924.n42 gnd 0.844371f
C1366 a_n3827_n3924.t21 gnd 0.930864f
C1367 a_n3827_n3924.n43 gnd 0.871367f
C1368 a_n3827_n3924.t29 gnd 0.089565f
C1369 a_n3827_n3924.t34 gnd 0.089565f
C1370 a_n3827_n3924.n44 gnd 0.731494f
C1371 a_n3827_n3924.n45 gnd 0.368632f
C1372 a_n3827_n3924.t27 gnd 0.089565f
C1373 a_n3827_n3924.t31 gnd 0.089565f
C1374 a_n3827_n3924.n46 gnd 0.731494f
C1375 a_n3827_n3924.n47 gnd 0.368632f
C1376 a_n3827_n3924.t24 gnd 0.089565f
C1377 a_n3827_n3924.t28 gnd 0.089565f
C1378 a_n3827_n3924.n48 gnd 0.731494f
C1379 a_n3827_n3924.n49 gnd 0.368632f
C1380 a_n3827_n3924.n50 gnd 0.368631f
C1381 a_n3827_n3924.n51 gnd 0.731495f
C1382 a_n3827_n3924.t39 gnd 0.089565f
C1383 plus.n0 gnd 0.022316f
C1384 plus.t6 gnd 0.405822f
C1385 plus.t12 gnd 0.37524f
C1386 plus.n1 gnd 0.151764f
C1387 plus.n2 gnd 0.022316f
C1388 plus.t8 gnd 0.37524f
C1389 plus.n3 gnd 0.018483f
C1390 plus.n4 gnd 0.022316f
C1391 plus.t7 gnd 0.37524f
C1392 plus.t19 gnd 0.37524f
C1393 plus.n5 gnd 0.151764f
C1394 plus.n6 gnd 0.022316f
C1395 plus.t18 gnd 0.37524f
C1396 plus.n7 gnd 0.151764f
C1397 plus.n8 gnd 0.022316f
C1398 plus.t24 gnd 0.37524f
C1399 plus.n9 gnd 0.018483f
C1400 plus.n10 gnd 0.022316f
C1401 plus.t22 gnd 0.37524f
C1402 plus.t9 gnd 0.37524f
C1403 plus.n11 gnd 0.174522f
C1404 plus.t14 gnd 0.420545f
C1405 plus.n12 gnd 0.176756f
C1406 plus.n13 gnd 0.09525f
C1407 plus.n14 gnd 0.028177f
C1408 plus.n15 gnd 0.025671f
C1409 plus.n16 gnd 0.151764f
C1410 plus.n17 gnd 0.027388f
C1411 plus.n18 gnd 0.022316f
C1412 plus.n19 gnd 0.022316f
C1413 plus.n20 gnd 0.022316f
C1414 plus.n21 gnd 0.028929f
C1415 plus.n22 gnd 0.151764f
C1416 plus.n23 gnd 0.027341f
C1417 plus.n24 gnd 0.026506f
C1418 plus.n25 gnd 0.022316f
C1419 plus.n26 gnd 0.022316f
C1420 plus.n27 gnd 0.028389f
C1421 plus.n28 gnd 0.018024f
C1422 plus.n29 gnd 0.028389f
C1423 plus.n30 gnd 0.022316f
C1424 plus.n31 gnd 0.022316f
C1425 plus.n32 gnd 0.026506f
C1426 plus.n33 gnd 0.027341f
C1427 plus.n34 gnd 0.151764f
C1428 plus.n35 gnd 0.028929f
C1429 plus.n36 gnd 0.022316f
C1430 plus.n37 gnd 0.022316f
C1431 plus.n38 gnd 0.022316f
C1432 plus.n39 gnd 0.027388f
C1433 plus.n40 gnd 0.151764f
C1434 plus.n41 gnd 0.025671f
C1435 plus.n42 gnd 0.028177f
C1436 plus.n43 gnd 0.022316f
C1437 plus.n44 gnd 0.022316f
C1438 plus.n45 gnd 0.029122f
C1439 plus.n46 gnd 0.008643f
C1440 plus.n47 gnd 0.175992f
C1441 plus.n48 gnd 0.25608f
C1442 plus.n49 gnd 0.022316f
C1443 plus.t10 gnd 0.37524f
C1444 plus.n50 gnd 0.151764f
C1445 plus.n51 gnd 0.022316f
C1446 plus.t15 gnd 0.37524f
C1447 plus.n52 gnd 0.018483f
C1448 plus.n53 gnd 0.022316f
C1449 plus.t13 gnd 0.37524f
C1450 plus.t17 gnd 0.37524f
C1451 plus.n54 gnd 0.151764f
C1452 plus.n55 gnd 0.022316f
C1453 plus.t16 gnd 0.37524f
C1454 plus.n56 gnd 0.151764f
C1455 plus.n57 gnd 0.022316f
C1456 plus.t20 gnd 0.37524f
C1457 plus.n58 gnd 0.018483f
C1458 plus.n59 gnd 0.022316f
C1459 plus.t21 gnd 0.37524f
C1460 plus.t5 gnd 0.37524f
C1461 plus.n60 gnd 0.174522f
C1462 plus.t11 gnd 0.420545f
C1463 plus.n61 gnd 0.176756f
C1464 plus.n62 gnd 0.09525f
C1465 plus.n63 gnd 0.028177f
C1466 plus.n64 gnd 0.025671f
C1467 plus.n65 gnd 0.151764f
C1468 plus.n66 gnd 0.027388f
C1469 plus.n67 gnd 0.022316f
C1470 plus.n68 gnd 0.022316f
C1471 plus.n69 gnd 0.022316f
C1472 plus.n70 gnd 0.028929f
C1473 plus.n71 gnd 0.151764f
C1474 plus.n72 gnd 0.027341f
C1475 plus.n73 gnd 0.026506f
C1476 plus.n74 gnd 0.022316f
C1477 plus.n75 gnd 0.022316f
C1478 plus.n76 gnd 0.028389f
C1479 plus.n77 gnd 0.018024f
C1480 plus.n78 gnd 0.028389f
C1481 plus.n79 gnd 0.022316f
C1482 plus.n80 gnd 0.022316f
C1483 plus.n81 gnd 0.026506f
C1484 plus.n82 gnd 0.027341f
C1485 plus.n83 gnd 0.151764f
C1486 plus.n84 gnd 0.028929f
C1487 plus.n85 gnd 0.022316f
C1488 plus.n86 gnd 0.022316f
C1489 plus.n87 gnd 0.022316f
C1490 plus.n88 gnd 0.027388f
C1491 plus.n89 gnd 0.151764f
C1492 plus.n90 gnd 0.025671f
C1493 plus.n91 gnd 0.028177f
C1494 plus.n92 gnd 0.022316f
C1495 plus.n93 gnd 0.022316f
C1496 plus.n94 gnd 0.029122f
C1497 plus.n95 gnd 0.008643f
C1498 plus.t23 gnd 0.405822f
C1499 plus.n96 gnd 0.175992f
C1500 plus.n97 gnd 0.745335f
C1501 plus.n98 gnd 1.11209f
C1502 plus.t1 gnd 0.038524f
C1503 plus.t3 gnd 0.006879f
C1504 plus.t2 gnd 0.006879f
C1505 plus.n99 gnd 0.022311f
C1506 plus.n100 gnd 0.173202f
C1507 plus.t4 gnd 0.006879f
C1508 plus.t0 gnd 0.006879f
C1509 plus.n101 gnd 0.022311f
C1510 plus.n102 gnd 0.130009f
C1511 plus.n103 gnd 2.81918f
C1512 a_n2472_13878.t25 gnd 0.187389f
C1513 a_n2472_13878.t21 gnd 0.187389f
C1514 a_n2472_13878.t27 gnd 0.187389f
C1515 a_n2472_13878.n0 gnd 1.47796f
C1516 a_n2472_13878.t8 gnd 0.187389f
C1517 a_n2472_13878.t18 gnd 0.187389f
C1518 a_n2472_13878.n1 gnd 1.47552f
C1519 a_n2472_13878.n2 gnd 1.32632f
C1520 a_n2472_13878.t23 gnd 0.187389f
C1521 a_n2472_13878.t15 gnd 0.187389f
C1522 a_n2472_13878.n3 gnd 1.47709f
C1523 a_n2472_13878.t20 gnd 0.187389f
C1524 a_n2472_13878.t14 gnd 0.187389f
C1525 a_n2472_13878.n4 gnd 1.47552f
C1526 a_n2472_13878.n5 gnd 2.06176f
C1527 a_n2472_13878.t10 gnd 0.187389f
C1528 a_n2472_13878.t12 gnd 0.187389f
C1529 a_n2472_13878.n6 gnd 1.47552f
C1530 a_n2472_13878.n7 gnd 1.00568f
C1531 a_n2472_13878.t22 gnd 0.187389f
C1532 a_n2472_13878.t11 gnd 0.187389f
C1533 a_n2472_13878.n8 gnd 1.47552f
C1534 a_n2472_13878.n9 gnd 1.00568f
C1535 a_n2472_13878.t19 gnd 0.187389f
C1536 a_n2472_13878.t9 gnd 0.187389f
C1537 a_n2472_13878.n10 gnd 1.47552f
C1538 a_n2472_13878.n11 gnd 4.40118f
C1539 a_n2472_13878.t1 gnd 1.75461f
C1540 a_n2472_13878.t4 gnd 0.187389f
C1541 a_n2472_13878.t5 gnd 0.187389f
C1542 a_n2472_13878.n12 gnd 1.31997f
C1543 a_n2472_13878.n13 gnd 1.47487f
C1544 a_n2472_13878.t0 gnd 1.75112f
C1545 a_n2472_13878.n14 gnd 0.742173f
C1546 a_n2472_13878.t3 gnd 1.75112f
C1547 a_n2472_13878.n15 gnd 0.742173f
C1548 a_n2472_13878.t6 gnd 0.187389f
C1549 a_n2472_13878.t7 gnd 0.187389f
C1550 a_n2472_13878.n16 gnd 1.31997f
C1551 a_n2472_13878.n17 gnd 0.749361f
C1552 a_n2472_13878.t2 gnd 1.75112f
C1553 a_n2472_13878.n18 gnd 2.43496f
C1554 a_n2472_13878.n19 gnd 3.22551f
C1555 a_n2472_13878.t24 gnd 0.187389f
C1556 a_n2472_13878.t13 gnd 0.187389f
C1557 a_n2472_13878.n20 gnd 1.47552f
C1558 a_n2472_13878.n21 gnd 2.21835f
C1559 a_n2472_13878.t16 gnd 0.187389f
C1560 a_n2472_13878.t17 gnd 0.187389f
C1561 a_n2472_13878.n22 gnd 1.47552f
C1562 a_n2472_13878.n23 gnd 0.653766f
C1563 a_n2472_13878.n24 gnd 0.653763f
C1564 a_n2472_13878.n25 gnd 1.47553f
C1565 a_n2472_13878.t26 gnd 0.187389f
C1566 a_n2650_13878.n0 gnd 0.89022f
C1567 a_n2650_13878.n1 gnd 3.61027f
C1568 a_n2650_13878.n2 gnd 3.33797f
C1569 a_n2650_13878.n3 gnd 3.94237f
C1570 a_n2650_13878.n4 gnd 0.783099f
C1571 a_n2650_13878.n5 gnd 0.199822f
C1572 a_n2650_13878.n6 gnd 0.147172f
C1573 a_n2650_13878.n7 gnd 0.231308f
C1574 a_n2650_13878.n8 gnd 0.178659f
C1575 a_n2650_13878.n9 gnd 0.199822f
C1576 a_n2650_13878.n10 gnd 0.147172f
C1577 a_n2650_13878.n11 gnd 0.835748f
C1578 a_n2650_13878.n12 gnd 0.210597f
C1579 a_n2650_13878.n13 gnd 0.679581f
C1580 a_n2650_13878.n14 gnd 0.210597f
C1581 a_n2650_13878.n15 gnd 0.490668f
C1582 a_n2650_13878.n16 gnd 0.210597f
C1583 a_n2650_13878.n17 gnd 0.543317f
C1584 a_n2650_13878.n18 gnd 0.210597f
C1585 a_n2650_13878.n19 gnd 0.871815f
C1586 a_n2650_13878.n20 gnd 0.210597f
C1587 a_n2650_13878.n21 gnd 2.91769f
C1588 a_n2650_13878.n22 gnd 0.783179f
C1589 a_n2650_13878.n23 gnd 0.210597f
C1590 a_n2650_13878.n24 gnd 0.911906f
C1591 a_n2650_13878.n25 gnd 0.210597f
C1592 a_n2650_13878.n26 gnd 0.490668f
C1593 a_n2650_13878.n27 gnd 1.73382f
C1594 a_n2650_13878.n28 gnd 1.16828f
C1595 a_n2650_13878.n29 gnd 2.18252f
C1596 a_n2650_13878.n30 gnd 1.14968f
C1597 a_n2650_13878.n31 gnd 1.16827f
C1598 a_n2650_13878.n32 gnd 0.438019f
C1599 a_n2650_13878.n33 gnd 0.278198f
C1600 a_n2650_13878.n34 gnd 0.00845f
C1601 a_n2650_13878.n35 gnd 4.07e-19
C1602 a_n2650_13878.n37 gnd 0.008154f
C1603 a_n2650_13878.n38 gnd 0.011856f
C1604 a_n2650_13878.n39 gnd 0.007844f
C1605 a_n2650_13878.n40 gnd 1.53361f
C1606 a_n2650_13878.n41 gnd 0.278198f
C1607 a_n2650_13878.n42 gnd 0.00845f
C1608 a_n2650_13878.n43 gnd 4.07e-19
C1609 a_n2650_13878.n45 gnd 0.008154f
C1610 a_n2650_13878.n46 gnd 0.011856f
C1611 a_n2650_13878.n47 gnd 0.00845f
C1612 a_n2650_13878.n48 gnd 4.07e-19
C1613 a_n2650_13878.n50 gnd 0.008154f
C1614 a_n2650_13878.n51 gnd 0.011856f
C1615 a_n2650_13878.n52 gnd 0.007844f
C1616 a_n2650_13878.n53 gnd 0.278198f
C1617 a_n2650_13878.n54 gnd 0.00845f
C1618 a_n2650_13878.n55 gnd 4.07e-19
C1619 a_n2650_13878.n57 gnd 0.008154f
C1620 a_n2650_13878.n58 gnd 0.011856f
C1621 a_n2650_13878.n59 gnd 0.007844f
C1622 a_n2650_13878.n60 gnd 0.278198f
C1623 a_n2650_13878.n61 gnd 0.008154f
C1624 a_n2650_13878.n62 gnd 0.278198f
C1625 a_n2650_13878.n63 gnd 0.008154f
C1626 a_n2650_13878.n64 gnd 0.278198f
C1627 a_n2650_13878.n65 gnd 0.008154f
C1628 a_n2650_13878.n66 gnd 0.278198f
C1629 a_n2650_13878.n67 gnd 0.008154f
C1630 a_n2650_13878.n68 gnd 0.278198f
C1631 a_n2650_13878.n69 gnd 0.007844f
C1632 a_n2650_13878.t36 gnd 0.146072f
C1633 a_n2650_13878.t30 gnd 1.36775f
C1634 a_n2650_13878.t44 gnd 0.146072f
C1635 a_n2650_13878.t48 gnd 0.146072f
C1636 a_n2650_13878.n70 gnd 1.02893f
C1637 a_n2650_13878.t21 gnd 0.679457f
C1638 a_n2650_13878.n71 gnd 0.295192f
C1639 a_n2650_13878.t27 gnd 0.679457f
C1640 a_n2650_13878.t47 gnd 0.679457f
C1641 a_n2650_13878.n72 gnd 0.298598f
C1642 a_n2650_13878.t29 gnd 0.679457f
C1643 a_n2650_13878.t72 gnd 0.679457f
C1644 a_n2650_13878.n73 gnd 0.295192f
C1645 a_n2650_13878.t87 gnd 0.679457f
C1646 a_n2650_13878.t90 gnd 0.679457f
C1647 a_n2650_13878.n74 gnd 0.298598f
C1648 a_n2650_13878.t66 gnd 0.679457f
C1649 a_n2650_13878.t11 gnd 0.679457f
C1650 a_n2650_13878.t17 gnd 0.679457f
C1651 a_n2650_13878.t45 gnd 0.679457f
C1652 a_n2650_13878.n75 gnd 0.298598f
C1653 a_n2650_13878.t31 gnd 0.679457f
C1654 a_n2650_13878.t39 gnd 0.679457f
C1655 a_n2650_13878.t33 gnd 0.679457f
C1656 a_n2650_13878.n76 gnd 0.294939f
C1657 a_n2650_13878.t13 gnd 0.679457f
C1658 a_n2650_13878.t37 gnd 0.679457f
C1659 a_n2650_13878.t23 gnd 0.679457f
C1660 a_n2650_13878.n77 gnd 0.298717f
C1661 a_n2650_13878.t8 gnd 0.113612f
C1662 a_n2650_13878.t57 gnd 0.113612f
C1663 a_n2650_13878.n78 gnd 1.00687f
C1664 a_n2650_13878.t7 gnd 0.113612f
C1665 a_n2650_13878.t49 gnd 0.113612f
C1666 a_n2650_13878.n79 gnd 1.00391f
C1667 a_n2650_13878.t52 gnd 0.113612f
C1668 a_n2650_13878.t3 gnd 0.113612f
C1669 a_n2650_13878.n80 gnd 1.00391f
C1670 a_n2650_13878.t50 gnd 0.113612f
C1671 a_n2650_13878.t54 gnd 0.113612f
C1672 a_n2650_13878.n81 gnd 1.00687f
C1673 a_n2650_13878.t56 gnd 0.113612f
C1674 a_n2650_13878.t53 gnd 0.113612f
C1675 a_n2650_13878.n82 gnd 1.00391f
C1676 a_n2650_13878.t55 gnd 0.113612f
C1677 a_n2650_13878.t59 gnd 0.113612f
C1678 a_n2650_13878.n83 gnd 1.00391f
C1679 a_n2650_13878.t58 gnd 0.113612f
C1680 a_n2650_13878.t1 gnd 0.113612f
C1681 a_n2650_13878.n84 gnd 1.00391f
C1682 a_n2650_13878.t4 gnd 0.113612f
C1683 a_n2650_13878.t0 gnd 0.113612f
C1684 a_n2650_13878.n85 gnd 1.00391f
C1685 a_n2650_13878.t5 gnd 0.113612f
C1686 a_n2650_13878.t2 gnd 0.113612f
C1687 a_n2650_13878.n86 gnd 1.00687f
C1688 a_n2650_13878.t51 gnd 0.113612f
C1689 a_n2650_13878.t6 gnd 0.113612f
C1690 a_n2650_13878.n87 gnd 1.00391f
C1691 a_n2650_13878.t94 gnd 0.679457f
C1692 a_n2650_13878.t73 gnd 0.679457f
C1693 a_n2650_13878.t78 gnd 0.679457f
C1694 a_n2650_13878.n88 gnd 0.298598f
C1695 a_n2650_13878.t67 gnd 0.679457f
C1696 a_n2650_13878.t83 gnd 0.679457f
C1697 a_n2650_13878.t91 gnd 0.679457f
C1698 a_n2650_13878.n89 gnd 0.294939f
C1699 a_n2650_13878.t92 gnd 0.679457f
C1700 a_n2650_13878.t62 gnd 0.679457f
C1701 a_n2650_13878.t75 gnd 0.679457f
C1702 a_n2650_13878.n90 gnd 0.298717f
C1703 a_n2650_13878.t65 gnd 0.690842f
C1704 a_n2650_13878.n91 gnd 0.295192f
C1705 a_n2650_13878.n92 gnd 0.289745f
C1706 a_n2650_13878.n93 gnd 0.298732f
C1707 a_n2650_13878.n94 gnd 0.301285f
C1708 a_n2650_13878.n95 gnd 0.294614f
C1709 a_n2650_13878.n96 gnd 0.289583f
C1710 a_n2650_13878.t25 gnd 0.690842f
C1711 a_n2650_13878.n97 gnd 0.295192f
C1712 a_n2650_13878.n98 gnd 0.289745f
C1713 a_n2650_13878.n99 gnd 0.298732f
C1714 a_n2650_13878.n100 gnd 0.301285f
C1715 a_n2650_13878.n101 gnd 0.294614f
C1716 a_n2650_13878.n102 gnd 0.289583f
C1717 a_n2650_13878.t26 gnd 1.36775f
C1718 a_n2650_13878.t38 gnd 0.146072f
C1719 a_n2650_13878.t24 gnd 0.146072f
C1720 a_n2650_13878.n103 gnd 1.02893f
C1721 a_n2650_13878.t34 gnd 0.146072f
C1722 a_n2650_13878.t14 gnd 0.146072f
C1723 a_n2650_13878.n104 gnd 1.02893f
C1724 a_n2650_13878.t32 gnd 0.146072f
C1725 a_n2650_13878.t40 gnd 0.146072f
C1726 a_n2650_13878.n105 gnd 1.02893f
C1727 a_n2650_13878.t18 gnd 0.146072f
C1728 a_n2650_13878.t46 gnd 0.146072f
C1729 a_n2650_13878.n106 gnd 1.02893f
C1730 a_n2650_13878.t12 gnd 1.36502f
C1731 a_n2650_13878.n107 gnd 1.41042f
C1732 a_n2650_13878.n108 gnd 0.918226f
C1733 a_n2650_13878.t71 gnd 0.679457f
C1734 a_n2650_13878.t81 gnd 0.679457f
C1735 a_n2650_13878.t95 gnd 0.679457f
C1736 a_n2650_13878.n109 gnd 0.298732f
C1737 a_n2650_13878.t84 gnd 0.679457f
C1738 a_n2650_13878.t68 gnd 0.679457f
C1739 a_n2650_13878.t69 gnd 0.679457f
C1740 a_n2650_13878.n110 gnd 0.298732f
C1741 a_n2650_13878.t88 gnd 0.679457f
C1742 a_n2650_13878.t77 gnd 0.679457f
C1743 a_n2650_13878.t76 gnd 0.679457f
C1744 a_n2650_13878.n111 gnd 0.298732f
C1745 a_n2650_13878.t80 gnd 0.679457f
C1746 a_n2650_13878.t70 gnd 0.679457f
C1747 a_n2650_13878.t60 gnd 0.679457f
C1748 a_n2650_13878.n112 gnd 0.298732f
C1749 a_n2650_13878.t85 gnd 0.690842f
C1750 a_n2650_13878.n113 gnd 0.294939f
C1751 a_n2650_13878.n114 gnd 0.289583f
C1752 a_n2650_13878.t93 gnd 0.690842f
C1753 a_n2650_13878.n115 gnd 0.294939f
C1754 a_n2650_13878.n116 gnd 0.289583f
C1755 a_n2650_13878.t79 gnd 0.690842f
C1756 a_n2650_13878.n117 gnd 0.294939f
C1757 a_n2650_13878.n118 gnd 0.289583f
C1758 a_n2650_13878.t74 gnd 0.690842f
C1759 a_n2650_13878.n119 gnd 0.294939f
C1760 a_n2650_13878.n120 gnd 0.289583f
C1761 a_n2650_13878.n121 gnd 1.20992f
C1762 a_n2650_13878.n122 gnd 0.289583f
C1763 a_n2650_13878.t89 gnd 0.679457f
C1764 a_n2650_13878.n123 gnd 0.294614f
C1765 a_n2650_13878.t64 gnd 0.679457f
C1766 a_n2650_13878.n124 gnd 0.301285f
C1767 a_n2650_13878.t86 gnd 0.679457f
C1768 a_n2650_13878.n125 gnd 0.298732f
C1769 a_n2650_13878.n126 gnd 0.294939f
C1770 a_n2650_13878.t61 gnd 0.679457f
C1771 a_n2650_13878.n127 gnd 0.289745f
C1772 a_n2650_13878.t82 gnd 0.679457f
C1773 a_n2650_13878.n128 gnd 0.298717f
C1774 a_n2650_13878.t63 gnd 0.690842f
C1775 a_n2650_13878.n129 gnd 0.289583f
C1776 a_n2650_13878.t43 gnd 0.679457f
C1777 a_n2650_13878.n130 gnd 0.294614f
C1778 a_n2650_13878.t35 gnd 0.679457f
C1779 a_n2650_13878.n131 gnd 0.301285f
C1780 a_n2650_13878.t9 gnd 0.679457f
C1781 a_n2650_13878.n132 gnd 0.298732f
C1782 a_n2650_13878.n133 gnd 0.294939f
C1783 a_n2650_13878.t15 gnd 0.679457f
C1784 a_n2650_13878.n134 gnd 0.289745f
C1785 a_n2650_13878.t41 gnd 0.679457f
C1786 a_n2650_13878.n135 gnd 0.298717f
C1787 a_n2650_13878.t19 gnd 0.690842f
C1788 a_n2650_13878.n136 gnd 1.24181f
C1789 a_n2650_13878.t20 gnd 1.36502f
C1790 a_n2650_13878.t22 gnd 0.146072f
C1791 a_n2650_13878.t42 gnd 0.146072f
C1792 a_n2650_13878.n137 gnd 1.02893f
C1793 a_n2650_13878.t28 gnd 0.146072f
C1794 a_n2650_13878.t16 gnd 0.146072f
C1795 a_n2650_13878.n138 gnd 1.02893f
C1796 a_n2650_13878.n139 gnd 1.02894f
C1797 a_n2650_13878.t10 gnd 0.146072f
C1798 CSoutput.n0 gnd 0.048277f
C1799 CSoutput.t197 gnd 0.319339f
C1800 CSoutput.n1 gnd 0.144197f
C1801 CSoutput.n2 gnd 0.048277f
C1802 CSoutput.t203 gnd 0.319339f
C1803 CSoutput.n3 gnd 0.038263f
C1804 CSoutput.n4 gnd 0.048277f
C1805 CSoutput.t192 gnd 0.319339f
C1806 CSoutput.n5 gnd 0.032995f
C1807 CSoutput.n6 gnd 0.048277f
C1808 CSoutput.t200 gnd 0.319339f
C1809 CSoutput.t184 gnd 0.319339f
C1810 CSoutput.n7 gnd 0.142626f
C1811 CSoutput.n8 gnd 0.048277f
C1812 CSoutput.t205 gnd 0.319339f
C1813 CSoutput.n9 gnd 0.031459f
C1814 CSoutput.n10 gnd 0.048277f
C1815 CSoutput.t193 gnd 0.319339f
C1816 CSoutput.t204 gnd 0.319339f
C1817 CSoutput.n11 gnd 0.142626f
C1818 CSoutput.n12 gnd 0.048277f
C1819 CSoutput.t201 gnd 0.319339f
C1820 CSoutput.n13 gnd 0.032995f
C1821 CSoutput.n14 gnd 0.048277f
C1822 CSoutput.t191 gnd 0.319339f
C1823 CSoutput.t194 gnd 0.319339f
C1824 CSoutput.n15 gnd 0.142626f
C1825 CSoutput.n16 gnd 0.048277f
C1826 CSoutput.t198 gnd 0.319339f
C1827 CSoutput.n17 gnd 0.03524f
C1828 CSoutput.t188 gnd 0.381619f
C1829 CSoutput.t190 gnd 0.319339f
C1830 CSoutput.n18 gnd 0.182078f
C1831 CSoutput.n19 gnd 0.176679f
C1832 CSoutput.n20 gnd 0.204968f
C1833 CSoutput.n21 gnd 0.048277f
C1834 CSoutput.n22 gnd 0.040292f
C1835 CSoutput.n23 gnd 0.142626f
C1836 CSoutput.n24 gnd 0.03884f
C1837 CSoutput.n25 gnd 0.038263f
C1838 CSoutput.n26 gnd 0.048277f
C1839 CSoutput.n27 gnd 0.048277f
C1840 CSoutput.n28 gnd 0.039982f
C1841 CSoutput.n29 gnd 0.033946f
C1842 CSoutput.n30 gnd 0.145801f
C1843 CSoutput.n31 gnd 0.034414f
C1844 CSoutput.n32 gnd 0.048277f
C1845 CSoutput.n33 gnd 0.048277f
C1846 CSoutput.n34 gnd 0.048277f
C1847 CSoutput.n35 gnd 0.039556f
C1848 CSoutput.n36 gnd 0.142626f
C1849 CSoutput.n37 gnd 0.03783f
C1850 CSoutput.n38 gnd 0.039274f
C1851 CSoutput.n39 gnd 0.048277f
C1852 CSoutput.n40 gnd 0.048277f
C1853 CSoutput.n41 gnd 0.040284f
C1854 CSoutput.n42 gnd 0.03682f
C1855 CSoutput.n43 gnd 0.142626f
C1856 CSoutput.n44 gnd 0.037753f
C1857 CSoutput.n45 gnd 0.048277f
C1858 CSoutput.n46 gnd 0.048277f
C1859 CSoutput.n47 gnd 0.048277f
C1860 CSoutput.n48 gnd 0.037753f
C1861 CSoutput.n49 gnd 0.142626f
C1862 CSoutput.n50 gnd 0.03682f
C1863 CSoutput.n51 gnd 0.040284f
C1864 CSoutput.n52 gnd 0.048277f
C1865 CSoutput.n53 gnd 0.048277f
C1866 CSoutput.n54 gnd 0.039274f
C1867 CSoutput.n55 gnd 0.03783f
C1868 CSoutput.n56 gnd 0.142626f
C1869 CSoutput.n57 gnd 0.039556f
C1870 CSoutput.n58 gnd 0.048277f
C1871 CSoutput.n59 gnd 0.048277f
C1872 CSoutput.n60 gnd 0.048277f
C1873 CSoutput.n61 gnd 0.034414f
C1874 CSoutput.n62 gnd 0.145801f
C1875 CSoutput.n63 gnd 0.033946f
C1876 CSoutput.t186 gnd 0.319339f
C1877 CSoutput.n64 gnd 0.142626f
C1878 CSoutput.n65 gnd 0.039982f
C1879 CSoutput.n66 gnd 0.048277f
C1880 CSoutput.n67 gnd 0.048277f
C1881 CSoutput.n68 gnd 0.048277f
C1882 CSoutput.n69 gnd 0.03884f
C1883 CSoutput.n70 gnd 0.142626f
C1884 CSoutput.n71 gnd 0.040292f
C1885 CSoutput.n72 gnd 0.03524f
C1886 CSoutput.n73 gnd 0.048277f
C1887 CSoutput.n74 gnd 0.048277f
C1888 CSoutput.n75 gnd 0.036546f
C1889 CSoutput.n76 gnd 0.021705f
C1890 CSoutput.t189 gnd 0.3588f
C1891 CSoutput.n77 gnd 0.178238f
C1892 CSoutput.n78 gnd 0.762662f
C1893 CSoutput.t60 gnd 0.060218f
C1894 CSoutput.t118 gnd 0.060218f
C1895 CSoutput.n79 gnd 0.46623f
C1896 CSoutput.t67 gnd 0.060218f
C1897 CSoutput.t93 gnd 0.060218f
C1898 CSoutput.n80 gnd 0.465398f
C1899 CSoutput.n81 gnd 0.472379f
C1900 CSoutput.t172 gnd 0.060218f
C1901 CSoutput.t111 gnd 0.060218f
C1902 CSoutput.n82 gnd 0.465398f
C1903 CSoutput.n83 gnd 0.232768f
C1904 CSoutput.t69 gnd 0.060218f
C1905 CSoutput.t151 gnd 0.060218f
C1906 CSoutput.n84 gnd 0.465398f
C1907 CSoutput.n85 gnd 0.232768f
C1908 CSoutput.t76 gnd 0.060218f
C1909 CSoutput.t133 gnd 0.060218f
C1910 CSoutput.n86 gnd 0.465398f
C1911 CSoutput.n87 gnd 0.232768f
C1912 CSoutput.t98 gnd 0.060218f
C1913 CSoutput.t119 gnd 0.060218f
C1914 CSoutput.n88 gnd 0.465398f
C1915 CSoutput.n89 gnd 0.232768f
C1916 CSoutput.t114 gnd 0.060218f
C1917 CSoutput.t160 gnd 0.060218f
C1918 CSoutput.n90 gnd 0.465398f
C1919 CSoutput.n91 gnd 0.232768f
C1920 CSoutput.t86 gnd 0.060218f
C1921 CSoutput.t138 gnd 0.060218f
C1922 CSoutput.n92 gnd 0.465398f
C1923 CSoutput.n93 gnd 0.232768f
C1924 CSoutput.t107 gnd 0.060218f
C1925 CSoutput.t153 gnd 0.060218f
C1926 CSoutput.n94 gnd 0.465398f
C1927 CSoutput.n95 gnd 0.232768f
C1928 CSoutput.t123 gnd 0.060218f
C1929 CSoutput.t168 gnd 0.060218f
C1930 CSoutput.n96 gnd 0.465398f
C1931 CSoutput.n97 gnd 0.426843f
C1932 CSoutput.t81 gnd 0.060218f
C1933 CSoutput.t161 gnd 0.060218f
C1934 CSoutput.n98 gnd 0.46623f
C1935 CSoutput.t131 gnd 0.060218f
C1936 CSoutput.t129 gnd 0.060218f
C1937 CSoutput.n99 gnd 0.465398f
C1938 CSoutput.n100 gnd 0.472379f
C1939 CSoutput.t115 gnd 0.060218f
C1940 CSoutput.t78 gnd 0.060218f
C1941 CSoutput.n101 gnd 0.465398f
C1942 CSoutput.n102 gnd 0.232768f
C1943 CSoutput.t59 gnd 0.060218f
C1944 CSoutput.t117 gnd 0.060218f
C1945 CSoutput.n103 gnd 0.465398f
C1946 CSoutput.n104 gnd 0.232768f
C1947 CSoutput.t112 gnd 0.060218f
C1948 CSoutput.t75 gnd 0.060218f
C1949 CSoutput.n105 gnd 0.465398f
C1950 CSoutput.n106 gnd 0.232768f
C1951 CSoutput.t57 gnd 0.060218f
C1952 CSoutput.t55 gnd 0.060218f
C1953 CSoutput.n107 gnd 0.465398f
C1954 CSoutput.n108 gnd 0.232768f
C1955 CSoutput.t134 gnd 0.060218f
C1956 CSoutput.t94 gnd 0.060218f
C1957 CSoutput.n109 gnd 0.465398f
C1958 CSoutput.n110 gnd 0.232768f
C1959 CSoutput.t88 gnd 0.060218f
C1960 CSoutput.t54 gnd 0.060218f
C1961 CSoutput.n111 gnd 0.465398f
C1962 CSoutput.n112 gnd 0.232768f
C1963 CSoutput.t157 gnd 0.060218f
C1964 CSoutput.t130 gnd 0.060218f
C1965 CSoutput.n113 gnd 0.465398f
C1966 CSoutput.n114 gnd 0.232768f
C1967 CSoutput.t116 gnd 0.060218f
C1968 CSoutput.t79 gnd 0.060218f
C1969 CSoutput.n115 gnd 0.465398f
C1970 CSoutput.n116 gnd 0.347116f
C1971 CSoutput.n117 gnd 0.437711f
C1972 CSoutput.t99 gnd 0.060218f
C1973 CSoutput.t173 gnd 0.060218f
C1974 CSoutput.n118 gnd 0.46623f
C1975 CSoutput.t142 gnd 0.060218f
C1976 CSoutput.t140 gnd 0.060218f
C1977 CSoutput.n119 gnd 0.465398f
C1978 CSoutput.n120 gnd 0.472379f
C1979 CSoutput.t125 gnd 0.060218f
C1980 CSoutput.t95 gnd 0.060218f
C1981 CSoutput.n121 gnd 0.465398f
C1982 CSoutput.n122 gnd 0.232768f
C1983 CSoutput.t72 gnd 0.060218f
C1984 CSoutput.t127 gnd 0.060218f
C1985 CSoutput.n123 gnd 0.465398f
C1986 CSoutput.n124 gnd 0.232768f
C1987 CSoutput.t124 gnd 0.060218f
C1988 CSoutput.t92 gnd 0.060218f
C1989 CSoutput.n125 gnd 0.465398f
C1990 CSoutput.n126 gnd 0.232768f
C1991 CSoutput.t71 gnd 0.060218f
C1992 CSoutput.t70 gnd 0.060218f
C1993 CSoutput.n127 gnd 0.465398f
C1994 CSoutput.n128 gnd 0.232768f
C1995 CSoutput.t143 gnd 0.060218f
C1996 CSoutput.t108 gnd 0.060218f
C1997 CSoutput.n129 gnd 0.465398f
C1998 CSoutput.n130 gnd 0.232768f
C1999 CSoutput.t103 gnd 0.060218f
C2000 CSoutput.t66 gnd 0.060218f
C2001 CSoutput.n131 gnd 0.465398f
C2002 CSoutput.n132 gnd 0.232768f
C2003 CSoutput.t169 gnd 0.060218f
C2004 CSoutput.t141 gnd 0.060218f
C2005 CSoutput.n133 gnd 0.465398f
C2006 CSoutput.n134 gnd 0.232768f
C2007 CSoutput.t126 gnd 0.060218f
C2008 CSoutput.t96 gnd 0.060218f
C2009 CSoutput.n135 gnd 0.465398f
C2010 CSoutput.n136 gnd 0.347116f
C2011 CSoutput.n137 gnd 0.489249f
C2012 CSoutput.n138 gnd 9.722839f
C2013 CSoutput.n140 gnd 0.854004f
C2014 CSoutput.n141 gnd 0.640503f
C2015 CSoutput.n142 gnd 0.854004f
C2016 CSoutput.n143 gnd 0.854004f
C2017 CSoutput.n144 gnd 2.29924f
C2018 CSoutput.n145 gnd 0.854004f
C2019 CSoutput.n146 gnd 0.854004f
C2020 CSoutput.t185 gnd 1.06751f
C2021 CSoutput.n147 gnd 0.854004f
C2022 CSoutput.n148 gnd 0.854004f
C2023 CSoutput.n152 gnd 0.854004f
C2024 CSoutput.n156 gnd 0.854004f
C2025 CSoutput.n157 gnd 0.854004f
C2026 CSoutput.n159 gnd 0.854004f
C2027 CSoutput.n164 gnd 0.854004f
C2028 CSoutput.n166 gnd 0.854004f
C2029 CSoutput.n167 gnd 0.854004f
C2030 CSoutput.n169 gnd 0.854004f
C2031 CSoutput.n170 gnd 0.854004f
C2032 CSoutput.n172 gnd 0.854004f
C2033 CSoutput.t196 gnd 14.2703f
C2034 CSoutput.n174 gnd 0.854004f
C2035 CSoutput.n175 gnd 0.640503f
C2036 CSoutput.n176 gnd 0.854004f
C2037 CSoutput.n177 gnd 0.854004f
C2038 CSoutput.n178 gnd 2.29924f
C2039 CSoutput.n179 gnd 0.854004f
C2040 CSoutput.n180 gnd 0.854004f
C2041 CSoutput.t199 gnd 1.06751f
C2042 CSoutput.n181 gnd 0.854004f
C2043 CSoutput.n182 gnd 0.854004f
C2044 CSoutput.n186 gnd 0.854004f
C2045 CSoutput.n190 gnd 0.854004f
C2046 CSoutput.n191 gnd 0.854004f
C2047 CSoutput.n193 gnd 0.854004f
C2048 CSoutput.n198 gnd 0.854004f
C2049 CSoutput.n200 gnd 0.854004f
C2050 CSoutput.n201 gnd 0.854004f
C2051 CSoutput.n203 gnd 0.854004f
C2052 CSoutput.n204 gnd 0.854004f
C2053 CSoutput.n206 gnd 0.854004f
C2054 CSoutput.n207 gnd 0.640503f
C2055 CSoutput.n209 gnd 0.854004f
C2056 CSoutput.n210 gnd 0.640503f
C2057 CSoutput.n211 gnd 0.854004f
C2058 CSoutput.n212 gnd 0.854004f
C2059 CSoutput.n213 gnd 2.29924f
C2060 CSoutput.n214 gnd 0.854004f
C2061 CSoutput.n215 gnd 0.854004f
C2062 CSoutput.t195 gnd 1.06751f
C2063 CSoutput.n216 gnd 0.854004f
C2064 CSoutput.n217 gnd 2.29924f
C2065 CSoutput.n219 gnd 0.854004f
C2066 CSoutput.n220 gnd 0.854004f
C2067 CSoutput.n222 gnd 0.854004f
C2068 CSoutput.n223 gnd 0.854004f
C2069 CSoutput.t202 gnd 14.0378f
C2070 CSoutput.t187 gnd 14.2703f
C2071 CSoutput.n229 gnd 2.67914f
C2072 CSoutput.n230 gnd 10.9138f
C2073 CSoutput.n231 gnd 11.3705f
C2074 CSoutput.n236 gnd 2.90223f
C2075 CSoutput.n242 gnd 0.854004f
C2076 CSoutput.n244 gnd 0.854004f
C2077 CSoutput.n246 gnd 0.854004f
C2078 CSoutput.n248 gnd 0.854004f
C2079 CSoutput.n250 gnd 0.854004f
C2080 CSoutput.n256 gnd 0.854004f
C2081 CSoutput.n263 gnd 1.56677f
C2082 CSoutput.n264 gnd 1.56677f
C2083 CSoutput.n265 gnd 0.854004f
C2084 CSoutput.n266 gnd 0.854004f
C2085 CSoutput.n268 gnd 0.640503f
C2086 CSoutput.n269 gnd 0.548533f
C2087 CSoutput.n271 gnd 0.640503f
C2088 CSoutput.n272 gnd 0.548533f
C2089 CSoutput.n273 gnd 0.640503f
C2090 CSoutput.n275 gnd 0.854004f
C2091 CSoutput.n277 gnd 2.29924f
C2092 CSoutput.n278 gnd 2.67914f
C2093 CSoutput.n279 gnd 10.0379f
C2094 CSoutput.n281 gnd 0.640503f
C2095 CSoutput.n282 gnd 1.64805f
C2096 CSoutput.n283 gnd 0.640503f
C2097 CSoutput.n285 gnd 0.854004f
C2098 CSoutput.n287 gnd 2.29924f
C2099 CSoutput.n288 gnd 5.00812f
C2100 CSoutput.t144 gnd 0.060218f
C2101 CSoutput.t58 gnd 0.060218f
C2102 CSoutput.n289 gnd 0.46623f
C2103 CSoutput.t91 gnd 0.060218f
C2104 CSoutput.t65 gnd 0.060218f
C2105 CSoutput.n290 gnd 0.465398f
C2106 CSoutput.n291 gnd 0.472379f
C2107 CSoutput.t110 gnd 0.060218f
C2108 CSoutput.t85 gnd 0.060218f
C2109 CSoutput.n292 gnd 0.465398f
C2110 CSoutput.n293 gnd 0.232768f
C2111 CSoutput.t150 gnd 0.060218f
C2112 CSoutput.t68 gnd 0.060218f
C2113 CSoutput.n294 gnd 0.465398f
C2114 CSoutput.n295 gnd 0.232768f
C2115 CSoutput.t132 gnd 0.060218f
C2116 CSoutput.t73 gnd 0.060218f
C2117 CSoutput.n296 gnd 0.465398f
C2118 CSoutput.n297 gnd 0.232768f
C2119 CSoutput.t146 gnd 0.060218f
C2120 CSoutput.t97 gnd 0.060218f
C2121 CSoutput.n298 gnd 0.465398f
C2122 CSoutput.n299 gnd 0.232768f
C2123 CSoutput.t159 gnd 0.060218f
C2124 CSoutput.t113 gnd 0.060218f
C2125 CSoutput.n300 gnd 0.465398f
C2126 CSoutput.n301 gnd 0.232768f
C2127 CSoutput.t137 gnd 0.060218f
C2128 CSoutput.t87 gnd 0.060218f
C2129 CSoutput.n302 gnd 0.465398f
C2130 CSoutput.n303 gnd 0.232768f
C2131 CSoutput.t152 gnd 0.060218f
C2132 CSoutput.t105 gnd 0.060218f
C2133 CSoutput.n304 gnd 0.465398f
C2134 CSoutput.n305 gnd 0.232768f
C2135 CSoutput.t167 gnd 0.060218f
C2136 CSoutput.t121 gnd 0.060218f
C2137 CSoutput.n306 gnd 0.465398f
C2138 CSoutput.n307 gnd 0.426843f
C2139 CSoutput.t90 gnd 0.060218f
C2140 CSoutput.t158 gnd 0.060218f
C2141 CSoutput.n308 gnd 0.46623f
C2142 CSoutput.t82 gnd 0.060218f
C2143 CSoutput.t84 gnd 0.060218f
C2144 CSoutput.n309 gnd 0.465398f
C2145 CSoutput.n310 gnd 0.472379f
C2146 CSoutput.t155 gnd 0.060218f
C2147 CSoutput.t156 gnd 0.060218f
C2148 CSoutput.n311 gnd 0.465398f
C2149 CSoutput.n312 gnd 0.232768f
C2150 CSoutput.t64 gnd 0.060218f
C2151 CSoutput.t139 gnd 0.060218f
C2152 CSoutput.n313 gnd 0.465398f
C2153 CSoutput.n314 gnd 0.232768f
C2154 CSoutput.t149 gnd 0.060218f
C2155 CSoutput.t61 gnd 0.060218f
C2156 CSoutput.n315 gnd 0.465398f
C2157 CSoutput.n316 gnd 0.232768f
C2158 CSoutput.t109 gnd 0.060218f
C2159 CSoutput.t136 gnd 0.060218f
C2160 CSoutput.n317 gnd 0.465398f
C2161 CSoutput.n318 gnd 0.232768f
C2162 CSoutput.t163 gnd 0.060218f
C2163 CSoutput.t89 gnd 0.060218f
C2164 CSoutput.n319 gnd 0.465398f
C2165 CSoutput.n320 gnd 0.232768f
C2166 CSoutput.t135 gnd 0.060218f
C2167 CSoutput.t171 gnd 0.060218f
C2168 CSoutput.n321 gnd 0.465398f
C2169 CSoutput.n322 gnd 0.232768f
C2170 CSoutput.t83 gnd 0.060218f
C2171 CSoutput.t120 gnd 0.060218f
C2172 CSoutput.n323 gnd 0.465398f
C2173 CSoutput.n324 gnd 0.232768f
C2174 CSoutput.t154 gnd 0.060218f
C2175 CSoutput.t63 gnd 0.060218f
C2176 CSoutput.n325 gnd 0.465398f
C2177 CSoutput.n326 gnd 0.347116f
C2178 CSoutput.n327 gnd 0.437711f
C2179 CSoutput.t106 gnd 0.060218f
C2180 CSoutput.t170 gnd 0.060218f
C2181 CSoutput.n328 gnd 0.46623f
C2182 CSoutput.t100 gnd 0.060218f
C2183 CSoutput.t102 gnd 0.060218f
C2184 CSoutput.n329 gnd 0.465398f
C2185 CSoutput.n330 gnd 0.472379f
C2186 CSoutput.t164 gnd 0.060218f
C2187 CSoutput.t166 gnd 0.060218f
C2188 CSoutput.n331 gnd 0.465398f
C2189 CSoutput.n332 gnd 0.232768f
C2190 CSoutput.t80 gnd 0.060218f
C2191 CSoutput.t148 gnd 0.060218f
C2192 CSoutput.n333 gnd 0.465398f
C2193 CSoutput.n334 gnd 0.232768f
C2194 CSoutput.t162 gnd 0.060218f
C2195 CSoutput.t74 gnd 0.060218f
C2196 CSoutput.n335 gnd 0.465398f
C2197 CSoutput.n336 gnd 0.232768f
C2198 CSoutput.t122 gnd 0.060218f
C2199 CSoutput.t147 gnd 0.060218f
C2200 CSoutput.n337 gnd 0.465398f
C2201 CSoutput.n338 gnd 0.232768f
C2202 CSoutput.t56 gnd 0.060218f
C2203 CSoutput.t104 gnd 0.060218f
C2204 CSoutput.n339 gnd 0.465398f
C2205 CSoutput.n340 gnd 0.232768f
C2206 CSoutput.t145 gnd 0.060218f
C2207 CSoutput.t62 gnd 0.060218f
C2208 CSoutput.n341 gnd 0.465398f
C2209 CSoutput.n342 gnd 0.232768f
C2210 CSoutput.t101 gnd 0.060218f
C2211 CSoutput.t128 gnd 0.060218f
C2212 CSoutput.n343 gnd 0.465398f
C2213 CSoutput.n344 gnd 0.232768f
C2214 CSoutput.t165 gnd 0.060218f
C2215 CSoutput.t77 gnd 0.060218f
C2216 CSoutput.n345 gnd 0.465397f
C2217 CSoutput.n346 gnd 0.347118f
C2218 CSoutput.n347 gnd 0.489249f
C2219 CSoutput.n348 gnd 13.6148f
C2220 CSoutput.t4 gnd 0.052691f
C2221 CSoutput.t23 gnd 0.052691f
C2222 CSoutput.n349 gnd 0.467154f
C2223 CSoutput.t176 gnd 0.052691f
C2224 CSoutput.t16 gnd 0.052691f
C2225 CSoutput.n350 gnd 0.465596f
C2226 CSoutput.n351 gnd 0.433848f
C2227 CSoutput.t0 gnd 0.052691f
C2228 CSoutput.t180 gnd 0.052691f
C2229 CSoutput.n352 gnd 0.465596f
C2230 CSoutput.n353 gnd 0.213867f
C2231 CSoutput.t51 gnd 0.052691f
C2232 CSoutput.t19 gnd 0.052691f
C2233 CSoutput.n354 gnd 0.465596f
C2234 CSoutput.n355 gnd 0.213867f
C2235 CSoutput.t35 gnd 0.052691f
C2236 CSoutput.t175 gnd 0.052691f
C2237 CSoutput.n356 gnd 0.465596f
C2238 CSoutput.n357 gnd 0.213867f
C2239 CSoutput.t45 gnd 0.052691f
C2240 CSoutput.t5 gnd 0.052691f
C2241 CSoutput.n358 gnd 0.465596f
C2242 CSoutput.n359 gnd 0.213867f
C2243 CSoutput.t53 gnd 0.052691f
C2244 CSoutput.t37 gnd 0.052691f
C2245 CSoutput.n360 gnd 0.465596f
C2246 CSoutput.n361 gnd 0.213867f
C2247 CSoutput.t1 gnd 0.052691f
C2248 CSoutput.t41 gnd 0.052691f
C2249 CSoutput.n362 gnd 0.465596f
C2250 CSoutput.n363 gnd 0.394414f
C2251 CSoutput.t17 gnd 0.052691f
C2252 CSoutput.t24 gnd 0.052691f
C2253 CSoutput.n364 gnd 0.467154f
C2254 CSoutput.t29 gnd 0.052691f
C2255 CSoutput.t20 gnd 0.052691f
C2256 CSoutput.n365 gnd 0.465596f
C2257 CSoutput.n366 gnd 0.433848f
C2258 CSoutput.t181 gnd 0.052691f
C2259 CSoutput.t52 gnd 0.052691f
C2260 CSoutput.n367 gnd 0.465596f
C2261 CSoutput.n368 gnd 0.213867f
C2262 CSoutput.t21 gnd 0.052691f
C2263 CSoutput.t22 gnd 0.052691f
C2264 CSoutput.n369 gnd 0.465596f
C2265 CSoutput.n370 gnd 0.213867f
C2266 CSoutput.t36 gnd 0.052691f
C2267 CSoutput.t38 gnd 0.052691f
C2268 CSoutput.n371 gnd 0.465596f
C2269 CSoutput.n372 gnd 0.213867f
C2270 CSoutput.t7 gnd 0.052691f
C2271 CSoutput.t49 gnd 0.052691f
C2272 CSoutput.n373 gnd 0.465596f
C2273 CSoutput.n374 gnd 0.213867f
C2274 CSoutput.t42 gnd 0.052691f
C2275 CSoutput.t40 gnd 0.052691f
C2276 CSoutput.n375 gnd 0.465596f
C2277 CSoutput.n376 gnd 0.213867f
C2278 CSoutput.t43 gnd 0.052691f
C2279 CSoutput.t31 gnd 0.052691f
C2280 CSoutput.n377 gnd 0.465596f
C2281 CSoutput.n378 gnd 0.324696f
C2282 CSoutput.n379 gnd 0.603309f
C2283 CSoutput.n380 gnd 13.9433f
C2284 CSoutput.t9 gnd 0.052691f
C2285 CSoutput.t28 gnd 0.052691f
C2286 CSoutput.n381 gnd 0.467154f
C2287 CSoutput.t30 gnd 0.052691f
C2288 CSoutput.t46 gnd 0.052691f
C2289 CSoutput.n382 gnd 0.465596f
C2290 CSoutput.n383 gnd 0.433848f
C2291 CSoutput.t47 gnd 0.052691f
C2292 CSoutput.t174 gnd 0.052691f
C2293 CSoutput.n384 gnd 0.465596f
C2294 CSoutput.n385 gnd 0.213867f
C2295 CSoutput.t15 gnd 0.052691f
C2296 CSoutput.t44 gnd 0.052691f
C2297 CSoutput.n386 gnd 0.465596f
C2298 CSoutput.n387 gnd 0.213867f
C2299 CSoutput.t11 gnd 0.052691f
C2300 CSoutput.t14 gnd 0.052691f
C2301 CSoutput.n388 gnd 0.465596f
C2302 CSoutput.n389 gnd 0.213867f
C2303 CSoutput.t178 gnd 0.052691f
C2304 CSoutput.t33 gnd 0.052691f
C2305 CSoutput.n390 gnd 0.465596f
C2306 CSoutput.n391 gnd 0.213867f
C2307 CSoutput.t12 gnd 0.052691f
C2308 CSoutput.t25 gnd 0.052691f
C2309 CSoutput.n392 gnd 0.465596f
C2310 CSoutput.n393 gnd 0.213867f
C2311 CSoutput.t183 gnd 0.052691f
C2312 CSoutput.t50 gnd 0.052691f
C2313 CSoutput.n394 gnd 0.465596f
C2314 CSoutput.n395 gnd 0.394414f
C2315 CSoutput.t26 gnd 0.052691f
C2316 CSoutput.t2 gnd 0.052691f
C2317 CSoutput.n396 gnd 0.467154f
C2318 CSoutput.t6 gnd 0.052691f
C2319 CSoutput.t13 gnd 0.052691f
C2320 CSoutput.n397 gnd 0.465596f
C2321 CSoutput.n398 gnd 0.433848f
C2322 CSoutput.t177 gnd 0.052691f
C2323 CSoutput.t3 gnd 0.052691f
C2324 CSoutput.n399 gnd 0.465596f
C2325 CSoutput.n400 gnd 0.213867f
C2326 CSoutput.t18 gnd 0.052691f
C2327 CSoutput.t48 gnd 0.052691f
C2328 CSoutput.n401 gnd 0.465596f
C2329 CSoutput.n402 gnd 0.213867f
C2330 CSoutput.t8 gnd 0.052691f
C2331 CSoutput.t27 gnd 0.052691f
C2332 CSoutput.n403 gnd 0.465596f
C2333 CSoutput.n404 gnd 0.213867f
C2334 CSoutput.t182 gnd 0.052691f
C2335 CSoutput.t34 gnd 0.052691f
C2336 CSoutput.n405 gnd 0.465596f
C2337 CSoutput.n406 gnd 0.213867f
C2338 CSoutput.t179 gnd 0.052691f
C2339 CSoutput.t39 gnd 0.052691f
C2340 CSoutput.n407 gnd 0.465596f
C2341 CSoutput.n408 gnd 0.213867f
C2342 CSoutput.t10 gnd 0.052691f
C2343 CSoutput.t32 gnd 0.052691f
C2344 CSoutput.n409 gnd 0.465596f
C2345 CSoutput.n410 gnd 0.324696f
C2346 CSoutput.n411 gnd 0.603309f
C2347 CSoutput.n412 gnd 8.38815f
C2348 CSoutput.n413 gnd 15.4765f
C2349 vdd.t110 gnd 0.037975f
C2350 vdd.t104 gnd 0.037975f
C2351 vdd.n0 gnd 0.299515f
C2352 vdd.t2 gnd 0.037975f
C2353 vdd.t303 gnd 0.037975f
C2354 vdd.n1 gnd 0.29902f
C2355 vdd.n2 gnd 0.275754f
C2356 vdd.t119 gnd 0.037975f
C2357 vdd.t138 gnd 0.037975f
C2358 vdd.n3 gnd 0.29902f
C2359 vdd.n4 gnd 0.139459f
C2360 vdd.t140 gnd 0.037975f
C2361 vdd.t129 gnd 0.037975f
C2362 vdd.n5 gnd 0.29902f
C2363 vdd.n6 gnd 0.130857f
C2364 vdd.t123 gnd 0.037975f
C2365 vdd.t121 gnd 0.037975f
C2366 vdd.n7 gnd 0.299515f
C2367 vdd.t102 gnd 0.037975f
C2368 vdd.t108 gnd 0.037975f
C2369 vdd.n8 gnd 0.29902f
C2370 vdd.n9 gnd 0.275754f
C2371 vdd.t4 gnd 0.037975f
C2372 vdd.t133 gnd 0.037975f
C2373 vdd.n10 gnd 0.29902f
C2374 vdd.n11 gnd 0.139459f
C2375 vdd.t126 gnd 0.037975f
C2376 vdd.t6 gnd 0.037975f
C2377 vdd.n12 gnd 0.29902f
C2378 vdd.n13 gnd 0.130857f
C2379 vdd.n14 gnd 0.092513f
C2380 vdd.t301 gnd 0.021097f
C2381 vdd.t16 gnd 0.021097f
C2382 vdd.n15 gnd 0.194191f
C2383 vdd.t12 gnd 0.021097f
C2384 vdd.t113 gnd 0.021097f
C2385 vdd.n16 gnd 0.193623f
C2386 vdd.n17 gnd 0.336964f
C2387 vdd.t116 gnd 0.021097f
C2388 vdd.t98 gnd 0.021097f
C2389 vdd.n18 gnd 0.193623f
C2390 vdd.n19 gnd 0.139406f
C2391 vdd.t13 gnd 0.021097f
C2392 vdd.t17 gnd 0.021097f
C2393 vdd.n20 gnd 0.194191f
C2394 vdd.t115 gnd 0.021097f
C2395 vdd.t100 gnd 0.021097f
C2396 vdd.n21 gnd 0.193623f
C2397 vdd.n22 gnd 0.336964f
C2398 vdd.t18 gnd 0.021097f
C2399 vdd.t112 gnd 0.021097f
C2400 vdd.n23 gnd 0.193623f
C2401 vdd.n24 gnd 0.139406f
C2402 vdd.t135 gnd 0.021097f
C2403 vdd.t99 gnd 0.021097f
C2404 vdd.n25 gnd 0.193623f
C2405 vdd.t136 gnd 0.021097f
C2406 vdd.t134 gnd 0.021097f
C2407 vdd.n26 gnd 0.193623f
C2408 vdd.n27 gnd 22.5087f
C2409 vdd.n28 gnd 8.71067f
C2410 vdd.n29 gnd 0.005754f
C2411 vdd.n30 gnd 0.00534f
C2412 vdd.n31 gnd 0.002954f
C2413 vdd.n32 gnd 0.006782f
C2414 vdd.n33 gnd 0.002869f
C2415 vdd.n34 gnd 0.003038f
C2416 vdd.n35 gnd 0.00534f
C2417 vdd.n36 gnd 0.002869f
C2418 vdd.n37 gnd 0.006782f
C2419 vdd.n38 gnd 0.003038f
C2420 vdd.n39 gnd 0.00534f
C2421 vdd.n40 gnd 0.002869f
C2422 vdd.n41 gnd 0.005086f
C2423 vdd.n42 gnd 0.005102f
C2424 vdd.t270 gnd 0.01457f
C2425 vdd.n43 gnd 0.032418f
C2426 vdd.n44 gnd 0.168712f
C2427 vdd.n45 gnd 0.002869f
C2428 vdd.n46 gnd 0.003038f
C2429 vdd.n47 gnd 0.006782f
C2430 vdd.n48 gnd 0.006782f
C2431 vdd.n49 gnd 0.003038f
C2432 vdd.n50 gnd 0.002869f
C2433 vdd.n51 gnd 0.00534f
C2434 vdd.n52 gnd 0.00534f
C2435 vdd.n53 gnd 0.002869f
C2436 vdd.n54 gnd 0.003038f
C2437 vdd.n55 gnd 0.006782f
C2438 vdd.n56 gnd 0.006782f
C2439 vdd.n57 gnd 0.003038f
C2440 vdd.n58 gnd 0.002869f
C2441 vdd.n59 gnd 0.00534f
C2442 vdd.n60 gnd 0.00534f
C2443 vdd.n61 gnd 0.002869f
C2444 vdd.n62 gnd 0.003038f
C2445 vdd.n63 gnd 0.006782f
C2446 vdd.n64 gnd 0.006782f
C2447 vdd.n65 gnd 0.016034f
C2448 vdd.n66 gnd 0.002954f
C2449 vdd.n67 gnd 0.002869f
C2450 vdd.n68 gnd 0.013801f
C2451 vdd.n69 gnd 0.009635f
C2452 vdd.t150 gnd 0.033756f
C2453 vdd.t202 gnd 0.033756f
C2454 vdd.n70 gnd 0.231991f
C2455 vdd.n71 gnd 0.182426f
C2456 vdd.t164 gnd 0.033756f
C2457 vdd.t228 gnd 0.033756f
C2458 vdd.n72 gnd 0.231991f
C2459 vdd.n73 gnd 0.147217f
C2460 vdd.t193 gnd 0.033756f
C2461 vdd.t276 gnd 0.033756f
C2462 vdd.n74 gnd 0.231991f
C2463 vdd.n75 gnd 0.147217f
C2464 vdd.t169 gnd 0.033756f
C2465 vdd.t257 gnd 0.033756f
C2466 vdd.n76 gnd 0.231991f
C2467 vdd.n77 gnd 0.147217f
C2468 vdd.t174 gnd 0.033756f
C2469 vdd.t272 gnd 0.033756f
C2470 vdd.n78 gnd 0.231991f
C2471 vdd.n79 gnd 0.147217f
C2472 vdd.t211 gnd 0.033756f
C2473 vdd.t284 gnd 0.033756f
C2474 vdd.n80 gnd 0.231991f
C2475 vdd.n81 gnd 0.147217f
C2476 vdd.t231 gnd 0.033756f
C2477 vdd.t263 gnd 0.033756f
C2478 vdd.n82 gnd 0.231991f
C2479 vdd.n83 gnd 0.147217f
C2480 vdd.t196 gnd 0.033756f
C2481 vdd.t278 gnd 0.033756f
C2482 vdd.n84 gnd 0.231991f
C2483 vdd.n85 gnd 0.147217f
C2484 vdd.t220 gnd 0.033756f
C2485 vdd.t294 gnd 0.033756f
C2486 vdd.n86 gnd 0.231991f
C2487 vdd.n87 gnd 0.147217f
C2488 vdd.n88 gnd 0.005754f
C2489 vdd.n89 gnd 0.00534f
C2490 vdd.n90 gnd 0.002954f
C2491 vdd.n91 gnd 0.006782f
C2492 vdd.n92 gnd 0.002869f
C2493 vdd.n93 gnd 0.003038f
C2494 vdd.n94 gnd 0.00534f
C2495 vdd.n95 gnd 0.002869f
C2496 vdd.n96 gnd 0.006782f
C2497 vdd.n97 gnd 0.003038f
C2498 vdd.n98 gnd 0.00534f
C2499 vdd.n99 gnd 0.002869f
C2500 vdd.n100 gnd 0.005086f
C2501 vdd.n101 gnd 0.005102f
C2502 vdd.t244 gnd 0.01457f
C2503 vdd.n102 gnd 0.032418f
C2504 vdd.n103 gnd 0.168712f
C2505 vdd.n104 gnd 0.002869f
C2506 vdd.n105 gnd 0.003038f
C2507 vdd.n106 gnd 0.006782f
C2508 vdd.n107 gnd 0.006782f
C2509 vdd.n108 gnd 0.003038f
C2510 vdd.n109 gnd 0.002869f
C2511 vdd.n110 gnd 0.00534f
C2512 vdd.n111 gnd 0.00534f
C2513 vdd.n112 gnd 0.002869f
C2514 vdd.n113 gnd 0.003038f
C2515 vdd.n114 gnd 0.006782f
C2516 vdd.n115 gnd 0.006782f
C2517 vdd.n116 gnd 0.003038f
C2518 vdd.n117 gnd 0.002869f
C2519 vdd.n118 gnd 0.00534f
C2520 vdd.n119 gnd 0.00534f
C2521 vdd.n120 gnd 0.002869f
C2522 vdd.n121 gnd 0.003038f
C2523 vdd.n122 gnd 0.006782f
C2524 vdd.n123 gnd 0.006782f
C2525 vdd.n124 gnd 0.016034f
C2526 vdd.n125 gnd 0.002954f
C2527 vdd.n126 gnd 0.002869f
C2528 vdd.n127 gnd 0.013801f
C2529 vdd.n128 gnd 0.009333f
C2530 vdd.n129 gnd 0.10953f
C2531 vdd.n130 gnd 0.005754f
C2532 vdd.n131 gnd 0.00534f
C2533 vdd.n132 gnd 0.002954f
C2534 vdd.n133 gnd 0.006782f
C2535 vdd.n134 gnd 0.002869f
C2536 vdd.n135 gnd 0.003038f
C2537 vdd.n136 gnd 0.00534f
C2538 vdd.n137 gnd 0.002869f
C2539 vdd.n138 gnd 0.006782f
C2540 vdd.n139 gnd 0.003038f
C2541 vdd.n140 gnd 0.00534f
C2542 vdd.n141 gnd 0.002869f
C2543 vdd.n142 gnd 0.005086f
C2544 vdd.n143 gnd 0.005102f
C2545 vdd.t201 gnd 0.01457f
C2546 vdd.n144 gnd 0.032418f
C2547 vdd.n145 gnd 0.168712f
C2548 vdd.n146 gnd 0.002869f
C2549 vdd.n147 gnd 0.003038f
C2550 vdd.n148 gnd 0.006782f
C2551 vdd.n149 gnd 0.006782f
C2552 vdd.n150 gnd 0.003038f
C2553 vdd.n151 gnd 0.002869f
C2554 vdd.n152 gnd 0.00534f
C2555 vdd.n153 gnd 0.00534f
C2556 vdd.n154 gnd 0.002869f
C2557 vdd.n155 gnd 0.003038f
C2558 vdd.n156 gnd 0.006782f
C2559 vdd.n157 gnd 0.006782f
C2560 vdd.n158 gnd 0.003038f
C2561 vdd.n159 gnd 0.002869f
C2562 vdd.n160 gnd 0.00534f
C2563 vdd.n161 gnd 0.00534f
C2564 vdd.n162 gnd 0.002869f
C2565 vdd.n163 gnd 0.003038f
C2566 vdd.n164 gnd 0.006782f
C2567 vdd.n165 gnd 0.006782f
C2568 vdd.n166 gnd 0.016034f
C2569 vdd.n167 gnd 0.002954f
C2570 vdd.n168 gnd 0.002869f
C2571 vdd.n169 gnd 0.013801f
C2572 vdd.n170 gnd 0.009635f
C2573 vdd.t286 gnd 0.033756f
C2574 vdd.t188 gnd 0.033756f
C2575 vdd.n171 gnd 0.231991f
C2576 vdd.n172 gnd 0.182426f
C2577 vdd.t191 gnd 0.033756f
C2578 vdd.t282 gnd 0.033756f
C2579 vdd.n173 gnd 0.231991f
C2580 vdd.n174 gnd 0.147217f
C2581 vdd.t283 gnd 0.033756f
C2582 vdd.t162 gnd 0.033756f
C2583 vdd.n175 gnd 0.231991f
C2584 vdd.n176 gnd 0.147217f
C2585 vdd.t265 gnd 0.033756f
C2586 vdd.t275 gnd 0.033756f
C2587 vdd.n177 gnd 0.231991f
C2588 vdd.n178 gnd 0.147217f
C2589 vdd.t156 gnd 0.033756f
C2590 vdd.t226 gnd 0.033756f
C2591 vdd.n179 gnd 0.231991f
C2592 vdd.n180 gnd 0.147217f
C2593 vdd.t262 gnd 0.033756f
C2594 vdd.t290 gnd 0.033756f
C2595 vdd.n181 gnd 0.231991f
C2596 vdd.n182 gnd 0.147217f
C2597 vdd.t199 gnd 0.033756f
C2598 vdd.t261 gnd 0.033756f
C2599 vdd.n183 gnd 0.231991f
C2600 vdd.n184 gnd 0.147217f
C2601 vdd.t298 gnd 0.033756f
C2602 vdd.t190 gnd 0.033756f
C2603 vdd.n185 gnd 0.231991f
C2604 vdd.n186 gnd 0.147217f
C2605 vdd.t242 gnd 0.033756f
C2606 vdd.t281 gnd 0.033756f
C2607 vdd.n187 gnd 0.231991f
C2608 vdd.n188 gnd 0.147217f
C2609 vdd.n189 gnd 0.005754f
C2610 vdd.n190 gnd 0.00534f
C2611 vdd.n191 gnd 0.002954f
C2612 vdd.n192 gnd 0.006782f
C2613 vdd.n193 gnd 0.002869f
C2614 vdd.n194 gnd 0.003038f
C2615 vdd.n195 gnd 0.00534f
C2616 vdd.n196 gnd 0.002869f
C2617 vdd.n197 gnd 0.006782f
C2618 vdd.n198 gnd 0.003038f
C2619 vdd.n199 gnd 0.00534f
C2620 vdd.n200 gnd 0.002869f
C2621 vdd.n201 gnd 0.005086f
C2622 vdd.n202 gnd 0.005102f
C2623 vdd.t160 gnd 0.01457f
C2624 vdd.n203 gnd 0.032418f
C2625 vdd.n204 gnd 0.168712f
C2626 vdd.n205 gnd 0.002869f
C2627 vdd.n206 gnd 0.003038f
C2628 vdd.n207 gnd 0.006782f
C2629 vdd.n208 gnd 0.006782f
C2630 vdd.n209 gnd 0.003038f
C2631 vdd.n210 gnd 0.002869f
C2632 vdd.n211 gnd 0.00534f
C2633 vdd.n212 gnd 0.00534f
C2634 vdd.n213 gnd 0.002869f
C2635 vdd.n214 gnd 0.003038f
C2636 vdd.n215 gnd 0.006782f
C2637 vdd.n216 gnd 0.006782f
C2638 vdd.n217 gnd 0.003038f
C2639 vdd.n218 gnd 0.002869f
C2640 vdd.n219 gnd 0.00534f
C2641 vdd.n220 gnd 0.00534f
C2642 vdd.n221 gnd 0.002869f
C2643 vdd.n222 gnd 0.003038f
C2644 vdd.n223 gnd 0.006782f
C2645 vdd.n224 gnd 0.006782f
C2646 vdd.n225 gnd 0.016034f
C2647 vdd.n226 gnd 0.002954f
C2648 vdd.n227 gnd 0.002869f
C2649 vdd.n228 gnd 0.013801f
C2650 vdd.n229 gnd 0.009333f
C2651 vdd.n230 gnd 0.065159f
C2652 vdd.n231 gnd 0.234786f
C2653 vdd.n232 gnd 0.005754f
C2654 vdd.n233 gnd 0.00534f
C2655 vdd.n234 gnd 0.002954f
C2656 vdd.n235 gnd 0.006782f
C2657 vdd.n236 gnd 0.002869f
C2658 vdd.n237 gnd 0.003038f
C2659 vdd.n238 gnd 0.00534f
C2660 vdd.n239 gnd 0.002869f
C2661 vdd.n240 gnd 0.006782f
C2662 vdd.n241 gnd 0.003038f
C2663 vdd.n242 gnd 0.00534f
C2664 vdd.n243 gnd 0.002869f
C2665 vdd.n244 gnd 0.005086f
C2666 vdd.n245 gnd 0.005102f
C2667 vdd.t221 gnd 0.01457f
C2668 vdd.n246 gnd 0.032418f
C2669 vdd.n247 gnd 0.168712f
C2670 vdd.n248 gnd 0.002869f
C2671 vdd.n249 gnd 0.003038f
C2672 vdd.n250 gnd 0.006782f
C2673 vdd.n251 gnd 0.006782f
C2674 vdd.n252 gnd 0.003038f
C2675 vdd.n253 gnd 0.002869f
C2676 vdd.n254 gnd 0.00534f
C2677 vdd.n255 gnd 0.00534f
C2678 vdd.n256 gnd 0.002869f
C2679 vdd.n257 gnd 0.003038f
C2680 vdd.n258 gnd 0.006782f
C2681 vdd.n259 gnd 0.006782f
C2682 vdd.n260 gnd 0.003038f
C2683 vdd.n261 gnd 0.002869f
C2684 vdd.n262 gnd 0.00534f
C2685 vdd.n263 gnd 0.00534f
C2686 vdd.n264 gnd 0.002869f
C2687 vdd.n265 gnd 0.003038f
C2688 vdd.n266 gnd 0.006782f
C2689 vdd.n267 gnd 0.006782f
C2690 vdd.n268 gnd 0.016034f
C2691 vdd.n269 gnd 0.002954f
C2692 vdd.n270 gnd 0.002869f
C2693 vdd.n271 gnd 0.013801f
C2694 vdd.n272 gnd 0.009635f
C2695 vdd.t297 gnd 0.033756f
C2696 vdd.t214 gnd 0.033756f
C2697 vdd.n273 gnd 0.231991f
C2698 vdd.n274 gnd 0.182426f
C2699 vdd.t216 gnd 0.033756f
C2700 vdd.t291 gnd 0.033756f
C2701 vdd.n275 gnd 0.231991f
C2702 vdd.n276 gnd 0.147217f
C2703 vdd.t293 gnd 0.033756f
C2704 vdd.t185 gnd 0.033756f
C2705 vdd.n277 gnd 0.231991f
C2706 vdd.n278 gnd 0.147217f
C2707 vdd.t274 gnd 0.033756f
C2708 vdd.t289 gnd 0.033756f
C2709 vdd.n279 gnd 0.231991f
C2710 vdd.n280 gnd 0.147217f
C2711 vdd.t175 gnd 0.033756f
C2712 vdd.t245 gnd 0.033756f
C2713 vdd.n281 gnd 0.231991f
C2714 vdd.n282 gnd 0.147217f
C2715 vdd.t273 gnd 0.033756f
C2716 vdd.t146 gnd 0.033756f
C2717 vdd.n283 gnd 0.231991f
C2718 vdd.n284 gnd 0.147217f
C2719 vdd.t218 gnd 0.033756f
C2720 vdd.t271 gnd 0.033756f
C2721 vdd.n285 gnd 0.231991f
C2722 vdd.n286 gnd 0.147217f
C2723 vdd.t158 gnd 0.033756f
C2724 vdd.t215 gnd 0.033756f
C2725 vdd.n287 gnd 0.231991f
C2726 vdd.n288 gnd 0.147217f
C2727 vdd.t251 gnd 0.033756f
C2728 vdd.t292 gnd 0.033756f
C2729 vdd.n289 gnd 0.231991f
C2730 vdd.n290 gnd 0.147217f
C2731 vdd.n291 gnd 0.005754f
C2732 vdd.n292 gnd 0.00534f
C2733 vdd.n293 gnd 0.002954f
C2734 vdd.n294 gnd 0.006782f
C2735 vdd.n295 gnd 0.002869f
C2736 vdd.n296 gnd 0.003038f
C2737 vdd.n297 gnd 0.00534f
C2738 vdd.n298 gnd 0.002869f
C2739 vdd.n299 gnd 0.006782f
C2740 vdd.n300 gnd 0.003038f
C2741 vdd.n301 gnd 0.00534f
C2742 vdd.n302 gnd 0.002869f
C2743 vdd.n303 gnd 0.005086f
C2744 vdd.n304 gnd 0.005102f
C2745 vdd.t180 gnd 0.01457f
C2746 vdd.n305 gnd 0.032418f
C2747 vdd.n306 gnd 0.168712f
C2748 vdd.n307 gnd 0.002869f
C2749 vdd.n308 gnd 0.003038f
C2750 vdd.n309 gnd 0.006782f
C2751 vdd.n310 gnd 0.006782f
C2752 vdd.n311 gnd 0.003038f
C2753 vdd.n312 gnd 0.002869f
C2754 vdd.n313 gnd 0.00534f
C2755 vdd.n314 gnd 0.00534f
C2756 vdd.n315 gnd 0.002869f
C2757 vdd.n316 gnd 0.003038f
C2758 vdd.n317 gnd 0.006782f
C2759 vdd.n318 gnd 0.006782f
C2760 vdd.n319 gnd 0.003038f
C2761 vdd.n320 gnd 0.002869f
C2762 vdd.n321 gnd 0.00534f
C2763 vdd.n322 gnd 0.00534f
C2764 vdd.n323 gnd 0.002869f
C2765 vdd.n324 gnd 0.003038f
C2766 vdd.n325 gnd 0.006782f
C2767 vdd.n326 gnd 0.006782f
C2768 vdd.n327 gnd 0.016034f
C2769 vdd.n328 gnd 0.002954f
C2770 vdd.n329 gnd 0.002869f
C2771 vdd.n330 gnd 0.013801f
C2772 vdd.n331 gnd 0.009333f
C2773 vdd.n332 gnd 0.065159f
C2774 vdd.n333 gnd 0.268779f
C2775 vdd.n334 gnd 0.008058f
C2776 vdd.n335 gnd 0.010485f
C2777 vdd.n336 gnd 0.008439f
C2778 vdd.n337 gnd 0.008439f
C2779 vdd.n338 gnd 0.010485f
C2780 vdd.n339 gnd 0.010485f
C2781 vdd.n340 gnd 0.76611f
C2782 vdd.n341 gnd 0.010485f
C2783 vdd.n342 gnd 0.010485f
C2784 vdd.n343 gnd 0.010485f
C2785 vdd.n344 gnd 0.830399f
C2786 vdd.n345 gnd 0.010485f
C2787 vdd.n346 gnd 0.010485f
C2788 vdd.n347 gnd 0.010485f
C2789 vdd.n348 gnd 0.010485f
C2790 vdd.n349 gnd 0.008439f
C2791 vdd.n350 gnd 0.010485f
C2792 vdd.t145 gnd 0.535742f
C2793 vdd.n351 gnd 0.010485f
C2794 vdd.n352 gnd 0.010485f
C2795 vdd.n353 gnd 0.010485f
C2796 vdd.t260 gnd 0.535742f
C2797 vdd.n354 gnd 0.010485f
C2798 vdd.n355 gnd 0.010485f
C2799 vdd.n356 gnd 0.010485f
C2800 vdd.n357 gnd 0.010485f
C2801 vdd.n358 gnd 0.010485f
C2802 vdd.n359 gnd 0.008439f
C2803 vdd.n360 gnd 0.010485f
C2804 vdd.n361 gnd 0.605388f
C2805 vdd.n362 gnd 0.010485f
C2806 vdd.n363 gnd 0.010485f
C2807 vdd.n364 gnd 0.010485f
C2808 vdd.t189 gnd 0.535742f
C2809 vdd.n365 gnd 0.010485f
C2810 vdd.n366 gnd 0.010485f
C2811 vdd.n367 gnd 0.010485f
C2812 vdd.n368 gnd 0.010485f
C2813 vdd.n369 gnd 0.010485f
C2814 vdd.n370 gnd 0.008439f
C2815 vdd.n371 gnd 0.010485f
C2816 vdd.t219 gnd 0.535742f
C2817 vdd.n372 gnd 0.010485f
C2818 vdd.n373 gnd 0.010485f
C2819 vdd.n374 gnd 0.010485f
C2820 vdd.n375 gnd 0.626818f
C2821 vdd.n376 gnd 0.010485f
C2822 vdd.n377 gnd 0.010485f
C2823 vdd.n378 gnd 0.010485f
C2824 vdd.n379 gnd 0.010485f
C2825 vdd.n380 gnd 0.010485f
C2826 vdd.n381 gnd 0.008439f
C2827 vdd.n382 gnd 0.010485f
C2828 vdd.t159 gnd 0.535742f
C2829 vdd.n383 gnd 0.010485f
C2830 vdd.n384 gnd 0.010485f
C2831 vdd.n385 gnd 0.010485f
C2832 vdd.n386 gnd 0.541099f
C2833 vdd.n387 gnd 0.010485f
C2834 vdd.n388 gnd 0.010485f
C2835 vdd.n389 gnd 0.010485f
C2836 vdd.n390 gnd 0.010485f
C2837 vdd.n391 gnd 0.025363f
C2838 vdd.n392 gnd 0.025907f
C2839 vdd.t34 gnd 0.535742f
C2840 vdd.n393 gnd 0.025363f
C2841 vdd.n425 gnd 0.010485f
C2842 vdd.t62 gnd 0.128989f
C2843 vdd.t61 gnd 0.137854f
C2844 vdd.t60 gnd 0.168458f
C2845 vdd.n426 gnd 0.215939f
C2846 vdd.n427 gnd 0.182272f
C2847 vdd.n428 gnd 0.01384f
C2848 vdd.n429 gnd 0.010485f
C2849 vdd.n430 gnd 0.008439f
C2850 vdd.n431 gnd 0.010485f
C2851 vdd.n432 gnd 0.008439f
C2852 vdd.n433 gnd 0.010485f
C2853 vdd.n434 gnd 0.008439f
C2854 vdd.n435 gnd 0.010485f
C2855 vdd.n436 gnd 0.008439f
C2856 vdd.n437 gnd 0.010485f
C2857 vdd.n438 gnd 0.008439f
C2858 vdd.n439 gnd 0.010485f
C2859 vdd.t36 gnd 0.128989f
C2860 vdd.t35 gnd 0.137854f
C2861 vdd.t33 gnd 0.168458f
C2862 vdd.n440 gnd 0.215939f
C2863 vdd.n441 gnd 0.182272f
C2864 vdd.n442 gnd 0.008439f
C2865 vdd.n443 gnd 0.010485f
C2866 vdd.n444 gnd 0.008439f
C2867 vdd.n445 gnd 0.010485f
C2868 vdd.n446 gnd 0.008439f
C2869 vdd.n447 gnd 0.010485f
C2870 vdd.n448 gnd 0.008439f
C2871 vdd.n449 gnd 0.010485f
C2872 vdd.n450 gnd 0.008439f
C2873 vdd.n451 gnd 0.010485f
C2874 vdd.t53 gnd 0.128989f
C2875 vdd.t52 gnd 0.137854f
C2876 vdd.t51 gnd 0.168458f
C2877 vdd.n452 gnd 0.215939f
C2878 vdd.n453 gnd 0.182272f
C2879 vdd.n454 gnd 0.018059f
C2880 vdd.n455 gnd 0.010485f
C2881 vdd.n456 gnd 0.008439f
C2882 vdd.n457 gnd 0.010485f
C2883 vdd.n458 gnd 0.008439f
C2884 vdd.n459 gnd 0.010485f
C2885 vdd.n460 gnd 0.008439f
C2886 vdd.n461 gnd 0.010485f
C2887 vdd.n462 gnd 0.008439f
C2888 vdd.n463 gnd 0.010485f
C2889 vdd.n464 gnd 0.025907f
C2890 vdd.n465 gnd 0.007004f
C2891 vdd.n466 gnd 0.008439f
C2892 vdd.n467 gnd 0.010485f
C2893 vdd.n468 gnd 0.010485f
C2894 vdd.n469 gnd 0.008439f
C2895 vdd.n470 gnd 0.010485f
C2896 vdd.n471 gnd 0.010485f
C2897 vdd.n472 gnd 0.010485f
C2898 vdd.n473 gnd 0.010485f
C2899 vdd.n474 gnd 0.010485f
C2900 vdd.n475 gnd 0.008439f
C2901 vdd.n476 gnd 0.008439f
C2902 vdd.n477 gnd 0.010485f
C2903 vdd.n478 gnd 0.010485f
C2904 vdd.n479 gnd 0.008439f
C2905 vdd.n480 gnd 0.010485f
C2906 vdd.n481 gnd 0.010485f
C2907 vdd.n482 gnd 0.010485f
C2908 vdd.n483 gnd 0.010485f
C2909 vdd.n484 gnd 0.010485f
C2910 vdd.n485 gnd 0.008439f
C2911 vdd.n486 gnd 0.008439f
C2912 vdd.n487 gnd 0.010485f
C2913 vdd.n488 gnd 0.010485f
C2914 vdd.n489 gnd 0.008439f
C2915 vdd.n490 gnd 0.010485f
C2916 vdd.n491 gnd 0.010485f
C2917 vdd.n492 gnd 0.010485f
C2918 vdd.n493 gnd 0.010485f
C2919 vdd.n494 gnd 0.010485f
C2920 vdd.n495 gnd 0.008439f
C2921 vdd.n496 gnd 0.008439f
C2922 vdd.n497 gnd 0.010485f
C2923 vdd.n498 gnd 0.010485f
C2924 vdd.n499 gnd 0.008439f
C2925 vdd.n500 gnd 0.010485f
C2926 vdd.n501 gnd 0.010485f
C2927 vdd.n502 gnd 0.010485f
C2928 vdd.n503 gnd 0.010485f
C2929 vdd.n504 gnd 0.010485f
C2930 vdd.n505 gnd 0.008439f
C2931 vdd.n506 gnd 0.008439f
C2932 vdd.n507 gnd 0.010485f
C2933 vdd.n508 gnd 0.010485f
C2934 vdd.n509 gnd 0.007046f
C2935 vdd.n510 gnd 0.010485f
C2936 vdd.n511 gnd 0.010485f
C2937 vdd.n512 gnd 0.010485f
C2938 vdd.n513 gnd 0.010485f
C2939 vdd.n514 gnd 0.010485f
C2940 vdd.n515 gnd 0.007046f
C2941 vdd.n516 gnd 0.008439f
C2942 vdd.n517 gnd 0.010485f
C2943 vdd.n518 gnd 0.010485f
C2944 vdd.n519 gnd 0.008439f
C2945 vdd.n520 gnd 0.010485f
C2946 vdd.n521 gnd 0.010485f
C2947 vdd.n522 gnd 0.010485f
C2948 vdd.n523 gnd 0.010485f
C2949 vdd.n524 gnd 0.010485f
C2950 vdd.n525 gnd 0.008439f
C2951 vdd.n526 gnd 0.008439f
C2952 vdd.n527 gnd 0.010485f
C2953 vdd.n528 gnd 0.010485f
C2954 vdd.n529 gnd 0.008439f
C2955 vdd.n530 gnd 0.010485f
C2956 vdd.n531 gnd 0.010485f
C2957 vdd.n532 gnd 0.010485f
C2958 vdd.n533 gnd 0.010485f
C2959 vdd.n534 gnd 0.010485f
C2960 vdd.n535 gnd 0.008439f
C2961 vdd.n536 gnd 0.008439f
C2962 vdd.n537 gnd 0.010485f
C2963 vdd.n538 gnd 0.010485f
C2964 vdd.n539 gnd 0.008439f
C2965 vdd.n540 gnd 0.010485f
C2966 vdd.n541 gnd 0.010485f
C2967 vdd.n542 gnd 0.010485f
C2968 vdd.n543 gnd 0.010485f
C2969 vdd.n544 gnd 0.010485f
C2970 vdd.n545 gnd 0.008439f
C2971 vdd.n546 gnd 0.008439f
C2972 vdd.n547 gnd 0.010485f
C2973 vdd.n548 gnd 0.010485f
C2974 vdd.n549 gnd 0.008439f
C2975 vdd.n550 gnd 0.010485f
C2976 vdd.n551 gnd 0.010485f
C2977 vdd.n552 gnd 0.010485f
C2978 vdd.n553 gnd 0.010485f
C2979 vdd.n554 gnd 0.010485f
C2980 vdd.n555 gnd 0.008439f
C2981 vdd.n556 gnd 0.008439f
C2982 vdd.n557 gnd 0.010485f
C2983 vdd.n558 gnd 0.010485f
C2984 vdd.n559 gnd 0.008439f
C2985 vdd.n560 gnd 0.010485f
C2986 vdd.n561 gnd 0.010485f
C2987 vdd.n562 gnd 0.010485f
C2988 vdd.n563 gnd 0.010485f
C2989 vdd.n564 gnd 0.010485f
C2990 vdd.n565 gnd 0.005738f
C2991 vdd.n566 gnd 0.018059f
C2992 vdd.n567 gnd 0.010485f
C2993 vdd.n568 gnd 0.010485f
C2994 vdd.n569 gnd 0.008354f
C2995 vdd.n570 gnd 0.010485f
C2996 vdd.n571 gnd 0.010485f
C2997 vdd.n572 gnd 0.010485f
C2998 vdd.n573 gnd 0.010485f
C2999 vdd.n574 gnd 0.010485f
C3000 vdd.n575 gnd 0.008439f
C3001 vdd.n576 gnd 0.008439f
C3002 vdd.n577 gnd 0.010485f
C3003 vdd.n578 gnd 0.010485f
C3004 vdd.n579 gnd 0.008439f
C3005 vdd.n580 gnd 0.010485f
C3006 vdd.n581 gnd 0.010485f
C3007 vdd.n582 gnd 0.010485f
C3008 vdd.n583 gnd 0.010485f
C3009 vdd.n584 gnd 0.010485f
C3010 vdd.n585 gnd 0.008439f
C3011 vdd.n586 gnd 0.008439f
C3012 vdd.n587 gnd 0.010485f
C3013 vdd.n588 gnd 0.010485f
C3014 vdd.n589 gnd 0.008439f
C3015 vdd.n590 gnd 0.010485f
C3016 vdd.n591 gnd 0.010485f
C3017 vdd.n592 gnd 0.010485f
C3018 vdd.n593 gnd 0.010485f
C3019 vdd.n594 gnd 0.010485f
C3020 vdd.n595 gnd 0.008439f
C3021 vdd.n596 gnd 0.008439f
C3022 vdd.n597 gnd 0.010485f
C3023 vdd.n598 gnd 0.010485f
C3024 vdd.n599 gnd 0.008439f
C3025 vdd.n600 gnd 0.010485f
C3026 vdd.n601 gnd 0.010485f
C3027 vdd.n602 gnd 0.010485f
C3028 vdd.n603 gnd 0.010485f
C3029 vdd.n604 gnd 0.010485f
C3030 vdd.n605 gnd 0.008439f
C3031 vdd.n606 gnd 0.008439f
C3032 vdd.n607 gnd 0.010485f
C3033 vdd.n608 gnd 0.010485f
C3034 vdd.n609 gnd 0.008439f
C3035 vdd.n610 gnd 0.010485f
C3036 vdd.n611 gnd 0.010485f
C3037 vdd.n612 gnd 0.010485f
C3038 vdd.n613 gnd 0.010485f
C3039 vdd.n614 gnd 0.010485f
C3040 vdd.n615 gnd 0.008439f
C3041 vdd.n616 gnd 0.010485f
C3042 vdd.n617 gnd 0.008439f
C3043 vdd.n618 gnd 0.00443f
C3044 vdd.n619 gnd 0.010485f
C3045 vdd.n620 gnd 0.010485f
C3046 vdd.n621 gnd 0.008439f
C3047 vdd.n622 gnd 0.010485f
C3048 vdd.n623 gnd 0.008439f
C3049 vdd.n624 gnd 0.010485f
C3050 vdd.n625 gnd 0.008439f
C3051 vdd.n626 gnd 0.010485f
C3052 vdd.n627 gnd 0.008439f
C3053 vdd.n628 gnd 0.010485f
C3054 vdd.n629 gnd 0.008439f
C3055 vdd.n630 gnd 0.010485f
C3056 vdd.n631 gnd 0.008439f
C3057 vdd.n632 gnd 0.010485f
C3058 vdd.n633 gnd 0.583958f
C3059 vdd.t155 gnd 0.535742f
C3060 vdd.n634 gnd 0.010485f
C3061 vdd.n635 gnd 0.008439f
C3062 vdd.n636 gnd 0.010485f
C3063 vdd.n637 gnd 0.008439f
C3064 vdd.n638 gnd 0.010485f
C3065 vdd.t168 gnd 0.535742f
C3066 vdd.n639 gnd 0.010485f
C3067 vdd.n640 gnd 0.008439f
C3068 vdd.n641 gnd 0.010485f
C3069 vdd.n642 gnd 0.008439f
C3070 vdd.n643 gnd 0.010485f
C3071 vdd.t161 gnd 0.535742f
C3072 vdd.n644 gnd 0.669677f
C3073 vdd.n645 gnd 0.010485f
C3074 vdd.n646 gnd 0.008439f
C3075 vdd.n647 gnd 0.010485f
C3076 vdd.n648 gnd 0.008439f
C3077 vdd.n649 gnd 0.010485f
C3078 vdd.t192 gnd 0.535742f
C3079 vdd.n650 gnd 0.010485f
C3080 vdd.n651 gnd 0.008439f
C3081 vdd.n652 gnd 0.010485f
C3082 vdd.n653 gnd 0.008439f
C3083 vdd.n654 gnd 0.010485f
C3084 vdd.n655 gnd 0.744681f
C3085 vdd.n656 gnd 0.889331f
C3086 vdd.t227 gnd 0.535742f
C3087 vdd.n657 gnd 0.010485f
C3088 vdd.n658 gnd 0.008439f
C3089 vdd.n659 gnd 0.010485f
C3090 vdd.n660 gnd 0.008439f
C3091 vdd.n661 gnd 0.010485f
C3092 vdd.n662 gnd 0.562529f
C3093 vdd.n663 gnd 0.010485f
C3094 vdd.n664 gnd 0.008439f
C3095 vdd.n665 gnd 0.010485f
C3096 vdd.n666 gnd 0.008439f
C3097 vdd.n667 gnd 0.010485f
C3098 vdd.t149 gnd 0.535742f
C3099 vdd.t187 gnd 0.535742f
C3100 vdd.n668 gnd 0.010485f
C3101 vdd.n669 gnd 0.008439f
C3102 vdd.n670 gnd 0.010485f
C3103 vdd.n671 gnd 0.008439f
C3104 vdd.n672 gnd 0.010485f
C3105 vdd.t200 gnd 0.535742f
C3106 vdd.n673 gnd 0.010485f
C3107 vdd.n674 gnd 0.008439f
C3108 vdd.n675 gnd 0.010485f
C3109 vdd.n676 gnd 0.008439f
C3110 vdd.n677 gnd 0.010485f
C3111 vdd.n678 gnd 1.07148f
C3112 vdd.n679 gnd 0.873259f
C3113 vdd.n680 gnd 0.010485f
C3114 vdd.n681 gnd 0.008439f
C3115 vdd.n682 gnd 0.025363f
C3116 vdd.n683 gnd 0.007004f
C3117 vdd.n684 gnd 0.025363f
C3118 vdd.t22 gnd 0.535742f
C3119 vdd.n685 gnd 0.025363f
C3120 vdd.n686 gnd 0.007004f
C3121 vdd.n687 gnd 0.009017f
C3122 vdd.t45 gnd 0.128989f
C3123 vdd.t46 gnd 0.137854f
C3124 vdd.t44 gnd 0.168458f
C3125 vdd.n688 gnd 0.215939f
C3126 vdd.n689 gnd 0.181428f
C3127 vdd.n690 gnd 0.012996f
C3128 vdd.n691 gnd 0.010485f
C3129 vdd.n692 gnd 10.897f
C3130 vdd.n723 gnd 1.47329f
C3131 vdd.n724 gnd 0.010485f
C3132 vdd.n725 gnd 0.010485f
C3133 vdd.n726 gnd 0.025907f
C3134 vdd.n727 gnd 0.009017f
C3135 vdd.n728 gnd 0.010485f
C3136 vdd.n729 gnd 0.008439f
C3137 vdd.n730 gnd 0.00671f
C3138 vdd.n731 gnd 0.033466f
C3139 vdd.n732 gnd 0.008439f
C3140 vdd.n733 gnd 0.010485f
C3141 vdd.n734 gnd 0.010485f
C3142 vdd.n735 gnd 0.010485f
C3143 vdd.n736 gnd 0.010485f
C3144 vdd.n737 gnd 0.010485f
C3145 vdd.n738 gnd 0.010485f
C3146 vdd.n739 gnd 0.010485f
C3147 vdd.n740 gnd 0.010485f
C3148 vdd.n741 gnd 0.010485f
C3149 vdd.n742 gnd 0.010485f
C3150 vdd.n743 gnd 0.010485f
C3151 vdd.n744 gnd 0.010485f
C3152 vdd.n745 gnd 0.010485f
C3153 vdd.n746 gnd 0.010485f
C3154 vdd.n747 gnd 0.007046f
C3155 vdd.n748 gnd 0.010485f
C3156 vdd.n749 gnd 0.010485f
C3157 vdd.n750 gnd 0.010485f
C3158 vdd.n751 gnd 0.010485f
C3159 vdd.n752 gnd 0.010485f
C3160 vdd.n753 gnd 0.010485f
C3161 vdd.n754 gnd 0.010485f
C3162 vdd.n755 gnd 0.010485f
C3163 vdd.n756 gnd 0.010485f
C3164 vdd.n757 gnd 0.010485f
C3165 vdd.n758 gnd 0.010485f
C3166 vdd.n759 gnd 0.010485f
C3167 vdd.n760 gnd 0.010485f
C3168 vdd.n761 gnd 0.010485f
C3169 vdd.n762 gnd 0.010485f
C3170 vdd.n763 gnd 0.010485f
C3171 vdd.n764 gnd 0.010485f
C3172 vdd.n765 gnd 0.010485f
C3173 vdd.n766 gnd 0.010485f
C3174 vdd.n767 gnd 0.008354f
C3175 vdd.t23 gnd 0.128989f
C3176 vdd.t24 gnd 0.137854f
C3177 vdd.t21 gnd 0.168458f
C3178 vdd.n768 gnd 0.215939f
C3179 vdd.n769 gnd 0.181428f
C3180 vdd.n770 gnd 0.010485f
C3181 vdd.n771 gnd 0.010485f
C3182 vdd.n772 gnd 0.010485f
C3183 vdd.n773 gnd 0.010485f
C3184 vdd.n774 gnd 0.010485f
C3185 vdd.n775 gnd 0.010485f
C3186 vdd.n776 gnd 0.010485f
C3187 vdd.n777 gnd 0.010485f
C3188 vdd.n778 gnd 0.010485f
C3189 vdd.n779 gnd 0.010485f
C3190 vdd.n780 gnd 0.010485f
C3191 vdd.n781 gnd 0.010485f
C3192 vdd.n782 gnd 0.010485f
C3193 vdd.n783 gnd 0.00671f
C3194 vdd.n785 gnd 0.00713f
C3195 vdd.n786 gnd 0.00713f
C3196 vdd.n787 gnd 0.00713f
C3197 vdd.n788 gnd 0.00713f
C3198 vdd.n789 gnd 0.00713f
C3199 vdd.n790 gnd 0.00713f
C3200 vdd.n792 gnd 0.00713f
C3201 vdd.n793 gnd 0.00713f
C3202 vdd.n795 gnd 0.00713f
C3203 vdd.n796 gnd 0.00519f
C3204 vdd.n798 gnd 0.00713f
C3205 vdd.t28 gnd 0.288105f
C3206 vdd.t27 gnd 0.294911f
C3207 vdd.t25 gnd 0.188086f
C3208 vdd.n799 gnd 0.10165f
C3209 vdd.n800 gnd 0.057659f
C3210 vdd.n801 gnd 0.010189f
C3211 vdd.n802 gnd 0.016345f
C3212 vdd.n804 gnd 0.00713f
C3213 vdd.n805 gnd 0.728608f
C3214 vdd.n806 gnd 0.015441f
C3215 vdd.n807 gnd 0.015441f
C3216 vdd.n808 gnd 0.00713f
C3217 vdd.n809 gnd 0.016433f
C3218 vdd.n810 gnd 0.00713f
C3219 vdd.n811 gnd 0.00713f
C3220 vdd.n812 gnd 0.00713f
C3221 vdd.n813 gnd 0.00713f
C3222 vdd.n814 gnd 0.00713f
C3223 vdd.n816 gnd 0.00713f
C3224 vdd.n817 gnd 0.00713f
C3225 vdd.n819 gnd 0.00713f
C3226 vdd.n820 gnd 0.00713f
C3227 vdd.n822 gnd 0.00713f
C3228 vdd.n823 gnd 0.00713f
C3229 vdd.n825 gnd 0.00713f
C3230 vdd.n826 gnd 0.00713f
C3231 vdd.n828 gnd 0.00713f
C3232 vdd.n829 gnd 0.00713f
C3233 vdd.n831 gnd 0.00713f
C3234 vdd.t56 gnd 0.288105f
C3235 vdd.t55 gnd 0.294911f
C3236 vdd.t54 gnd 0.188086f
C3237 vdd.n832 gnd 0.10165f
C3238 vdd.n833 gnd 0.057659f
C3239 vdd.n834 gnd 0.00713f
C3240 vdd.n836 gnd 0.00713f
C3241 vdd.n837 gnd 0.00713f
C3242 vdd.t26 gnd 0.364304f
C3243 vdd.n838 gnd 0.00713f
C3244 vdd.n839 gnd 0.00713f
C3245 vdd.n840 gnd 0.00713f
C3246 vdd.n841 gnd 0.00713f
C3247 vdd.n842 gnd 0.00713f
C3248 vdd.n843 gnd 0.728608f
C3249 vdd.n844 gnd 0.00713f
C3250 vdd.n845 gnd 0.00713f
C3251 vdd.n846 gnd 0.594673f
C3252 vdd.n847 gnd 0.00713f
C3253 vdd.n848 gnd 0.00713f
C3254 vdd.n849 gnd 0.00713f
C3255 vdd.n850 gnd 0.00713f
C3256 vdd.n851 gnd 0.728608f
C3257 vdd.n852 gnd 0.00713f
C3258 vdd.n853 gnd 0.00713f
C3259 vdd.n854 gnd 0.00713f
C3260 vdd.n855 gnd 0.00713f
C3261 vdd.n856 gnd 0.00713f
C3262 vdd.t9 gnd 0.364304f
C3263 vdd.n857 gnd 0.00713f
C3264 vdd.n858 gnd 0.00713f
C3265 vdd.n859 gnd 0.00713f
C3266 vdd.n860 gnd 0.00713f
C3267 vdd.n861 gnd 0.00713f
C3268 vdd.t111 gnd 0.364304f
C3269 vdd.n862 gnd 0.00713f
C3270 vdd.n863 gnd 0.00713f
C3271 vdd.n864 gnd 0.723251f
C3272 vdd.n865 gnd 0.00713f
C3273 vdd.n866 gnd 0.00713f
C3274 vdd.n867 gnd 0.00713f
C3275 vdd.t7 gnd 0.364304f
C3276 vdd.n868 gnd 0.00713f
C3277 vdd.n869 gnd 0.00713f
C3278 vdd.n870 gnd 0.562529f
C3279 vdd.n871 gnd 0.00713f
C3280 vdd.n872 gnd 0.00713f
C3281 vdd.n873 gnd 0.00713f
C3282 vdd.n874 gnd 0.487525f
C3283 vdd.n875 gnd 0.00713f
C3284 vdd.n876 gnd 0.00713f
C3285 vdd.n877 gnd 0.401806f
C3286 vdd.n878 gnd 0.00713f
C3287 vdd.n879 gnd 0.00713f
C3288 vdd.n880 gnd 0.00713f
C3289 vdd.n881 gnd 0.600031f
C3290 vdd.n882 gnd 0.00713f
C3291 vdd.n883 gnd 0.00713f
C3292 vdd.t114 gnd 0.364304f
C3293 vdd.n884 gnd 0.00713f
C3294 vdd.t42 gnd 0.294911f
C3295 vdd.t40 gnd 0.188086f
C3296 vdd.t43 gnd 0.294911f
C3297 vdd.n885 gnd 0.165752f
C3298 vdd.n886 gnd 0.00713f
C3299 vdd.n887 gnd 0.00713f
C3300 vdd.n888 gnd 0.728608f
C3301 vdd.n889 gnd 0.00713f
C3302 vdd.n890 gnd 0.00713f
C3303 vdd.t41 gnd 0.283943f
C3304 vdd.t97 gnd 0.128578f
C3305 vdd.n891 gnd 0.00713f
C3306 vdd.n892 gnd 0.00713f
C3307 vdd.n893 gnd 0.00713f
C3308 vdd.t14 gnd 0.364304f
C3309 vdd.n894 gnd 0.00713f
C3310 vdd.n895 gnd 0.00713f
C3311 vdd.n896 gnd 0.00713f
C3312 vdd.n897 gnd 0.00713f
C3313 vdd.n898 gnd 0.00713f
C3314 vdd.t15 gnd 0.364304f
C3315 vdd.n899 gnd 0.00713f
C3316 vdd.n900 gnd 0.00713f
C3317 vdd.n901 gnd 0.648247f
C3318 vdd.n902 gnd 0.00713f
C3319 vdd.n903 gnd 0.00713f
C3320 vdd.n904 gnd 0.00713f
C3321 vdd.n905 gnd 0.401806f
C3322 vdd.n906 gnd 0.00713f
C3323 vdd.n907 gnd 0.00713f
C3324 vdd.t120 gnd 0.364304f
C3325 vdd.n908 gnd 0.00713f
C3326 vdd.n909 gnd 0.00713f
C3327 vdd.n910 gnd 0.00713f
C3328 vdd.n911 gnd 0.562529f
C3329 vdd.n912 gnd 0.00713f
C3330 vdd.n913 gnd 0.00713f
C3331 vdd.t127 gnd 0.267871f
C3332 vdd.t122 gnd 0.326802f
C3333 vdd.n914 gnd 0.00713f
C3334 vdd.n915 gnd 0.00713f
C3335 vdd.n916 gnd 0.00713f
C3336 vdd.t107 gnd 0.364304f
C3337 vdd.n917 gnd 0.00713f
C3338 vdd.n918 gnd 0.00713f
C3339 vdd.t106 gnd 0.364304f
C3340 vdd.n919 gnd 0.00713f
C3341 vdd.n920 gnd 0.00713f
C3342 vdd.n921 gnd 0.00713f
C3343 vdd.t101 gnd 0.364304f
C3344 vdd.n922 gnd 0.00713f
C3345 vdd.n923 gnd 0.00713f
C3346 vdd.t0 gnd 0.364304f
C3347 vdd.n924 gnd 0.00713f
C3348 vdd.n925 gnd 0.00713f
C3349 vdd.n926 gnd 0.00713f
C3350 vdd.n927 gnd 0.728608f
C3351 vdd.n928 gnd 0.00713f
C3352 vdd.n929 gnd 0.00713f
C3353 vdd.n930 gnd 0.503597f
C3354 vdd.n931 gnd 0.00713f
C3355 vdd.n932 gnd 0.00713f
C3356 vdd.n933 gnd 0.00713f
C3357 vdd.t132 gnd 0.364304f
C3358 vdd.n934 gnd 0.00713f
C3359 vdd.n935 gnd 0.00713f
C3360 vdd.n936 gnd 0.00713f
C3361 vdd.n937 gnd 0.00713f
C3362 vdd.n938 gnd 0.00713f
C3363 vdd.t3 gnd 0.364304f
C3364 vdd.n939 gnd 0.00713f
C3365 vdd.n940 gnd 0.00713f
C3366 vdd.t72 gnd 0.364304f
C3367 vdd.n941 gnd 0.00713f
C3368 vdd.n942 gnd 0.016433f
C3369 vdd.n943 gnd 0.016433f
C3370 vdd.t5 gnd 0.64289f
C3371 vdd.n944 gnd 0.015441f
C3372 vdd.n945 gnd 0.015441f
C3373 vdd.n946 gnd 0.407164f
C3374 vdd.n947 gnd 0.016433f
C3375 vdd.n948 gnd 0.00713f
C3376 vdd.n949 gnd 0.00713f
C3377 vdd.t139 gnd 0.64289f
C3378 vdd.n967 gnd 0.016433f
C3379 vdd.n985 gnd 0.015441f
C3380 vdd.n986 gnd 0.00713f
C3381 vdd.n987 gnd 0.015441f
C3382 vdd.t93 gnd 0.288105f
C3383 vdd.t92 gnd 0.294911f
C3384 vdd.t91 gnd 0.188086f
C3385 vdd.n988 gnd 0.10165f
C3386 vdd.n989 gnd 0.057659f
C3387 vdd.n990 gnd 0.016345f
C3388 vdd.n991 gnd 0.00713f
C3389 vdd.n992 gnd 0.407164f
C3390 vdd.n993 gnd 0.015441f
C3391 vdd.n994 gnd 0.00713f
C3392 vdd.n995 gnd 0.016433f
C3393 vdd.n996 gnd 0.00713f
C3394 vdd.t70 gnd 0.288105f
C3395 vdd.t69 gnd 0.294911f
C3396 vdd.t67 gnd 0.188086f
C3397 vdd.n997 gnd 0.10165f
C3398 vdd.n998 gnd 0.057659f
C3399 vdd.n999 gnd 0.010189f
C3400 vdd.n1000 gnd 0.00713f
C3401 vdd.n1001 gnd 0.00713f
C3402 vdd.t68 gnd 0.364304f
C3403 vdd.n1002 gnd 0.00713f
C3404 vdd.t137 gnd 0.364304f
C3405 vdd.n1003 gnd 0.00713f
C3406 vdd.n1004 gnd 0.00713f
C3407 vdd.n1005 gnd 0.00713f
C3408 vdd.n1006 gnd 0.00713f
C3409 vdd.n1007 gnd 0.00713f
C3410 vdd.n1008 gnd 0.728608f
C3411 vdd.n1009 gnd 0.00713f
C3412 vdd.n1010 gnd 0.00713f
C3413 vdd.t118 gnd 0.364304f
C3414 vdd.n1011 gnd 0.00713f
C3415 vdd.n1012 gnd 0.00713f
C3416 vdd.n1013 gnd 0.00713f
C3417 vdd.n1014 gnd 0.00713f
C3418 vdd.n1015 gnd 0.503597f
C3419 vdd.n1016 gnd 0.00713f
C3420 vdd.n1017 gnd 0.00713f
C3421 vdd.n1018 gnd 0.00713f
C3422 vdd.n1019 gnd 0.00713f
C3423 vdd.n1020 gnd 0.00713f
C3424 vdd.t131 gnd 0.364304f
C3425 vdd.n1021 gnd 0.00713f
C3426 vdd.n1022 gnd 0.00713f
C3427 vdd.t302 gnd 0.364304f
C3428 vdd.n1023 gnd 0.00713f
C3429 vdd.n1024 gnd 0.00713f
C3430 vdd.n1025 gnd 0.00713f
C3431 vdd.t20 gnd 0.364304f
C3432 vdd.n1026 gnd 0.00713f
C3433 vdd.n1027 gnd 0.00713f
C3434 vdd.t1 gnd 0.364304f
C3435 vdd.n1028 gnd 0.00713f
C3436 vdd.n1029 gnd 0.00713f
C3437 vdd.n1030 gnd 0.00713f
C3438 vdd.t103 gnd 0.326802f
C3439 vdd.n1031 gnd 0.00713f
C3440 vdd.n1032 gnd 0.00713f
C3441 vdd.n1033 gnd 0.562529f
C3442 vdd.n1034 gnd 0.00713f
C3443 vdd.n1035 gnd 0.00713f
C3444 vdd.n1036 gnd 0.00713f
C3445 vdd.t109 gnd 0.364304f
C3446 vdd.n1037 gnd 0.00713f
C3447 vdd.n1038 gnd 0.00713f
C3448 vdd.t105 gnd 0.267871f
C3449 vdd.n1039 gnd 0.401806f
C3450 vdd.n1040 gnd 0.00713f
C3451 vdd.n1041 gnd 0.00713f
C3452 vdd.n1042 gnd 0.00713f
C3453 vdd.n1043 gnd 0.648247f
C3454 vdd.n1044 gnd 0.00713f
C3455 vdd.n1045 gnd 0.00713f
C3456 vdd.t124 gnd 0.364304f
C3457 vdd.n1046 gnd 0.00713f
C3458 vdd.n1047 gnd 0.00713f
C3459 vdd.n1048 gnd 0.00713f
C3460 vdd.n1049 gnd 0.728608f
C3461 vdd.n1050 gnd 0.00713f
C3462 vdd.n1051 gnd 0.00713f
C3463 vdd.t11 gnd 0.364304f
C3464 vdd.n1052 gnd 0.00713f
C3465 vdd.n1053 gnd 0.00713f
C3466 vdd.n1054 gnd 0.00713f
C3467 vdd.t10 gnd 0.128578f
C3468 vdd.n1055 gnd 0.00713f
C3469 vdd.n1056 gnd 0.00713f
C3470 vdd.n1057 gnd 0.00713f
C3471 vdd.t83 gnd 0.294911f
C3472 vdd.t81 gnd 0.188086f
C3473 vdd.t84 gnd 0.294911f
C3474 vdd.n1058 gnd 0.165752f
C3475 vdd.n1059 gnd 0.00713f
C3476 vdd.n1060 gnd 0.00713f
C3477 vdd.t8 gnd 0.364304f
C3478 vdd.n1061 gnd 0.00713f
C3479 vdd.n1062 gnd 0.00713f
C3480 vdd.t82 gnd 0.283943f
C3481 vdd.n1063 gnd 0.600031f
C3482 vdd.n1064 gnd 0.00713f
C3483 vdd.n1065 gnd 0.00713f
C3484 vdd.n1066 gnd 0.00713f
C3485 vdd.n1067 gnd 0.401806f
C3486 vdd.n1068 gnd 0.00713f
C3487 vdd.n1069 gnd 0.00713f
C3488 vdd.n1070 gnd 0.487525f
C3489 vdd.n1071 gnd 0.00713f
C3490 vdd.n1072 gnd 0.00713f
C3491 vdd.n1073 gnd 0.00713f
C3492 vdd.n1074 gnd 0.562529f
C3493 vdd.n1075 gnd 0.00713f
C3494 vdd.n1076 gnd 0.00713f
C3495 vdd.t130 gnd 0.364304f
C3496 vdd.n1077 gnd 0.00713f
C3497 vdd.n1078 gnd 0.00713f
C3498 vdd.n1079 gnd 0.00713f
C3499 vdd.n1080 gnd 0.723251f
C3500 vdd.n1081 gnd 0.00713f
C3501 vdd.n1082 gnd 0.00713f
C3502 vdd.t19 gnd 0.364304f
C3503 vdd.n1083 gnd 0.00713f
C3504 vdd.n1084 gnd 0.00713f
C3505 vdd.n1085 gnd 0.00713f
C3506 vdd.n1086 gnd 0.728608f
C3507 vdd.n1087 gnd 0.00713f
C3508 vdd.n1088 gnd 0.00713f
C3509 vdd.t117 gnd 0.364304f
C3510 vdd.n1089 gnd 0.00713f
C3511 vdd.n1090 gnd 0.00713f
C3512 vdd.n1091 gnd 0.00713f
C3513 vdd.n1092 gnd 0.728608f
C3514 vdd.n1093 gnd 0.00713f
C3515 vdd.n1094 gnd 0.00713f
C3516 vdd.n1095 gnd 0.00713f
C3517 vdd.n1096 gnd 0.00713f
C3518 vdd.n1097 gnd 0.00713f
C3519 vdd.n1098 gnd 0.594673f
C3520 vdd.n1099 gnd 0.00713f
C3521 vdd.n1100 gnd 0.00713f
C3522 vdd.n1101 gnd 0.00713f
C3523 vdd.n1102 gnd 0.00713f
C3524 vdd.n1103 gnd 0.00713f
C3525 vdd.n1104 gnd 0.728608f
C3526 vdd.n1105 gnd 0.00713f
C3527 vdd.n1106 gnd 0.00713f
C3528 vdd.t30 gnd 0.364304f
C3529 vdd.n1107 gnd 0.00713f
C3530 vdd.n1108 gnd 0.016433f
C3531 vdd.n1109 gnd 0.016433f
C3532 vdd.n1110 gnd 10.897f
C3533 vdd.n1111 gnd 0.015441f
C3534 vdd.n1112 gnd 0.015441f
C3535 vdd.n1113 gnd 0.016433f
C3536 vdd.n1114 gnd 0.00713f
C3537 vdd.n1116 gnd 0.00713f
C3538 vdd.n1117 gnd 0.00713f
C3539 vdd.n1118 gnd 0.00713f
C3540 vdd.n1119 gnd 0.00713f
C3541 vdd.n1120 gnd 0.00713f
C3542 vdd.n1121 gnd 0.00713f
C3543 vdd.n1122 gnd 0.037513f
C3544 vdd.n1123 gnd 0.00713f
C3545 vdd.n1124 gnd 0.00713f
C3546 vdd.n1125 gnd 0.00713f
C3547 vdd.n1126 gnd 0.00713f
C3548 vdd.n1127 gnd 0.00713f
C3549 vdd.n1128 gnd 0.00713f
C3550 vdd.n1129 gnd 0.00713f
C3551 vdd.t95 gnd 0.288105f
C3552 vdd.t96 gnd 0.294911f
C3553 vdd.t94 gnd 0.188086f
C3554 vdd.n1130 gnd 0.10165f
C3555 vdd.n1131 gnd 0.057659f
C3556 vdd.n1132 gnd 0.00713f
C3557 vdd.n1133 gnd 0.00713f
C3558 vdd.n1134 gnd 0.00713f
C3559 vdd.n1135 gnd 0.00713f
C3560 vdd.t31 gnd 0.288105f
C3561 vdd.t32 gnd 0.294911f
C3562 vdd.t29 gnd 0.188086f
C3563 vdd.n1136 gnd 0.10165f
C3564 vdd.n1137 gnd 0.057659f
C3565 vdd.n1138 gnd 0.00713f
C3566 vdd.n1139 gnd 0.00713f
C3567 vdd.n1140 gnd 0.00713f
C3568 vdd.n1141 gnd 0.00713f
C3569 vdd.n1142 gnd 0.00713f
C3570 vdd.n1143 gnd 0.00713f
C3571 vdd.n1144 gnd 0.00671f
C3572 vdd.n1147 gnd 0.025907f
C3573 vdd.n1148 gnd 0.008439f
C3574 vdd.n1149 gnd 0.010485f
C3575 vdd.n1151 gnd 0.010485f
C3576 vdd.n1152 gnd 0.007004f
C3577 vdd.t48 gnd 0.535742f
C3578 vdd.n1153 gnd 11.304099f
C3579 vdd.n1154 gnd 0.010485f
C3580 vdd.n1155 gnd 0.025907f
C3581 vdd.n1156 gnd 0.008439f
C3582 vdd.n1157 gnd 0.010485f
C3583 vdd.n1158 gnd 0.008439f
C3584 vdd.n1159 gnd 0.010485f
C3585 vdd.n1160 gnd 1.07148f
C3586 vdd.n1161 gnd 0.010485f
C3587 vdd.n1162 gnd 0.008439f
C3588 vdd.n1163 gnd 0.008439f
C3589 vdd.n1164 gnd 0.010485f
C3590 vdd.n1165 gnd 0.008439f
C3591 vdd.n1166 gnd 0.010485f
C3592 vdd.t240 gnd 0.535742f
C3593 vdd.n1167 gnd 0.010485f
C3594 vdd.n1168 gnd 0.008439f
C3595 vdd.n1169 gnd 0.010485f
C3596 vdd.n1170 gnd 0.008439f
C3597 vdd.n1171 gnd 0.010485f
C3598 vdd.t153 gnd 0.535742f
C3599 vdd.n1172 gnd 0.010485f
C3600 vdd.n1173 gnd 0.008439f
C3601 vdd.n1174 gnd 0.010485f
C3602 vdd.n1175 gnd 0.008439f
C3603 vdd.n1176 gnd 0.010485f
C3604 vdd.n1177 gnd 0.862544f
C3605 vdd.n1178 gnd 0.889331f
C3606 vdd.t204 gnd 0.535742f
C3607 vdd.n1179 gnd 0.010485f
C3608 vdd.n1180 gnd 0.008439f
C3609 vdd.n1181 gnd 0.010485f
C3610 vdd.n1182 gnd 0.008439f
C3611 vdd.n1183 gnd 0.010485f
C3612 vdd.n1184 gnd 0.680392f
C3613 vdd.n1185 gnd 0.010485f
C3614 vdd.n1186 gnd 0.008439f
C3615 vdd.n1187 gnd 0.010485f
C3616 vdd.n1188 gnd 0.008439f
C3617 vdd.n1189 gnd 0.010485f
C3618 vdd.t234 gnd 0.535742f
C3619 vdd.t181 gnd 0.535742f
C3620 vdd.n1190 gnd 0.010485f
C3621 vdd.n1191 gnd 0.008439f
C3622 vdd.n1192 gnd 0.010485f
C3623 vdd.n1193 gnd 0.008439f
C3624 vdd.n1194 gnd 0.010485f
C3625 vdd.t238 gnd 0.535742f
C3626 vdd.n1195 gnd 0.010485f
C3627 vdd.n1196 gnd 0.008439f
C3628 vdd.n1197 gnd 0.010485f
C3629 vdd.n1198 gnd 0.008439f
C3630 vdd.n1199 gnd 0.010485f
C3631 vdd.t151 gnd 0.535742f
C3632 vdd.n1200 gnd 0.755396f
C3633 vdd.n1201 gnd 0.010485f
C3634 vdd.n1202 gnd 0.008439f
C3635 vdd.n1203 gnd 0.010485f
C3636 vdd.n1204 gnd 0.008439f
C3637 vdd.n1205 gnd 0.010485f
C3638 vdd.n1206 gnd 0.841114f
C3639 vdd.n1207 gnd 0.010485f
C3640 vdd.n1208 gnd 0.008439f
C3641 vdd.n1209 gnd 0.010485f
C3642 vdd.n1210 gnd 0.008439f
C3643 vdd.n1211 gnd 0.010485f
C3644 vdd.n1212 gnd 0.658962f
C3645 vdd.t178 gnd 0.535742f
C3646 vdd.n1213 gnd 0.010485f
C3647 vdd.n1214 gnd 0.008439f
C3648 vdd.n1215 gnd 0.010485f
C3649 vdd.n1216 gnd 0.008439f
C3650 vdd.n1217 gnd 0.010485f
C3651 vdd.t147 gnd 0.535742f
C3652 vdd.n1218 gnd 0.010485f
C3653 vdd.n1219 gnd 0.008439f
C3654 vdd.n1220 gnd 0.010485f
C3655 vdd.n1221 gnd 0.008439f
C3656 vdd.n1222 gnd 0.010485f
C3657 vdd.t206 gnd 0.535742f
C3658 vdd.n1223 gnd 0.594673f
C3659 vdd.n1224 gnd 0.010485f
C3660 vdd.n1225 gnd 0.008439f
C3661 vdd.n1226 gnd 0.010485f
C3662 vdd.n1227 gnd 0.008439f
C3663 vdd.n1228 gnd 0.010485f
C3664 vdd.t232 gnd 0.535742f
C3665 vdd.n1229 gnd 0.010485f
C3666 vdd.n1230 gnd 0.008439f
C3667 vdd.n1231 gnd 0.010485f
C3668 vdd.n1232 gnd 0.008439f
C3669 vdd.n1233 gnd 0.010485f
C3670 vdd.n1234 gnd 0.819685f
C3671 vdd.n1235 gnd 0.889331f
C3672 vdd.t141 gnd 0.535742f
C3673 vdd.n1236 gnd 0.010485f
C3674 vdd.n1237 gnd 0.008439f
C3675 vdd.n1238 gnd 0.010485f
C3676 vdd.n1239 gnd 0.008439f
C3677 vdd.n1240 gnd 0.010485f
C3678 vdd.n1241 gnd 0.637532f
C3679 vdd.n1242 gnd 0.010485f
C3680 vdd.n1243 gnd 0.008439f
C3681 vdd.n1244 gnd 0.010485f
C3682 vdd.n1245 gnd 0.008439f
C3683 vdd.n1246 gnd 0.010485f
C3684 vdd.t222 gnd 0.535742f
C3685 vdd.t253 gnd 0.535742f
C3686 vdd.n1247 gnd 0.010485f
C3687 vdd.n1248 gnd 0.008439f
C3688 vdd.n1249 gnd 0.010485f
C3689 vdd.n1250 gnd 0.008439f
C3690 vdd.n1251 gnd 0.010485f
C3691 vdd.t183 gnd 0.535742f
C3692 vdd.n1252 gnd 0.010485f
C3693 vdd.n1253 gnd 0.008439f
C3694 vdd.n1254 gnd 0.010485f
C3695 vdd.n1255 gnd 0.008439f
C3696 vdd.n1256 gnd 0.010485f
C3697 vdd.t236 gnd 0.535742f
C3698 vdd.n1257 gnd 0.798255f
C3699 vdd.n1258 gnd 0.010485f
C3700 vdd.n1259 gnd 0.008439f
C3701 vdd.n1260 gnd 0.010485f
C3702 vdd.n1261 gnd 0.008439f
C3703 vdd.n1262 gnd 0.010485f
C3704 vdd.n1263 gnd 1.07148f
C3705 vdd.n1264 gnd 0.010485f
C3706 vdd.n1265 gnd 0.008439f
C3707 vdd.n1266 gnd 0.025363f
C3708 vdd.n1267 gnd 0.007004f
C3709 vdd.n1268 gnd 0.025363f
C3710 vdd.t64 gnd 0.535742f
C3711 vdd.n1269 gnd 0.025363f
C3712 vdd.n1270 gnd 0.007004f
C3713 vdd.n1271 gnd 0.010485f
C3714 vdd.n1272 gnd 0.008439f
C3715 vdd.n1273 gnd 0.010485f
C3716 vdd.n1304 gnd 0.025907f
C3717 vdd.n1305 gnd 1.58044f
C3718 vdd.n1306 gnd 0.010485f
C3719 vdd.n1307 gnd 0.008439f
C3720 vdd.n1308 gnd 0.010485f
C3721 vdd.n1309 gnd 0.010485f
C3722 vdd.n1310 gnd 0.010485f
C3723 vdd.n1311 gnd 0.010485f
C3724 vdd.n1312 gnd 0.010485f
C3725 vdd.n1313 gnd 0.008439f
C3726 vdd.n1314 gnd 0.010485f
C3727 vdd.n1315 gnd 0.010485f
C3728 vdd.n1316 gnd 0.010485f
C3729 vdd.n1317 gnd 0.010485f
C3730 vdd.n1318 gnd 0.010485f
C3731 vdd.n1319 gnd 0.008439f
C3732 vdd.n1320 gnd 0.010485f
C3733 vdd.n1321 gnd 0.010485f
C3734 vdd.n1322 gnd 0.010485f
C3735 vdd.n1323 gnd 0.010485f
C3736 vdd.n1324 gnd 0.010485f
C3737 vdd.n1325 gnd 0.008439f
C3738 vdd.n1326 gnd 0.010485f
C3739 vdd.n1327 gnd 0.010485f
C3740 vdd.n1328 gnd 0.010485f
C3741 vdd.n1329 gnd 0.010485f
C3742 vdd.n1330 gnd 0.010485f
C3743 vdd.t89 gnd 0.128989f
C3744 vdd.t90 gnd 0.137854f
C3745 vdd.t88 gnd 0.168458f
C3746 vdd.n1331 gnd 0.215939f
C3747 vdd.n1332 gnd 0.182272f
C3748 vdd.n1333 gnd 0.018059f
C3749 vdd.n1334 gnd 0.010485f
C3750 vdd.n1335 gnd 0.010485f
C3751 vdd.n1336 gnd 0.010485f
C3752 vdd.n1337 gnd 0.010485f
C3753 vdd.n1338 gnd 0.010485f
C3754 vdd.n1339 gnd 0.008439f
C3755 vdd.n1340 gnd 0.010485f
C3756 vdd.n1341 gnd 0.010485f
C3757 vdd.n1342 gnd 0.010485f
C3758 vdd.n1343 gnd 0.010485f
C3759 vdd.n1344 gnd 0.010485f
C3760 vdd.n1345 gnd 0.008439f
C3761 vdd.n1346 gnd 0.010485f
C3762 vdd.n1347 gnd 0.010485f
C3763 vdd.n1348 gnd 0.010485f
C3764 vdd.n1349 gnd 0.010485f
C3765 vdd.n1350 gnd 0.010485f
C3766 vdd.n1351 gnd 0.008439f
C3767 vdd.n1352 gnd 0.010485f
C3768 vdd.n1353 gnd 0.010485f
C3769 vdd.n1354 gnd 0.010485f
C3770 vdd.n1355 gnd 0.010485f
C3771 vdd.n1356 gnd 0.010485f
C3772 vdd.n1357 gnd 0.008439f
C3773 vdd.n1358 gnd 0.010485f
C3774 vdd.n1359 gnd 0.010485f
C3775 vdd.n1360 gnd 0.010485f
C3776 vdd.n1361 gnd 0.010485f
C3777 vdd.n1362 gnd 0.010485f
C3778 vdd.n1363 gnd 0.008439f
C3779 vdd.n1364 gnd 0.010485f
C3780 vdd.n1365 gnd 0.010485f
C3781 vdd.n1366 gnd 0.010485f
C3782 vdd.n1367 gnd 0.010485f
C3783 vdd.n1368 gnd 0.008439f
C3784 vdd.n1369 gnd 0.010485f
C3785 vdd.n1370 gnd 0.010485f
C3786 vdd.n1371 gnd 0.010485f
C3787 vdd.n1372 gnd 0.010485f
C3788 vdd.n1373 gnd 0.010485f
C3789 vdd.n1374 gnd 0.008439f
C3790 vdd.n1375 gnd 0.010485f
C3791 vdd.n1376 gnd 0.010485f
C3792 vdd.n1377 gnd 0.010485f
C3793 vdd.n1378 gnd 0.010485f
C3794 vdd.n1379 gnd 0.010485f
C3795 vdd.n1380 gnd 0.008439f
C3796 vdd.n1381 gnd 0.010485f
C3797 vdd.n1382 gnd 0.010485f
C3798 vdd.n1383 gnd 0.010485f
C3799 vdd.n1384 gnd 0.010485f
C3800 vdd.n1385 gnd 0.010485f
C3801 vdd.n1386 gnd 0.008439f
C3802 vdd.n1387 gnd 0.010485f
C3803 vdd.n1388 gnd 0.010485f
C3804 vdd.n1389 gnd 0.010485f
C3805 vdd.n1390 gnd 0.010485f
C3806 vdd.n1391 gnd 0.010485f
C3807 vdd.n1392 gnd 0.008439f
C3808 vdd.n1393 gnd 0.010485f
C3809 vdd.n1394 gnd 0.010485f
C3810 vdd.n1395 gnd 0.010485f
C3811 vdd.n1396 gnd 0.010485f
C3812 vdd.t65 gnd 0.128989f
C3813 vdd.t66 gnd 0.137854f
C3814 vdd.t63 gnd 0.168458f
C3815 vdd.n1397 gnd 0.215939f
C3816 vdd.n1398 gnd 0.182272f
C3817 vdd.n1399 gnd 0.01384f
C3818 vdd.n1400 gnd 0.004008f
C3819 vdd.n1401 gnd 0.025907f
C3820 vdd.n1402 gnd 0.010485f
C3821 vdd.n1403 gnd 0.00443f
C3822 vdd.n1404 gnd 0.008439f
C3823 vdd.n1405 gnd 0.008439f
C3824 vdd.n1406 gnd 0.010485f
C3825 vdd.n1407 gnd 0.010485f
C3826 vdd.n1408 gnd 0.010485f
C3827 vdd.n1409 gnd 0.008439f
C3828 vdd.n1410 gnd 0.008439f
C3829 vdd.n1411 gnd 0.008439f
C3830 vdd.n1412 gnd 0.010485f
C3831 vdd.n1413 gnd 0.010485f
C3832 vdd.n1414 gnd 0.010485f
C3833 vdd.n1415 gnd 0.008439f
C3834 vdd.n1416 gnd 0.008439f
C3835 vdd.n1417 gnd 0.008439f
C3836 vdd.n1418 gnd 0.010485f
C3837 vdd.n1419 gnd 0.010485f
C3838 vdd.n1420 gnd 0.010485f
C3839 vdd.n1421 gnd 0.008439f
C3840 vdd.n1422 gnd 0.008439f
C3841 vdd.n1423 gnd 0.008439f
C3842 vdd.n1424 gnd 0.010485f
C3843 vdd.n1425 gnd 0.010485f
C3844 vdd.n1426 gnd 0.010485f
C3845 vdd.n1427 gnd 0.008439f
C3846 vdd.n1428 gnd 0.008439f
C3847 vdd.n1429 gnd 0.008439f
C3848 vdd.n1430 gnd 0.010485f
C3849 vdd.n1431 gnd 0.010485f
C3850 vdd.n1432 gnd 0.010485f
C3851 vdd.n1433 gnd 0.008354f
C3852 vdd.n1434 gnd 0.010485f
C3853 vdd.t76 gnd 0.128989f
C3854 vdd.t77 gnd 0.137854f
C3855 vdd.t75 gnd 0.168458f
C3856 vdd.n1435 gnd 0.215939f
C3857 vdd.n1436 gnd 0.182272f
C3858 vdd.n1437 gnd 0.018059f
C3859 vdd.n1438 gnd 0.005738f
C3860 vdd.n1439 gnd 0.010485f
C3861 vdd.n1440 gnd 0.010485f
C3862 vdd.n1441 gnd 0.010485f
C3863 vdd.n1442 gnd 0.008439f
C3864 vdd.n1443 gnd 0.008439f
C3865 vdd.n1444 gnd 0.008439f
C3866 vdd.n1445 gnd 0.010485f
C3867 vdd.n1446 gnd 0.010485f
C3868 vdd.n1447 gnd 0.010485f
C3869 vdd.n1448 gnd 0.008439f
C3870 vdd.n1449 gnd 0.008439f
C3871 vdd.n1450 gnd 0.008439f
C3872 vdd.n1451 gnd 0.010485f
C3873 vdd.n1452 gnd 0.010485f
C3874 vdd.n1453 gnd 0.010485f
C3875 vdd.n1454 gnd 0.008439f
C3876 vdd.n1455 gnd 0.008439f
C3877 vdd.n1456 gnd 0.008439f
C3878 vdd.n1457 gnd 0.010485f
C3879 vdd.n1458 gnd 0.010485f
C3880 vdd.n1459 gnd 0.010485f
C3881 vdd.n1460 gnd 0.008439f
C3882 vdd.n1461 gnd 0.008439f
C3883 vdd.n1462 gnd 0.008439f
C3884 vdd.n1463 gnd 0.010485f
C3885 vdd.n1464 gnd 0.010485f
C3886 vdd.n1465 gnd 0.010485f
C3887 vdd.n1466 gnd 0.008439f
C3888 vdd.n1467 gnd 0.008439f
C3889 vdd.n1468 gnd 0.007046f
C3890 vdd.n1469 gnd 0.010485f
C3891 vdd.n1470 gnd 0.010485f
C3892 vdd.n1471 gnd 0.010485f
C3893 vdd.n1472 gnd 0.007046f
C3894 vdd.n1473 gnd 0.008439f
C3895 vdd.n1474 gnd 0.008439f
C3896 vdd.n1475 gnd 0.010485f
C3897 vdd.n1476 gnd 0.010485f
C3898 vdd.n1477 gnd 0.010485f
C3899 vdd.n1478 gnd 0.008439f
C3900 vdd.n1479 gnd 0.008439f
C3901 vdd.n1480 gnd 0.008439f
C3902 vdd.n1481 gnd 0.010485f
C3903 vdd.n1482 gnd 0.010485f
C3904 vdd.n1483 gnd 0.010485f
C3905 vdd.n1484 gnd 0.008439f
C3906 vdd.n1485 gnd 0.008439f
C3907 vdd.n1486 gnd 0.008439f
C3908 vdd.n1487 gnd 0.010485f
C3909 vdd.n1488 gnd 0.010485f
C3910 vdd.n1489 gnd 0.010485f
C3911 vdd.n1490 gnd 0.008439f
C3912 vdd.n1491 gnd 0.008439f
C3913 vdd.n1492 gnd 0.008439f
C3914 vdd.n1493 gnd 0.010485f
C3915 vdd.n1494 gnd 0.010485f
C3916 vdd.n1495 gnd 0.010485f
C3917 vdd.n1496 gnd 0.008439f
C3918 vdd.n1497 gnd 0.010485f
C3919 vdd.n1498 gnd 2.53941f
C3920 vdd.n1500 gnd 0.025907f
C3921 vdd.n1501 gnd 0.007004f
C3922 vdd.n1502 gnd 0.025907f
C3923 vdd.n1503 gnd 0.025363f
C3924 vdd.n1504 gnd 0.010485f
C3925 vdd.n1505 gnd 0.008439f
C3926 vdd.n1506 gnd 0.010485f
C3927 vdd.n1507 gnd 0.541099f
C3928 vdd.n1508 gnd 0.010485f
C3929 vdd.n1509 gnd 0.008439f
C3930 vdd.n1510 gnd 0.010485f
C3931 vdd.n1511 gnd 0.010485f
C3932 vdd.n1512 gnd 0.010485f
C3933 vdd.n1513 gnd 0.008439f
C3934 vdd.n1514 gnd 0.010485f
C3935 vdd.n1515 gnd 0.980407f
C3936 vdd.n1516 gnd 1.07148f
C3937 vdd.n1517 gnd 0.010485f
C3938 vdd.n1518 gnd 0.008439f
C3939 vdd.n1519 gnd 0.010485f
C3940 vdd.n1520 gnd 0.010485f
C3941 vdd.n1521 gnd 0.010485f
C3942 vdd.n1522 gnd 0.008439f
C3943 vdd.n1523 gnd 0.010485f
C3944 vdd.n1524 gnd 0.626818f
C3945 vdd.n1525 gnd 0.010485f
C3946 vdd.n1526 gnd 0.008439f
C3947 vdd.n1527 gnd 0.010485f
C3948 vdd.n1528 gnd 0.010485f
C3949 vdd.n1529 gnd 0.010485f
C3950 vdd.n1530 gnd 0.008439f
C3951 vdd.n1531 gnd 0.010485f
C3952 vdd.n1532 gnd 0.616103f
C3953 vdd.n1533 gnd 0.80897f
C3954 vdd.n1534 gnd 0.010485f
C3955 vdd.n1535 gnd 0.008439f
C3956 vdd.n1536 gnd 0.010485f
C3957 vdd.n1537 gnd 0.010485f
C3958 vdd.n1538 gnd 0.010485f
C3959 vdd.n1539 gnd 0.008439f
C3960 vdd.n1540 gnd 0.010485f
C3961 vdd.n1541 gnd 0.889331f
C3962 vdd.n1542 gnd 0.010485f
C3963 vdd.n1543 gnd 0.008439f
C3964 vdd.n1544 gnd 0.010485f
C3965 vdd.n1545 gnd 0.010485f
C3966 vdd.n1546 gnd 0.010485f
C3967 vdd.n1547 gnd 0.008439f
C3968 vdd.n1548 gnd 0.010485f
C3969 vdd.t194 gnd 0.535742f
C3970 vdd.n1549 gnd 0.78754f
C3971 vdd.n1550 gnd 0.010485f
C3972 vdd.n1551 gnd 0.008439f
C3973 vdd.n1552 gnd 0.010485f
C3974 vdd.n1553 gnd 0.010485f
C3975 vdd.n1554 gnd 0.010485f
C3976 vdd.n1555 gnd 0.008439f
C3977 vdd.n1556 gnd 0.010485f
C3978 vdd.n1557 gnd 0.605388f
C3979 vdd.n1558 gnd 0.010485f
C3980 vdd.n1559 gnd 0.008439f
C3981 vdd.n1560 gnd 0.010485f
C3982 vdd.n1561 gnd 0.010485f
C3983 vdd.n1562 gnd 0.010485f
C3984 vdd.n1563 gnd 0.008439f
C3985 vdd.n1564 gnd 0.010485f
C3986 vdd.n1565 gnd 0.776825f
C3987 vdd.n1566 gnd 0.648247f
C3988 vdd.n1567 gnd 0.010485f
C3989 vdd.n1568 gnd 0.008439f
C3990 vdd.n1569 gnd 0.010485f
C3991 vdd.n1570 gnd 0.010485f
C3992 vdd.n1571 gnd 0.010485f
C3993 vdd.n1572 gnd 0.008439f
C3994 vdd.n1573 gnd 0.010485f
C3995 vdd.n1574 gnd 0.830399f
C3996 vdd.n1575 gnd 0.010485f
C3997 vdd.n1576 gnd 0.008439f
C3998 vdd.n1577 gnd 0.010485f
C3999 vdd.n1578 gnd 0.010485f
C4000 vdd.n1579 gnd 0.010485f
C4001 vdd.n1580 gnd 0.008439f
C4002 vdd.n1581 gnd 0.010485f
C4003 vdd.t143 gnd 0.535742f
C4004 vdd.n1582 gnd 0.889331f
C4005 vdd.n1583 gnd 0.010485f
C4006 vdd.n1584 gnd 0.008439f
C4007 vdd.n1585 gnd 0.010485f
C4008 vdd.n1586 gnd 0.008058f
C4009 vdd.n1587 gnd 0.005754f
C4010 vdd.n1588 gnd 0.00534f
C4011 vdd.n1589 gnd 0.002954f
C4012 vdd.n1590 gnd 0.006782f
C4013 vdd.n1591 gnd 0.002869f
C4014 vdd.n1592 gnd 0.003038f
C4015 vdd.n1593 gnd 0.00534f
C4016 vdd.n1594 gnd 0.002869f
C4017 vdd.n1595 gnd 0.006782f
C4018 vdd.n1596 gnd 0.003038f
C4019 vdd.n1597 gnd 0.00534f
C4020 vdd.n1598 gnd 0.002869f
C4021 vdd.n1599 gnd 0.005086f
C4022 vdd.n1600 gnd 0.005102f
C4023 vdd.t241 gnd 0.01457f
C4024 vdd.n1601 gnd 0.032418f
C4025 vdd.n1602 gnd 0.168712f
C4026 vdd.n1603 gnd 0.002869f
C4027 vdd.n1604 gnd 0.003038f
C4028 vdd.n1605 gnd 0.006782f
C4029 vdd.n1606 gnd 0.006782f
C4030 vdd.n1607 gnd 0.003038f
C4031 vdd.n1608 gnd 0.002869f
C4032 vdd.n1609 gnd 0.00534f
C4033 vdd.n1610 gnd 0.00534f
C4034 vdd.n1611 gnd 0.002869f
C4035 vdd.n1612 gnd 0.003038f
C4036 vdd.n1613 gnd 0.006782f
C4037 vdd.n1614 gnd 0.006782f
C4038 vdd.n1615 gnd 0.003038f
C4039 vdd.n1616 gnd 0.002869f
C4040 vdd.n1617 gnd 0.00534f
C4041 vdd.n1618 gnd 0.00534f
C4042 vdd.n1619 gnd 0.002869f
C4043 vdd.n1620 gnd 0.003038f
C4044 vdd.n1621 gnd 0.006782f
C4045 vdd.n1622 gnd 0.006782f
C4046 vdd.n1623 gnd 0.016034f
C4047 vdd.n1624 gnd 0.002954f
C4048 vdd.n1625 gnd 0.002869f
C4049 vdd.n1626 gnd 0.013801f
C4050 vdd.n1627 gnd 0.009635f
C4051 vdd.t205 gnd 0.033756f
C4052 vdd.t154 gnd 0.033756f
C4053 vdd.n1628 gnd 0.231991f
C4054 vdd.n1629 gnd 0.182426f
C4055 vdd.t229 gnd 0.033756f
C4056 vdd.t167 gnd 0.033756f
C4057 vdd.n1630 gnd 0.231991f
C4058 vdd.n1631 gnd 0.147217f
C4059 vdd.t277 gnd 0.033756f
C4060 vdd.t299 gnd 0.033756f
C4061 vdd.n1632 gnd 0.231991f
C4062 vdd.n1633 gnd 0.147217f
C4063 vdd.t258 gnd 0.033756f
C4064 vdd.t170 gnd 0.033756f
C4065 vdd.n1634 gnd 0.231991f
C4066 vdd.n1635 gnd 0.147217f
C4067 vdd.t243 gnd 0.033756f
C4068 vdd.t179 gnd 0.033756f
C4069 vdd.n1636 gnd 0.231991f
C4070 vdd.n1637 gnd 0.147217f
C4071 vdd.t287 gnd 0.033756f
C4072 vdd.t212 gnd 0.033756f
C4073 vdd.n1638 gnd 0.231991f
C4074 vdd.n1639 gnd 0.147217f
C4075 vdd.t264 gnd 0.033756f
C4076 vdd.t233 gnd 0.033756f
C4077 vdd.n1640 gnd 0.231991f
C4078 vdd.n1641 gnd 0.147217f
C4079 vdd.t279 gnd 0.033756f
C4080 vdd.t195 gnd 0.033756f
C4081 vdd.n1642 gnd 0.231991f
C4082 vdd.n1643 gnd 0.147217f
C4083 vdd.t295 gnd 0.033756f
C4084 vdd.t223 gnd 0.033756f
C4085 vdd.n1644 gnd 0.231991f
C4086 vdd.n1645 gnd 0.147217f
C4087 vdd.n1646 gnd 0.005754f
C4088 vdd.n1647 gnd 0.00534f
C4089 vdd.n1648 gnd 0.002954f
C4090 vdd.n1649 gnd 0.006782f
C4091 vdd.n1650 gnd 0.002869f
C4092 vdd.n1651 gnd 0.003038f
C4093 vdd.n1652 gnd 0.00534f
C4094 vdd.n1653 gnd 0.002869f
C4095 vdd.n1654 gnd 0.006782f
C4096 vdd.n1655 gnd 0.003038f
C4097 vdd.n1656 gnd 0.00534f
C4098 vdd.n1657 gnd 0.002869f
C4099 vdd.n1658 gnd 0.005086f
C4100 vdd.n1659 gnd 0.005102f
C4101 vdd.t246 gnd 0.01457f
C4102 vdd.n1660 gnd 0.032418f
C4103 vdd.n1661 gnd 0.168712f
C4104 vdd.n1662 gnd 0.002869f
C4105 vdd.n1663 gnd 0.003038f
C4106 vdd.n1664 gnd 0.006782f
C4107 vdd.n1665 gnd 0.006782f
C4108 vdd.n1666 gnd 0.003038f
C4109 vdd.n1667 gnd 0.002869f
C4110 vdd.n1668 gnd 0.00534f
C4111 vdd.n1669 gnd 0.00534f
C4112 vdd.n1670 gnd 0.002869f
C4113 vdd.n1671 gnd 0.003038f
C4114 vdd.n1672 gnd 0.006782f
C4115 vdd.n1673 gnd 0.006782f
C4116 vdd.n1674 gnd 0.003038f
C4117 vdd.n1675 gnd 0.002869f
C4118 vdd.n1676 gnd 0.00534f
C4119 vdd.n1677 gnd 0.00534f
C4120 vdd.n1678 gnd 0.002869f
C4121 vdd.n1679 gnd 0.003038f
C4122 vdd.n1680 gnd 0.006782f
C4123 vdd.n1681 gnd 0.006782f
C4124 vdd.n1682 gnd 0.016034f
C4125 vdd.n1683 gnd 0.002954f
C4126 vdd.n1684 gnd 0.002869f
C4127 vdd.n1685 gnd 0.013801f
C4128 vdd.n1686 gnd 0.009333f
C4129 vdd.n1687 gnd 0.10953f
C4130 vdd.n1688 gnd 0.005754f
C4131 vdd.n1689 gnd 0.00534f
C4132 vdd.n1690 gnd 0.002954f
C4133 vdd.n1691 gnd 0.006782f
C4134 vdd.n1692 gnd 0.002869f
C4135 vdd.n1693 gnd 0.003038f
C4136 vdd.n1694 gnd 0.00534f
C4137 vdd.n1695 gnd 0.002869f
C4138 vdd.n1696 gnd 0.006782f
C4139 vdd.n1697 gnd 0.003038f
C4140 vdd.n1698 gnd 0.00534f
C4141 vdd.n1699 gnd 0.002869f
C4142 vdd.n1700 gnd 0.005086f
C4143 vdd.n1701 gnd 0.005102f
C4144 vdd.t288 gnd 0.01457f
C4145 vdd.n1702 gnd 0.032418f
C4146 vdd.n1703 gnd 0.168712f
C4147 vdd.n1704 gnd 0.002869f
C4148 vdd.n1705 gnd 0.003038f
C4149 vdd.n1706 gnd 0.006782f
C4150 vdd.n1707 gnd 0.006782f
C4151 vdd.n1708 gnd 0.003038f
C4152 vdd.n1709 gnd 0.002869f
C4153 vdd.n1710 gnd 0.00534f
C4154 vdd.n1711 gnd 0.00534f
C4155 vdd.n1712 gnd 0.002869f
C4156 vdd.n1713 gnd 0.003038f
C4157 vdd.n1714 gnd 0.006782f
C4158 vdd.n1715 gnd 0.006782f
C4159 vdd.n1716 gnd 0.003038f
C4160 vdd.n1717 gnd 0.002869f
C4161 vdd.n1718 gnd 0.00534f
C4162 vdd.n1719 gnd 0.00534f
C4163 vdd.n1720 gnd 0.002869f
C4164 vdd.n1721 gnd 0.003038f
C4165 vdd.n1722 gnd 0.006782f
C4166 vdd.n1723 gnd 0.006782f
C4167 vdd.n1724 gnd 0.016034f
C4168 vdd.n1725 gnd 0.002954f
C4169 vdd.n1726 gnd 0.002869f
C4170 vdd.n1727 gnd 0.013801f
C4171 vdd.n1728 gnd 0.009635f
C4172 vdd.t252 gnd 0.033756f
C4173 vdd.t186 gnd 0.033756f
C4174 vdd.n1729 gnd 0.231991f
C4175 vdd.n1730 gnd 0.182426f
C4176 vdd.t182 gnd 0.033756f
C4177 vdd.t255 gnd 0.033756f
C4178 vdd.n1731 gnd 0.231991f
C4179 vdd.n1732 gnd 0.147217f
C4180 vdd.t239 gnd 0.033756f
C4181 vdd.t235 gnd 0.033756f
C4182 vdd.n1733 gnd 0.231991f
C4183 vdd.n1734 gnd 0.147217f
C4184 vdd.t177 gnd 0.033756f
C4185 vdd.t152 gnd 0.033756f
C4186 vdd.n1735 gnd 0.231991f
C4187 vdd.n1736 gnd 0.147217f
C4188 vdd.t144 gnd 0.033756f
C4189 vdd.t230 gnd 0.033756f
C4190 vdd.n1737 gnd 0.231991f
C4191 vdd.n1738 gnd 0.147217f
C4192 vdd.t207 gnd 0.033756f
C4193 vdd.t148 gnd 0.033756f
C4194 vdd.n1739 gnd 0.231991f
C4195 vdd.n1740 gnd 0.147217f
C4196 vdd.t142 gnd 0.033756f
C4197 vdd.t259 gnd 0.033756f
C4198 vdd.n1741 gnd 0.231991f
C4199 vdd.n1742 gnd 0.147217f
C4200 vdd.t254 gnd 0.033756f
C4201 vdd.t197 gnd 0.033756f
C4202 vdd.n1743 gnd 0.231991f
C4203 vdd.n1744 gnd 0.147217f
C4204 vdd.t184 gnd 0.033756f
C4205 vdd.t285 gnd 0.033756f
C4206 vdd.n1745 gnd 0.231991f
C4207 vdd.n1746 gnd 0.147217f
C4208 vdd.n1747 gnd 0.005754f
C4209 vdd.n1748 gnd 0.00534f
C4210 vdd.n1749 gnd 0.002954f
C4211 vdd.n1750 gnd 0.006782f
C4212 vdd.n1751 gnd 0.002869f
C4213 vdd.n1752 gnd 0.003038f
C4214 vdd.n1753 gnd 0.00534f
C4215 vdd.n1754 gnd 0.002869f
C4216 vdd.n1755 gnd 0.006782f
C4217 vdd.n1756 gnd 0.003038f
C4218 vdd.n1757 gnd 0.00534f
C4219 vdd.n1758 gnd 0.002869f
C4220 vdd.n1759 gnd 0.005086f
C4221 vdd.n1760 gnd 0.005102f
C4222 vdd.t237 gnd 0.01457f
C4223 vdd.n1761 gnd 0.032418f
C4224 vdd.n1762 gnd 0.168712f
C4225 vdd.n1763 gnd 0.002869f
C4226 vdd.n1764 gnd 0.003038f
C4227 vdd.n1765 gnd 0.006782f
C4228 vdd.n1766 gnd 0.006782f
C4229 vdd.n1767 gnd 0.003038f
C4230 vdd.n1768 gnd 0.002869f
C4231 vdd.n1769 gnd 0.00534f
C4232 vdd.n1770 gnd 0.00534f
C4233 vdd.n1771 gnd 0.002869f
C4234 vdd.n1772 gnd 0.003038f
C4235 vdd.n1773 gnd 0.006782f
C4236 vdd.n1774 gnd 0.006782f
C4237 vdd.n1775 gnd 0.003038f
C4238 vdd.n1776 gnd 0.002869f
C4239 vdd.n1777 gnd 0.00534f
C4240 vdd.n1778 gnd 0.00534f
C4241 vdd.n1779 gnd 0.002869f
C4242 vdd.n1780 gnd 0.003038f
C4243 vdd.n1781 gnd 0.006782f
C4244 vdd.n1782 gnd 0.006782f
C4245 vdd.n1783 gnd 0.016034f
C4246 vdd.n1784 gnd 0.002954f
C4247 vdd.n1785 gnd 0.002869f
C4248 vdd.n1786 gnd 0.013801f
C4249 vdd.n1787 gnd 0.009333f
C4250 vdd.n1788 gnd 0.065159f
C4251 vdd.n1789 gnd 0.234786f
C4252 vdd.n1790 gnd 0.005754f
C4253 vdd.n1791 gnd 0.00534f
C4254 vdd.n1792 gnd 0.002954f
C4255 vdd.n1793 gnd 0.006782f
C4256 vdd.n1794 gnd 0.002869f
C4257 vdd.n1795 gnd 0.003038f
C4258 vdd.n1796 gnd 0.00534f
C4259 vdd.n1797 gnd 0.002869f
C4260 vdd.n1798 gnd 0.006782f
C4261 vdd.n1799 gnd 0.003038f
C4262 vdd.n1800 gnd 0.00534f
C4263 vdd.n1801 gnd 0.002869f
C4264 vdd.n1802 gnd 0.005086f
C4265 vdd.n1803 gnd 0.005102f
C4266 vdd.t300 gnd 0.01457f
C4267 vdd.n1804 gnd 0.032418f
C4268 vdd.n1805 gnd 0.168712f
C4269 vdd.n1806 gnd 0.002869f
C4270 vdd.n1807 gnd 0.003038f
C4271 vdd.n1808 gnd 0.006782f
C4272 vdd.n1809 gnd 0.006782f
C4273 vdd.n1810 gnd 0.003038f
C4274 vdd.n1811 gnd 0.002869f
C4275 vdd.n1812 gnd 0.00534f
C4276 vdd.n1813 gnd 0.00534f
C4277 vdd.n1814 gnd 0.002869f
C4278 vdd.n1815 gnd 0.003038f
C4279 vdd.n1816 gnd 0.006782f
C4280 vdd.n1817 gnd 0.006782f
C4281 vdd.n1818 gnd 0.003038f
C4282 vdd.n1819 gnd 0.002869f
C4283 vdd.n1820 gnd 0.00534f
C4284 vdd.n1821 gnd 0.00534f
C4285 vdd.n1822 gnd 0.002869f
C4286 vdd.n1823 gnd 0.003038f
C4287 vdd.n1824 gnd 0.006782f
C4288 vdd.n1825 gnd 0.006782f
C4289 vdd.n1826 gnd 0.016034f
C4290 vdd.n1827 gnd 0.002954f
C4291 vdd.n1828 gnd 0.002869f
C4292 vdd.n1829 gnd 0.013801f
C4293 vdd.n1830 gnd 0.009635f
C4294 vdd.t266 gnd 0.033756f
C4295 vdd.t213 gnd 0.033756f
C4296 vdd.n1831 gnd 0.231991f
C4297 vdd.n1832 gnd 0.182426f
C4298 vdd.t208 gnd 0.033756f
C4299 vdd.t268 gnd 0.033756f
C4300 vdd.n1833 gnd 0.231991f
C4301 vdd.n1834 gnd 0.147217f
C4302 vdd.t250 gnd 0.033756f
C4303 vdd.t248 gnd 0.033756f
C4304 vdd.n1835 gnd 0.231991f
C4305 vdd.n1836 gnd 0.147217f
C4306 vdd.t203 gnd 0.033756f
C4307 vdd.t173 gnd 0.033756f
C4308 vdd.n1837 gnd 0.231991f
C4309 vdd.n1838 gnd 0.147217f
C4310 vdd.t171 gnd 0.033756f
C4311 vdd.t247 gnd 0.033756f
C4312 vdd.n1839 gnd 0.231991f
C4313 vdd.n1840 gnd 0.147217f
C4314 vdd.t224 gnd 0.033756f
C4315 vdd.t172 gnd 0.033756f
C4316 vdd.n1841 gnd 0.231991f
C4317 vdd.n1842 gnd 0.147217f
C4318 vdd.t165 gnd 0.033756f
C4319 vdd.t269 gnd 0.033756f
C4320 vdd.n1843 gnd 0.231991f
C4321 vdd.n1844 gnd 0.147217f
C4322 vdd.t267 gnd 0.033756f
C4323 vdd.t217 gnd 0.033756f
C4324 vdd.n1845 gnd 0.231991f
C4325 vdd.n1846 gnd 0.147217f
C4326 vdd.t209 gnd 0.033756f
C4327 vdd.t296 gnd 0.033756f
C4328 vdd.n1847 gnd 0.231991f
C4329 vdd.n1848 gnd 0.147217f
C4330 vdd.n1849 gnd 0.005754f
C4331 vdd.n1850 gnd 0.00534f
C4332 vdd.n1851 gnd 0.002954f
C4333 vdd.n1852 gnd 0.006782f
C4334 vdd.n1853 gnd 0.002869f
C4335 vdd.n1854 gnd 0.003038f
C4336 vdd.n1855 gnd 0.00534f
C4337 vdd.n1856 gnd 0.002869f
C4338 vdd.n1857 gnd 0.006782f
C4339 vdd.n1858 gnd 0.003038f
C4340 vdd.n1859 gnd 0.00534f
C4341 vdd.n1860 gnd 0.002869f
C4342 vdd.n1861 gnd 0.005086f
C4343 vdd.n1862 gnd 0.005102f
C4344 vdd.t249 gnd 0.01457f
C4345 vdd.n1863 gnd 0.032418f
C4346 vdd.n1864 gnd 0.168712f
C4347 vdd.n1865 gnd 0.002869f
C4348 vdd.n1866 gnd 0.003038f
C4349 vdd.n1867 gnd 0.006782f
C4350 vdd.n1868 gnd 0.006782f
C4351 vdd.n1869 gnd 0.003038f
C4352 vdd.n1870 gnd 0.002869f
C4353 vdd.n1871 gnd 0.00534f
C4354 vdd.n1872 gnd 0.00534f
C4355 vdd.n1873 gnd 0.002869f
C4356 vdd.n1874 gnd 0.003038f
C4357 vdd.n1875 gnd 0.006782f
C4358 vdd.n1876 gnd 0.006782f
C4359 vdd.n1877 gnd 0.003038f
C4360 vdd.n1878 gnd 0.002869f
C4361 vdd.n1879 gnd 0.00534f
C4362 vdd.n1880 gnd 0.00534f
C4363 vdd.n1881 gnd 0.002869f
C4364 vdd.n1882 gnd 0.003038f
C4365 vdd.n1883 gnd 0.006782f
C4366 vdd.n1884 gnd 0.006782f
C4367 vdd.n1885 gnd 0.016034f
C4368 vdd.n1886 gnd 0.002954f
C4369 vdd.n1887 gnd 0.002869f
C4370 vdd.n1888 gnd 0.013801f
C4371 vdd.n1889 gnd 0.009333f
C4372 vdd.n1890 gnd 0.065159f
C4373 vdd.n1891 gnd 0.268779f
C4374 vdd.n1892 gnd 2.94641f
C4375 vdd.n1893 gnd 0.618425f
C4376 vdd.n1894 gnd 0.008058f
C4377 vdd.n1895 gnd 0.008439f
C4378 vdd.n1896 gnd 0.010485f
C4379 vdd.n1897 gnd 0.76611f
C4380 vdd.n1898 gnd 0.010485f
C4381 vdd.n1899 gnd 0.008439f
C4382 vdd.n1900 gnd 0.010485f
C4383 vdd.n1901 gnd 0.010485f
C4384 vdd.n1902 gnd 0.010485f
C4385 vdd.n1903 gnd 0.008439f
C4386 vdd.n1904 gnd 0.010485f
C4387 vdd.n1905 gnd 0.889331f
C4388 vdd.t176 gnd 0.535742f
C4389 vdd.n1906 gnd 0.583958f
C4390 vdd.n1907 gnd 0.010485f
C4391 vdd.n1908 gnd 0.008439f
C4392 vdd.n1909 gnd 0.010485f
C4393 vdd.n1910 gnd 0.010485f
C4394 vdd.n1911 gnd 0.010485f
C4395 vdd.n1912 gnd 0.008439f
C4396 vdd.n1913 gnd 0.010485f
C4397 vdd.n1914 gnd 0.669677f
C4398 vdd.n1915 gnd 0.010485f
C4399 vdd.n1916 gnd 0.008439f
C4400 vdd.n1917 gnd 0.010485f
C4401 vdd.n1918 gnd 0.010485f
C4402 vdd.n1919 gnd 0.010485f
C4403 vdd.n1920 gnd 0.008439f
C4404 vdd.n1921 gnd 0.010485f
C4405 vdd.n1922 gnd 0.573243f
C4406 vdd.n1923 gnd 0.851829f
C4407 vdd.n1924 gnd 0.010485f
C4408 vdd.n1925 gnd 0.008439f
C4409 vdd.n1926 gnd 0.010485f
C4410 vdd.n1927 gnd 0.010485f
C4411 vdd.n1928 gnd 0.010485f
C4412 vdd.n1929 gnd 0.008439f
C4413 vdd.n1930 gnd 0.010485f
C4414 vdd.n1931 gnd 0.889331f
C4415 vdd.n1932 gnd 0.010485f
C4416 vdd.n1933 gnd 0.008439f
C4417 vdd.n1934 gnd 0.010485f
C4418 vdd.n1935 gnd 0.010485f
C4419 vdd.n1936 gnd 0.010485f
C4420 vdd.n1937 gnd 0.008439f
C4421 vdd.n1938 gnd 0.010485f
C4422 vdd.t166 gnd 0.535742f
C4423 vdd.n1939 gnd 0.744681f
C4424 vdd.n1940 gnd 0.010485f
C4425 vdd.n1941 gnd 0.008439f
C4426 vdd.n1942 gnd 0.010485f
C4427 vdd.n1943 gnd 0.010485f
C4428 vdd.n1944 gnd 0.010485f
C4429 vdd.n1945 gnd 0.008439f
C4430 vdd.n1946 gnd 0.010485f
C4431 vdd.n1947 gnd 0.562529f
C4432 vdd.n1948 gnd 0.010485f
C4433 vdd.n1949 gnd 0.008439f
C4434 vdd.n1950 gnd 0.010485f
C4435 vdd.n1951 gnd 0.010485f
C4436 vdd.n1952 gnd 0.010485f
C4437 vdd.n1953 gnd 0.008439f
C4438 vdd.n1954 gnd 0.010485f
C4439 vdd.n1955 gnd 0.733966f
C4440 vdd.n1956 gnd 0.691107f
C4441 vdd.n1957 gnd 0.010485f
C4442 vdd.n1958 gnd 0.008439f
C4443 vdd.n1959 gnd 0.010485f
C4444 vdd.n1960 gnd 0.010485f
C4445 vdd.n1961 gnd 0.010485f
C4446 vdd.n1962 gnd 0.008439f
C4447 vdd.n1963 gnd 0.010485f
C4448 vdd.n1964 gnd 0.873259f
C4449 vdd.n1965 gnd 0.010485f
C4450 vdd.n1966 gnd 0.008439f
C4451 vdd.n1967 gnd 0.010485f
C4452 vdd.n1968 gnd 0.010485f
C4453 vdd.n1969 gnd 0.025363f
C4454 vdd.n1970 gnd 0.010485f
C4455 vdd.n1971 gnd 0.010485f
C4456 vdd.n1972 gnd 0.008439f
C4457 vdd.n1973 gnd 0.010485f
C4458 vdd.n1974 gnd 0.648247f
C4459 vdd.n1975 gnd 1.07148f
C4460 vdd.n1976 gnd 0.010485f
C4461 vdd.n1977 gnd 0.008439f
C4462 vdd.n1978 gnd 0.010485f
C4463 vdd.n1979 gnd 0.010485f
C4464 vdd.n1980 gnd 0.009017f
C4465 vdd.n1981 gnd 0.008439f
C4466 vdd.n1983 gnd 0.010485f
C4467 vdd.n1985 gnd 0.008439f
C4468 vdd.n1986 gnd 0.010485f
C4469 vdd.n1987 gnd 0.008439f
C4470 vdd.n1989 gnd 0.010485f
C4471 vdd.n1990 gnd 0.008439f
C4472 vdd.n1991 gnd 0.010485f
C4473 vdd.n1992 gnd 0.010485f
C4474 vdd.n1993 gnd 0.010485f
C4475 vdd.n1994 gnd 0.010485f
C4476 vdd.n1995 gnd 0.010485f
C4477 vdd.n1996 gnd 0.008439f
C4478 vdd.n1998 gnd 0.010485f
C4479 vdd.n1999 gnd 0.010485f
C4480 vdd.n2000 gnd 0.010485f
C4481 vdd.n2001 gnd 0.010485f
C4482 vdd.n2002 gnd 0.010485f
C4483 vdd.n2003 gnd 0.008439f
C4484 vdd.n2005 gnd 0.010485f
C4485 vdd.n2006 gnd 0.010485f
C4486 vdd.n2007 gnd 0.010485f
C4487 vdd.n2008 gnd 0.010485f
C4488 vdd.n2009 gnd 0.007046f
C4489 vdd.t80 gnd 0.128989f
C4490 vdd.t79 gnd 0.137854f
C4491 vdd.t78 gnd 0.168458f
C4492 vdd.n2010 gnd 0.215939f
C4493 vdd.n2011 gnd 0.181428f
C4494 vdd.n2013 gnd 0.010485f
C4495 vdd.n2014 gnd 0.010485f
C4496 vdd.n2015 gnd 0.008439f
C4497 vdd.n2016 gnd 0.010485f
C4498 vdd.n2018 gnd 0.010485f
C4499 vdd.n2019 gnd 0.010485f
C4500 vdd.n2020 gnd 0.010485f
C4501 vdd.n2021 gnd 0.010485f
C4502 vdd.n2022 gnd 0.008439f
C4503 vdd.n2024 gnd 0.010485f
C4504 vdd.n2025 gnd 0.010485f
C4505 vdd.n2026 gnd 0.010485f
C4506 vdd.n2027 gnd 0.010485f
C4507 vdd.n2028 gnd 0.010485f
C4508 vdd.n2029 gnd 0.008439f
C4509 vdd.n2031 gnd 0.010485f
C4510 vdd.n2032 gnd 0.010485f
C4511 vdd.n2033 gnd 0.010485f
C4512 vdd.n2034 gnd 0.010485f
C4513 vdd.n2035 gnd 0.010485f
C4514 vdd.n2036 gnd 0.008439f
C4515 vdd.n2038 gnd 0.010485f
C4516 vdd.n2039 gnd 0.010485f
C4517 vdd.n2040 gnd 0.010485f
C4518 vdd.n2041 gnd 0.010485f
C4519 vdd.n2042 gnd 0.010485f
C4520 vdd.n2043 gnd 0.008439f
C4521 vdd.n2045 gnd 0.010485f
C4522 vdd.n2046 gnd 0.010485f
C4523 vdd.n2047 gnd 0.010485f
C4524 vdd.n2048 gnd 0.010485f
C4525 vdd.n2049 gnd 0.008354f
C4526 vdd.t59 gnd 0.128989f
C4527 vdd.t58 gnd 0.137854f
C4528 vdd.t57 gnd 0.168458f
C4529 vdd.n2050 gnd 0.215939f
C4530 vdd.n2051 gnd 0.181428f
C4531 vdd.n2053 gnd 0.010485f
C4532 vdd.n2054 gnd 0.010485f
C4533 vdd.n2055 gnd 0.008439f
C4534 vdd.n2056 gnd 0.010485f
C4535 vdd.n2058 gnd 0.010485f
C4536 vdd.n2059 gnd 0.010485f
C4537 vdd.n2060 gnd 0.010485f
C4538 vdd.n2061 gnd 0.010485f
C4539 vdd.n2062 gnd 0.008439f
C4540 vdd.n2064 gnd 0.010485f
C4541 vdd.n2065 gnd 0.010485f
C4542 vdd.n2066 gnd 0.010485f
C4543 vdd.n2067 gnd 0.010485f
C4544 vdd.n2068 gnd 0.010485f
C4545 vdd.n2069 gnd 0.008439f
C4546 vdd.n2071 gnd 0.010485f
C4547 vdd.n2072 gnd 0.010485f
C4548 vdd.n2073 gnd 0.010485f
C4549 vdd.n2074 gnd 0.010485f
C4550 vdd.n2075 gnd 0.010485f
C4551 vdd.n2076 gnd 0.010485f
C4552 vdd.n2077 gnd 0.008439f
C4553 vdd.n2079 gnd 0.010485f
C4554 vdd.n2081 gnd 0.010485f
C4555 vdd.n2082 gnd 0.008439f
C4556 vdd.n2083 gnd 0.008439f
C4557 vdd.n2084 gnd 0.010485f
C4558 vdd.n2086 gnd 0.010485f
C4559 vdd.n2087 gnd 0.008439f
C4560 vdd.n2088 gnd 0.008439f
C4561 vdd.n2089 gnd 0.010485f
C4562 vdd.n2091 gnd 0.010485f
C4563 vdd.n2092 gnd 0.010485f
C4564 vdd.n2093 gnd 0.008439f
C4565 vdd.n2094 gnd 0.008439f
C4566 vdd.n2095 gnd 0.008439f
C4567 vdd.n2096 gnd 0.010485f
C4568 vdd.n2098 gnd 0.010485f
C4569 vdd.n2099 gnd 0.010485f
C4570 vdd.n2100 gnd 0.008439f
C4571 vdd.n2101 gnd 0.008439f
C4572 vdd.n2102 gnd 0.008439f
C4573 vdd.n2103 gnd 0.010485f
C4574 vdd.n2105 gnd 0.010485f
C4575 vdd.n2106 gnd 0.010485f
C4576 vdd.n2107 gnd 0.008439f
C4577 vdd.n2108 gnd 0.008439f
C4578 vdd.n2109 gnd 0.008439f
C4579 vdd.n2110 gnd 0.010485f
C4580 vdd.n2112 gnd 0.010485f
C4581 vdd.n2113 gnd 0.010485f
C4582 vdd.n2114 gnd 0.008439f
C4583 vdd.n2115 gnd 0.010485f
C4584 vdd.n2116 gnd 0.010485f
C4585 vdd.n2117 gnd 0.010485f
C4586 vdd.n2118 gnd 0.017215f
C4587 vdd.n2119 gnd 0.005738f
C4588 vdd.n2120 gnd 0.008439f
C4589 vdd.n2121 gnd 0.010485f
C4590 vdd.n2123 gnd 0.010485f
C4591 vdd.n2124 gnd 0.010485f
C4592 vdd.n2125 gnd 0.008439f
C4593 vdd.n2126 gnd 0.008439f
C4594 vdd.n2127 gnd 0.008439f
C4595 vdd.n2128 gnd 0.010485f
C4596 vdd.n2130 gnd 0.010485f
C4597 vdd.n2131 gnd 0.010485f
C4598 vdd.n2132 gnd 0.008439f
C4599 vdd.n2133 gnd 0.008439f
C4600 vdd.n2134 gnd 0.008439f
C4601 vdd.n2135 gnd 0.010485f
C4602 vdd.n2137 gnd 0.010485f
C4603 vdd.n2138 gnd 0.010485f
C4604 vdd.n2139 gnd 0.008439f
C4605 vdd.n2140 gnd 0.008439f
C4606 vdd.n2141 gnd 0.008439f
C4607 vdd.n2142 gnd 0.010485f
C4608 vdd.n2144 gnd 0.010485f
C4609 vdd.n2145 gnd 0.010485f
C4610 vdd.n2146 gnd 0.008439f
C4611 vdd.n2147 gnd 0.008439f
C4612 vdd.n2148 gnd 0.008439f
C4613 vdd.n2149 gnd 0.010485f
C4614 vdd.n2151 gnd 0.010485f
C4615 vdd.n2152 gnd 0.010485f
C4616 vdd.n2153 gnd 0.008439f
C4617 vdd.n2154 gnd 0.010485f
C4618 vdd.n2155 gnd 0.010485f
C4619 vdd.n2156 gnd 0.010485f
C4620 vdd.n2157 gnd 0.017215f
C4621 vdd.n2158 gnd 0.007046f
C4622 vdd.n2159 gnd 0.008439f
C4623 vdd.n2160 gnd 0.010485f
C4624 vdd.n2162 gnd 0.010485f
C4625 vdd.n2163 gnd 0.010485f
C4626 vdd.n2164 gnd 0.008439f
C4627 vdd.n2165 gnd 0.008439f
C4628 vdd.n2166 gnd 0.008439f
C4629 vdd.n2167 gnd 0.010485f
C4630 vdd.n2169 gnd 0.010485f
C4631 vdd.n2170 gnd 0.010485f
C4632 vdd.n2171 gnd 0.008439f
C4633 vdd.n2172 gnd 0.008439f
C4634 vdd.n2173 gnd 0.008439f
C4635 vdd.n2174 gnd 0.010485f
C4636 vdd.n2176 gnd 0.010485f
C4637 vdd.n2177 gnd 0.010485f
C4638 vdd.n2179 gnd 0.010485f
C4639 vdd.n2180 gnd 0.008439f
C4640 vdd.n2181 gnd 0.00671f
C4641 vdd.n2182 gnd 0.95377f
C4642 vdd.n2184 gnd 0.008439f
C4643 vdd.n2185 gnd 0.008439f
C4644 vdd.n2186 gnd 0.010485f
C4645 vdd.n2188 gnd 0.010485f
C4646 vdd.n2189 gnd 0.010485f
C4647 vdd.n2190 gnd 0.008439f
C4648 vdd.n2191 gnd 0.007004f
C4649 vdd.n2192 gnd 0.025907f
C4650 vdd.n2193 gnd 0.025363f
C4651 vdd.n2194 gnd 0.007004f
C4652 vdd.n2195 gnd 0.025363f
C4653 vdd.n2196 gnd 1.47329f
C4654 vdd.n2197 gnd 0.025363f
C4655 vdd.n2198 gnd 0.025907f
C4656 vdd.n2199 gnd 0.004008f
C4657 vdd.t50 gnd 0.128989f
C4658 vdd.t49 gnd 0.137854f
C4659 vdd.t47 gnd 0.168458f
C4660 vdd.n2200 gnd 0.215939f
C4661 vdd.n2201 gnd 0.181428f
C4662 vdd.n2202 gnd 0.012996f
C4663 vdd.n2203 gnd 0.00443f
C4664 vdd.n2204 gnd 0.009017f
C4665 vdd.n2205 gnd 0.95377f
C4666 vdd.n2206 gnd 0.037513f
C4667 vdd.n2207 gnd 0.00713f
C4668 vdd.n2208 gnd 0.00713f
C4669 vdd.n2209 gnd 0.00713f
C4670 vdd.n2210 gnd 0.00713f
C4671 vdd.n2211 gnd 0.00713f
C4672 vdd.n2212 gnd 0.00713f
C4673 vdd.n2213 gnd 0.00713f
C4674 vdd.n2214 gnd 0.00713f
C4675 vdd.n2216 gnd 0.00713f
C4676 vdd.n2218 gnd 0.00713f
C4677 vdd.n2219 gnd 0.00713f
C4678 vdd.n2220 gnd 0.00713f
C4679 vdd.n2221 gnd 0.00713f
C4680 vdd.n2222 gnd 0.00713f
C4681 vdd.n2224 gnd 0.00713f
C4682 vdd.n2226 gnd 0.00713f
C4683 vdd.n2227 gnd 0.00713f
C4684 vdd.n2228 gnd 0.00713f
C4685 vdd.n2229 gnd 0.00713f
C4686 vdd.n2230 gnd 0.00713f
C4687 vdd.n2232 gnd 0.00713f
C4688 vdd.n2234 gnd 0.00713f
C4689 vdd.n2235 gnd 0.00713f
C4690 vdd.n2236 gnd 0.00713f
C4691 vdd.n2237 gnd 0.00713f
C4692 vdd.n2238 gnd 0.00713f
C4693 vdd.n2240 gnd 0.00713f
C4694 vdd.n2242 gnd 0.00713f
C4695 vdd.n2243 gnd 0.00713f
C4696 vdd.n2244 gnd 0.00713f
C4697 vdd.n2245 gnd 0.00713f
C4698 vdd.n2246 gnd 0.00713f
C4699 vdd.n2248 gnd 0.00713f
C4700 vdd.n2250 gnd 0.00713f
C4701 vdd.n2251 gnd 0.00713f
C4702 vdd.n2252 gnd 0.00713f
C4703 vdd.n2253 gnd 0.00713f
C4704 vdd.n2254 gnd 0.00713f
C4705 vdd.n2256 gnd 0.00713f
C4706 vdd.n2258 gnd 0.00713f
C4707 vdd.n2259 gnd 0.00713f
C4708 vdd.n2260 gnd 0.00713f
C4709 vdd.n2261 gnd 0.00713f
C4710 vdd.n2262 gnd 0.00713f
C4711 vdd.n2264 gnd 0.00713f
C4712 vdd.n2266 gnd 0.00713f
C4713 vdd.n2267 gnd 0.00713f
C4714 vdd.n2268 gnd 0.00713f
C4715 vdd.n2269 gnd 0.00713f
C4716 vdd.n2270 gnd 0.00713f
C4717 vdd.n2272 gnd 0.00713f
C4718 vdd.n2274 gnd 0.00713f
C4719 vdd.n2275 gnd 0.00713f
C4720 vdd.n2276 gnd 0.00519f
C4721 vdd.n2277 gnd 0.010189f
C4722 vdd.n2278 gnd 0.005504f
C4723 vdd.n2279 gnd 0.00713f
C4724 vdd.n2281 gnd 0.00713f
C4725 vdd.n2282 gnd 0.016433f
C4726 vdd.n2283 gnd 0.016433f
C4727 vdd.n2284 gnd 0.015441f
C4728 vdd.n2285 gnd 0.00713f
C4729 vdd.n2286 gnd 0.00713f
C4730 vdd.n2287 gnd 0.00713f
C4731 vdd.n2288 gnd 0.00713f
C4732 vdd.n2289 gnd 0.00713f
C4733 vdd.n2290 gnd 0.00713f
C4734 vdd.n2291 gnd 0.00713f
C4735 vdd.n2292 gnd 0.00713f
C4736 vdd.n2293 gnd 0.00713f
C4737 vdd.n2294 gnd 0.00713f
C4738 vdd.n2295 gnd 0.00713f
C4739 vdd.n2296 gnd 0.00713f
C4740 vdd.n2297 gnd 0.00713f
C4741 vdd.n2298 gnd 0.00713f
C4742 vdd.n2299 gnd 0.00713f
C4743 vdd.n2300 gnd 0.00713f
C4744 vdd.n2301 gnd 0.00713f
C4745 vdd.n2302 gnd 0.00713f
C4746 vdd.n2303 gnd 0.00713f
C4747 vdd.n2304 gnd 0.00713f
C4748 vdd.n2305 gnd 0.00713f
C4749 vdd.n2306 gnd 0.00713f
C4750 vdd.n2307 gnd 0.00713f
C4751 vdd.n2308 gnd 0.00713f
C4752 vdd.n2309 gnd 0.00713f
C4753 vdd.n2310 gnd 0.00713f
C4754 vdd.n2311 gnd 0.00713f
C4755 vdd.n2312 gnd 0.00713f
C4756 vdd.n2313 gnd 0.00713f
C4757 vdd.n2314 gnd 0.00713f
C4758 vdd.n2315 gnd 0.00713f
C4759 vdd.n2316 gnd 0.00713f
C4760 vdd.n2317 gnd 0.00713f
C4761 vdd.n2318 gnd 0.00713f
C4762 vdd.n2319 gnd 0.00713f
C4763 vdd.n2320 gnd 0.00713f
C4764 vdd.n2321 gnd 0.00713f
C4765 vdd.n2322 gnd 0.00713f
C4766 vdd.n2323 gnd 0.00713f
C4767 vdd.n2324 gnd 0.00713f
C4768 vdd.n2325 gnd 0.00713f
C4769 vdd.n2326 gnd 0.00713f
C4770 vdd.n2327 gnd 0.00713f
C4771 vdd.n2328 gnd 0.00713f
C4772 vdd.n2329 gnd 0.00713f
C4773 vdd.n2330 gnd 0.00713f
C4774 vdd.n2331 gnd 0.00713f
C4775 vdd.n2332 gnd 0.00713f
C4776 vdd.n2333 gnd 0.00713f
C4777 vdd.n2334 gnd 0.433951f
C4778 vdd.n2335 gnd 0.00713f
C4779 vdd.n2336 gnd 0.00713f
C4780 vdd.n2337 gnd 0.00713f
C4781 vdd.n2338 gnd 0.00713f
C4782 vdd.n2339 gnd 0.00713f
C4783 vdd.n2340 gnd 0.00713f
C4784 vdd.n2341 gnd 0.00713f
C4785 vdd.n2342 gnd 0.00713f
C4786 vdd.n2343 gnd 0.00713f
C4787 vdd.n2344 gnd 0.00713f
C4788 vdd.n2345 gnd 0.00713f
C4789 vdd.n2346 gnd 0.658962f
C4790 vdd.n2347 gnd 0.00713f
C4791 vdd.n2348 gnd 0.00713f
C4792 vdd.n2349 gnd 0.00713f
C4793 vdd.n2350 gnd 0.00713f
C4794 vdd.n2351 gnd 0.00713f
C4795 vdd.n2352 gnd 0.00713f
C4796 vdd.n2353 gnd 0.00713f
C4797 vdd.n2354 gnd 0.00713f
C4798 vdd.n2355 gnd 0.00713f
C4799 vdd.n2356 gnd 0.00713f
C4800 vdd.n2357 gnd 0.00713f
C4801 vdd.n2358 gnd 0.230369f
C4802 vdd.n2359 gnd 0.00713f
C4803 vdd.n2360 gnd 0.00713f
C4804 vdd.n2361 gnd 0.00713f
C4805 vdd.n2362 gnd 0.00713f
C4806 vdd.n2363 gnd 0.00713f
C4807 vdd.n2364 gnd 0.00713f
C4808 vdd.n2365 gnd 0.00713f
C4809 vdd.n2366 gnd 0.00713f
C4810 vdd.n2367 gnd 0.00713f
C4811 vdd.n2368 gnd 0.00713f
C4812 vdd.n2369 gnd 0.00713f
C4813 vdd.n2370 gnd 0.00713f
C4814 vdd.n2371 gnd 0.00713f
C4815 vdd.n2372 gnd 0.00713f
C4816 vdd.n2373 gnd 0.00713f
C4817 vdd.n2374 gnd 0.00713f
C4818 vdd.n2375 gnd 0.00713f
C4819 vdd.n2376 gnd 0.00713f
C4820 vdd.n2377 gnd 0.00713f
C4821 vdd.n2378 gnd 0.00713f
C4822 vdd.n2379 gnd 0.00713f
C4823 vdd.n2380 gnd 0.00713f
C4824 vdd.n2381 gnd 0.00713f
C4825 vdd.n2382 gnd 0.00713f
C4826 vdd.n2383 gnd 0.00713f
C4827 vdd.n2384 gnd 0.00713f
C4828 vdd.n2385 gnd 0.00713f
C4829 vdd.n2386 gnd 0.00713f
C4830 vdd.n2387 gnd 0.00713f
C4831 vdd.n2388 gnd 0.00713f
C4832 vdd.n2389 gnd 0.00713f
C4833 vdd.n2390 gnd 0.00713f
C4834 vdd.n2391 gnd 0.00713f
C4835 vdd.n2392 gnd 0.00713f
C4836 vdd.n2393 gnd 0.00713f
C4837 vdd.n2394 gnd 0.015441f
C4838 vdd.n2395 gnd 0.016433f
C4839 vdd.n2396 gnd 0.016433f
C4840 vdd.n2398 gnd 0.00713f
C4841 vdd.n2400 gnd 0.00713f
C4842 vdd.n2401 gnd 0.005504f
C4843 vdd.n2402 gnd 0.010189f
C4844 vdd.n2403 gnd 0.00519f
C4845 vdd.n2404 gnd 0.00713f
C4846 vdd.n2405 gnd 0.00713f
C4847 vdd.n2407 gnd 0.00713f
C4848 vdd.n2409 gnd 0.00713f
C4849 vdd.n2410 gnd 0.00713f
C4850 vdd.n2411 gnd 0.00713f
C4851 vdd.n2412 gnd 0.00713f
C4852 vdd.n2413 gnd 0.00713f
C4853 vdd.n2415 gnd 0.00713f
C4854 vdd.n2417 gnd 0.00713f
C4855 vdd.n2418 gnd 0.00713f
C4856 vdd.n2419 gnd 0.00713f
C4857 vdd.n2420 gnd 0.00713f
C4858 vdd.n2421 gnd 0.00713f
C4859 vdd.n2423 gnd 0.00713f
C4860 vdd.n2425 gnd 0.00713f
C4861 vdd.n2426 gnd 0.00713f
C4862 vdd.n2427 gnd 0.00713f
C4863 vdd.n2428 gnd 0.00713f
C4864 vdd.n2429 gnd 0.00713f
C4865 vdd.n2431 gnd 0.00713f
C4866 vdd.n2433 gnd 0.00713f
C4867 vdd.n2434 gnd 0.00713f
C4868 vdd.n2435 gnd 0.00713f
C4869 vdd.n2436 gnd 0.00713f
C4870 vdd.n2437 gnd 0.00713f
C4871 vdd.n2439 gnd 0.00713f
C4872 vdd.n2441 gnd 0.00713f
C4873 vdd.n2442 gnd 0.00713f
C4874 vdd.n2443 gnd 0.00713f
C4875 vdd.n2444 gnd 0.00713f
C4876 vdd.n2445 gnd 0.00713f
C4877 vdd.n2447 gnd 0.00713f
C4878 vdd.n2449 gnd 0.00713f
C4879 vdd.n2450 gnd 0.00713f
C4880 vdd.n2451 gnd 0.00713f
C4881 vdd.n2452 gnd 0.00713f
C4882 vdd.n2453 gnd 0.00713f
C4883 vdd.n2455 gnd 0.00713f
C4884 vdd.n2456 gnd 0.00713f
C4885 vdd.n2457 gnd 0.00713f
C4886 vdd.n2458 gnd 0.00713f
C4887 vdd.n2459 gnd 0.00713f
C4888 vdd.n2460 gnd 0.00713f
C4889 vdd.n2462 gnd 0.00713f
C4890 vdd.n2463 gnd 0.00713f
C4891 vdd.n2464 gnd 0.016433f
C4892 vdd.n2465 gnd 0.015441f
C4893 vdd.n2466 gnd 0.015441f
C4894 vdd.n2467 gnd 1.00719f
C4895 vdd.n2468 gnd 0.015441f
C4896 vdd.n2469 gnd 0.015441f
C4897 vdd.n2470 gnd 0.00713f
C4898 vdd.n2471 gnd 0.00713f
C4899 vdd.n2472 gnd 0.00713f
C4900 vdd.n2473 gnd 0.49824f
C4901 vdd.n2474 gnd 0.00713f
C4902 vdd.n2475 gnd 0.00713f
C4903 vdd.n2476 gnd 0.00713f
C4904 vdd.n2477 gnd 0.00713f
C4905 vdd.n2478 gnd 0.00713f
C4906 vdd.n2479 gnd 0.728608f
C4907 vdd.n2480 gnd 0.00713f
C4908 vdd.n2481 gnd 0.00713f
C4909 vdd.n2482 gnd 0.00713f
C4910 vdd.n2483 gnd 0.00713f
C4911 vdd.n2484 gnd 0.00713f
C4912 vdd.n2485 gnd 0.728608f
C4913 vdd.n2486 gnd 0.00713f
C4914 vdd.n2487 gnd 0.00713f
C4915 vdd.n2488 gnd 0.00713f
C4916 vdd.n2489 gnd 0.00713f
C4917 vdd.n2490 gnd 0.00713f
C4918 vdd.n2491 gnd 0.369662f
C4919 vdd.n2492 gnd 0.00713f
C4920 vdd.n2493 gnd 0.00713f
C4921 vdd.n2494 gnd 0.00713f
C4922 vdd.n2495 gnd 0.00713f
C4923 vdd.n2496 gnd 0.00713f
C4924 vdd.n2497 gnd 0.530384f
C4925 vdd.n2498 gnd 0.00713f
C4926 vdd.n2499 gnd 0.00713f
C4927 vdd.n2500 gnd 0.00713f
C4928 vdd.n2501 gnd 0.00713f
C4929 vdd.n2502 gnd 0.00713f
C4930 vdd.n2503 gnd 0.691107f
C4931 vdd.n2504 gnd 0.00713f
C4932 vdd.n2505 gnd 0.00713f
C4933 vdd.n2506 gnd 0.00713f
C4934 vdd.n2507 gnd 0.00713f
C4935 vdd.n2508 gnd 0.00713f
C4936 vdd.n2509 gnd 0.728608f
C4937 vdd.n2510 gnd 0.00713f
C4938 vdd.n2511 gnd 0.00713f
C4939 vdd.n2512 gnd 0.00713f
C4940 vdd.n2513 gnd 0.00713f
C4941 vdd.n2514 gnd 0.00713f
C4942 vdd.n2515 gnd 0.605388f
C4943 vdd.n2516 gnd 0.00713f
C4944 vdd.n2517 gnd 0.00713f
C4945 vdd.n2518 gnd 0.005871f
C4946 vdd.n2519 gnd 0.020653f
C4947 vdd.n2520 gnd 0.004823f
C4948 vdd.n2521 gnd 0.00713f
C4949 vdd.n2522 gnd 0.444665f
C4950 vdd.n2523 gnd 0.00713f
C4951 vdd.n2524 gnd 0.00713f
C4952 vdd.n2525 gnd 0.00713f
C4953 vdd.n2526 gnd 0.00713f
C4954 vdd.n2527 gnd 0.00713f
C4955 vdd.n2528 gnd 0.444665f
C4956 vdd.n2529 gnd 0.00713f
C4957 vdd.n2530 gnd 0.00713f
C4958 vdd.n2531 gnd 0.00713f
C4959 vdd.n2532 gnd 0.00713f
C4960 vdd.n2533 gnd 0.00713f
C4961 vdd.n2534 gnd 0.605388f
C4962 vdd.n2535 gnd 0.00713f
C4963 vdd.n2536 gnd 0.00713f
C4964 vdd.n2537 gnd 0.00713f
C4965 vdd.n2538 gnd 0.00713f
C4966 vdd.n2539 gnd 0.00713f
C4967 vdd.n2540 gnd 0.62146f
C4968 vdd.n2541 gnd 0.00713f
C4969 vdd.n2542 gnd 0.00713f
C4970 vdd.n2543 gnd 0.00713f
C4971 vdd.n2544 gnd 0.00713f
C4972 vdd.n2545 gnd 0.00713f
C4973 vdd.n2546 gnd 0.460738f
C4974 vdd.n2547 gnd 0.00713f
C4975 vdd.n2548 gnd 0.00713f
C4976 vdd.n2549 gnd 0.00713f
C4977 vdd.n2550 gnd 0.00713f
C4978 vdd.n2551 gnd 0.00713f
C4979 vdd.n2552 gnd 0.230369f
C4980 vdd.n2553 gnd 0.00713f
C4981 vdd.n2554 gnd 0.00713f
C4982 vdd.n2555 gnd 0.00713f
C4983 vdd.n2556 gnd 0.00713f
C4984 vdd.n2557 gnd 0.00713f
C4985 vdd.n2558 gnd 0.230369f
C4986 vdd.n2559 gnd 0.00713f
C4987 vdd.n2560 gnd 0.00713f
C4988 vdd.n2561 gnd 0.00713f
C4989 vdd.n2562 gnd 0.00713f
C4990 vdd.n2563 gnd 0.00713f
C4991 vdd.n2564 gnd 0.728608f
C4992 vdd.n2565 gnd 0.00713f
C4993 vdd.n2566 gnd 0.00713f
C4994 vdd.n2567 gnd 0.00713f
C4995 vdd.n2568 gnd 0.00713f
C4996 vdd.n2569 gnd 0.00713f
C4997 vdd.n2570 gnd 0.00713f
C4998 vdd.n2571 gnd 0.00713f
C4999 vdd.n2572 gnd 0.525027f
C5000 vdd.n2573 gnd 0.00713f
C5001 vdd.n2574 gnd 0.00713f
C5002 vdd.n2575 gnd 0.00713f
C5003 vdd.n2576 gnd 0.00713f
C5004 vdd.n2577 gnd 0.00713f
C5005 vdd.n2578 gnd 0.00713f
C5006 vdd.n2579 gnd 0.45538f
C5007 vdd.n2580 gnd 0.00713f
C5008 vdd.n2581 gnd 0.00713f
C5009 vdd.n2582 gnd 0.00713f
C5010 vdd.n2583 gnd 0.016345f
C5011 vdd.n2584 gnd 0.015529f
C5012 vdd.n2585 gnd 0.00713f
C5013 vdd.n2586 gnd 0.00713f
C5014 vdd.n2587 gnd 0.005504f
C5015 vdd.n2588 gnd 0.00713f
C5016 vdd.n2589 gnd 0.00713f
C5017 vdd.n2590 gnd 0.00519f
C5018 vdd.n2591 gnd 0.00713f
C5019 vdd.n2592 gnd 0.00713f
C5020 vdd.n2593 gnd 0.00713f
C5021 vdd.n2594 gnd 0.00713f
C5022 vdd.n2595 gnd 0.00713f
C5023 vdd.n2596 gnd 0.00713f
C5024 vdd.n2597 gnd 0.00713f
C5025 vdd.n2598 gnd 0.00713f
C5026 vdd.n2599 gnd 0.00713f
C5027 vdd.n2600 gnd 0.00713f
C5028 vdd.n2601 gnd 0.00713f
C5029 vdd.n2602 gnd 0.00713f
C5030 vdd.n2603 gnd 0.00713f
C5031 vdd.n2604 gnd 0.00713f
C5032 vdd.n2605 gnd 0.00713f
C5033 vdd.n2606 gnd 0.00713f
C5034 vdd.n2607 gnd 0.00713f
C5035 vdd.n2608 gnd 0.00713f
C5036 vdd.n2609 gnd 0.00713f
C5037 vdd.n2610 gnd 0.00713f
C5038 vdd.n2611 gnd 0.00713f
C5039 vdd.n2612 gnd 0.00713f
C5040 vdd.n2613 gnd 0.00713f
C5041 vdd.n2614 gnd 0.00713f
C5042 vdd.n2615 gnd 0.00713f
C5043 vdd.n2616 gnd 0.00713f
C5044 vdd.n2617 gnd 0.00713f
C5045 vdd.n2618 gnd 0.00713f
C5046 vdd.n2619 gnd 0.00713f
C5047 vdd.n2620 gnd 0.00713f
C5048 vdd.n2621 gnd 0.00713f
C5049 vdd.n2622 gnd 0.00713f
C5050 vdd.n2623 gnd 0.00713f
C5051 vdd.n2624 gnd 0.00713f
C5052 vdd.n2625 gnd 0.00713f
C5053 vdd.n2626 gnd 0.00713f
C5054 vdd.n2627 gnd 0.00713f
C5055 vdd.n2628 gnd 0.00713f
C5056 vdd.n2629 gnd 0.00713f
C5057 vdd.n2630 gnd 0.00713f
C5058 vdd.n2631 gnd 0.00713f
C5059 vdd.n2632 gnd 0.00713f
C5060 vdd.n2633 gnd 0.00713f
C5061 vdd.n2634 gnd 0.00713f
C5062 vdd.n2635 gnd 0.00713f
C5063 vdd.n2636 gnd 0.00713f
C5064 vdd.n2637 gnd 0.00713f
C5065 vdd.n2638 gnd 0.00713f
C5066 vdd.n2639 gnd 0.00713f
C5067 vdd.n2640 gnd 0.00713f
C5068 vdd.n2641 gnd 0.00713f
C5069 vdd.n2642 gnd 0.00713f
C5070 vdd.n2643 gnd 0.00713f
C5071 vdd.n2644 gnd 0.00713f
C5072 vdd.n2645 gnd 0.00713f
C5073 vdd.n2646 gnd 0.00713f
C5074 vdd.n2647 gnd 0.00713f
C5075 vdd.n2648 gnd 0.00713f
C5076 vdd.n2649 gnd 0.00713f
C5077 vdd.n2650 gnd 0.00713f
C5078 vdd.n2651 gnd 0.016433f
C5079 vdd.n2652 gnd 0.015441f
C5080 vdd.n2653 gnd 0.015441f
C5081 vdd.n2654 gnd 0.846472f
C5082 vdd.n2655 gnd 0.015441f
C5083 vdd.n2656 gnd 0.016433f
C5084 vdd.n2657 gnd 0.015529f
C5085 vdd.n2658 gnd 0.00713f
C5086 vdd.n2659 gnd 0.00713f
C5087 vdd.n2660 gnd 0.00713f
C5088 vdd.n2661 gnd 0.005504f
C5089 vdd.n2662 gnd 0.010189f
C5090 vdd.n2663 gnd 0.00519f
C5091 vdd.n2664 gnd 0.00713f
C5092 vdd.n2665 gnd 0.00713f
C5093 vdd.n2666 gnd 0.00713f
C5094 vdd.n2667 gnd 0.00713f
C5095 vdd.n2668 gnd 0.00713f
C5096 vdd.n2669 gnd 0.00713f
C5097 vdd.n2670 gnd 0.00713f
C5098 vdd.n2671 gnd 0.00713f
C5099 vdd.n2672 gnd 0.00713f
C5100 vdd.n2673 gnd 0.00713f
C5101 vdd.n2674 gnd 0.00713f
C5102 vdd.n2675 gnd 0.00713f
C5103 vdd.n2676 gnd 0.00713f
C5104 vdd.n2677 gnd 0.00713f
C5105 vdd.n2678 gnd 0.00713f
C5106 vdd.n2679 gnd 0.00713f
C5107 vdd.n2680 gnd 0.00713f
C5108 vdd.n2681 gnd 0.00713f
C5109 vdd.n2682 gnd 0.00713f
C5110 vdd.n2683 gnd 0.00713f
C5111 vdd.n2684 gnd 0.00713f
C5112 vdd.n2685 gnd 0.00713f
C5113 vdd.n2686 gnd 0.00713f
C5114 vdd.n2687 gnd 0.00713f
C5115 vdd.n2688 gnd 0.00713f
C5116 vdd.n2689 gnd 0.00713f
C5117 vdd.n2690 gnd 0.00713f
C5118 vdd.n2691 gnd 0.00713f
C5119 vdd.n2692 gnd 0.00713f
C5120 vdd.n2693 gnd 0.00713f
C5121 vdd.n2694 gnd 0.00713f
C5122 vdd.n2695 gnd 0.00713f
C5123 vdd.n2696 gnd 0.00713f
C5124 vdd.n2697 gnd 0.00713f
C5125 vdd.n2698 gnd 0.00713f
C5126 vdd.n2699 gnd 0.00713f
C5127 vdd.n2700 gnd 0.00713f
C5128 vdd.n2701 gnd 0.00713f
C5129 vdd.n2702 gnd 0.00713f
C5130 vdd.n2703 gnd 0.00713f
C5131 vdd.n2704 gnd 0.00713f
C5132 vdd.n2705 gnd 0.00713f
C5133 vdd.n2706 gnd 0.00713f
C5134 vdd.n2707 gnd 0.00713f
C5135 vdd.n2708 gnd 0.00713f
C5136 vdd.n2709 gnd 0.00713f
C5137 vdd.n2710 gnd 0.00713f
C5138 vdd.n2711 gnd 0.00713f
C5139 vdd.n2712 gnd 0.00713f
C5140 vdd.n2713 gnd 0.00713f
C5141 vdd.n2714 gnd 0.00713f
C5142 vdd.n2715 gnd 0.00713f
C5143 vdd.n2716 gnd 0.00713f
C5144 vdd.n2717 gnd 0.00713f
C5145 vdd.n2718 gnd 0.00713f
C5146 vdd.n2719 gnd 0.00713f
C5147 vdd.n2720 gnd 0.00713f
C5148 vdd.n2721 gnd 0.00713f
C5149 vdd.n2722 gnd 0.00713f
C5150 vdd.n2723 gnd 0.00713f
C5151 vdd.n2724 gnd 0.016433f
C5152 vdd.n2725 gnd 0.016433f
C5153 vdd.n2726 gnd 0.889331f
C5154 vdd.t128 gnd 3.16088f
C5155 vdd.t125 gnd 3.16088f
C5156 vdd.n2760 gnd 0.00713f
C5157 vdd.t86 gnd 0.288105f
C5158 vdd.t87 gnd 0.294911f
C5159 vdd.t85 gnd 0.188086f
C5160 vdd.n2761 gnd 0.10165f
C5161 vdd.n2762 gnd 0.057659f
C5162 vdd.n2763 gnd 0.010189f
C5163 vdd.n2764 gnd 0.00713f
C5164 vdd.n2765 gnd 0.00713f
C5165 vdd.n2766 gnd 0.00713f
C5166 vdd.n2767 gnd 0.00713f
C5167 vdd.n2768 gnd 0.00713f
C5168 vdd.n2769 gnd 0.00713f
C5169 vdd.n2770 gnd 0.00713f
C5170 vdd.n2771 gnd 0.00713f
C5171 vdd.n2772 gnd 0.00713f
C5172 vdd.n2773 gnd 0.00713f
C5173 vdd.n2774 gnd 0.00713f
C5174 vdd.n2775 gnd 0.00713f
C5175 vdd.n2776 gnd 0.00713f
C5176 vdd.n2777 gnd 0.00713f
C5177 vdd.n2778 gnd 0.00713f
C5178 vdd.n2779 gnd 0.00713f
C5179 vdd.n2780 gnd 0.00713f
C5180 vdd.n2781 gnd 0.00713f
C5181 vdd.n2782 gnd 0.00713f
C5182 vdd.n2783 gnd 0.00713f
C5183 vdd.n2784 gnd 0.00713f
C5184 vdd.n2785 gnd 0.00713f
C5185 vdd.n2786 gnd 0.00713f
C5186 vdd.n2787 gnd 0.00713f
C5187 vdd.n2788 gnd 0.00713f
C5188 vdd.n2789 gnd 0.00713f
C5189 vdd.n2790 gnd 0.00713f
C5190 vdd.n2791 gnd 0.00713f
C5191 vdd.n2792 gnd 0.00713f
C5192 vdd.n2793 gnd 0.00713f
C5193 vdd.n2794 gnd 0.00713f
C5194 vdd.n2795 gnd 0.00713f
C5195 vdd.n2796 gnd 0.00713f
C5196 vdd.n2797 gnd 0.00713f
C5197 vdd.n2798 gnd 0.00713f
C5198 vdd.n2799 gnd 0.00713f
C5199 vdd.n2800 gnd 0.00713f
C5200 vdd.n2801 gnd 0.00713f
C5201 vdd.n2802 gnd 0.00713f
C5202 vdd.n2803 gnd 0.00713f
C5203 vdd.n2804 gnd 0.00713f
C5204 vdd.n2805 gnd 0.00713f
C5205 vdd.n2806 gnd 0.00713f
C5206 vdd.n2807 gnd 0.00713f
C5207 vdd.n2808 gnd 0.00713f
C5208 vdd.n2809 gnd 0.00713f
C5209 vdd.n2810 gnd 0.00713f
C5210 vdd.n2811 gnd 0.00713f
C5211 vdd.n2812 gnd 0.00713f
C5212 vdd.n2813 gnd 0.00713f
C5213 vdd.n2814 gnd 0.00713f
C5214 vdd.n2815 gnd 0.00713f
C5215 vdd.n2816 gnd 0.00713f
C5216 vdd.n2817 gnd 0.00713f
C5217 vdd.n2818 gnd 0.00713f
C5218 vdd.n2819 gnd 0.00713f
C5219 vdd.n2820 gnd 0.00713f
C5220 vdd.n2821 gnd 0.00713f
C5221 vdd.n2822 gnd 0.00713f
C5222 vdd.n2823 gnd 0.00713f
C5223 vdd.n2824 gnd 0.00519f
C5224 vdd.n2825 gnd 0.00713f
C5225 vdd.n2826 gnd 0.00713f
C5226 vdd.n2827 gnd 0.005504f
C5227 vdd.n2828 gnd 0.00713f
C5228 vdd.n2829 gnd 0.00713f
C5229 vdd.t73 gnd 0.288105f
C5230 vdd.t74 gnd 0.294911f
C5231 vdd.t71 gnd 0.188086f
C5232 vdd.n2830 gnd 0.10165f
C5233 vdd.n2831 gnd 0.057659f
C5234 vdd.n2832 gnd 0.00713f
C5235 vdd.n2833 gnd 0.00713f
C5236 vdd.n2834 gnd 0.00713f
C5237 vdd.n2835 gnd 0.00713f
C5238 vdd.n2836 gnd 0.00713f
C5239 vdd.n2837 gnd 0.00713f
C5240 vdd.n2838 gnd 0.00713f
C5241 vdd.n2839 gnd 0.00713f
C5242 vdd.n2840 gnd 0.00713f
C5243 vdd.n2841 gnd 0.00713f
C5244 vdd.n2842 gnd 0.00713f
C5245 vdd.n2843 gnd 0.00713f
C5246 vdd.n2844 gnd 0.00713f
C5247 vdd.n2845 gnd 0.00713f
C5248 vdd.n2846 gnd 0.00713f
C5249 vdd.n2847 gnd 0.00713f
C5250 vdd.n2848 gnd 0.00713f
C5251 vdd.n2849 gnd 0.00713f
C5252 vdd.n2850 gnd 0.00713f
C5253 vdd.n2851 gnd 0.00713f
C5254 vdd.n2852 gnd 0.00713f
C5255 vdd.n2853 gnd 0.00713f
C5256 vdd.n2854 gnd 0.00713f
C5257 vdd.n2855 gnd 0.00713f
C5258 vdd.n2856 gnd 0.00713f
C5259 vdd.n2857 gnd 0.00713f
C5260 vdd.n2858 gnd 0.00713f
C5261 vdd.n2859 gnd 0.00713f
C5262 vdd.n2860 gnd 0.00713f
C5263 vdd.n2861 gnd 0.00713f
C5264 vdd.n2862 gnd 0.00713f
C5265 vdd.n2863 gnd 0.00713f
C5266 vdd.n2864 gnd 0.00713f
C5267 vdd.n2865 gnd 0.00713f
C5268 vdd.n2866 gnd 0.00713f
C5269 vdd.n2867 gnd 0.00713f
C5270 vdd.n2868 gnd 0.00713f
C5271 vdd.n2869 gnd 0.00713f
C5272 vdd.n2870 gnd 0.00713f
C5273 vdd.n2871 gnd 0.00713f
C5274 vdd.n2872 gnd 0.00713f
C5275 vdd.n2873 gnd 0.00713f
C5276 vdd.n2874 gnd 0.00713f
C5277 vdd.n2875 gnd 0.00713f
C5278 vdd.n2876 gnd 0.00713f
C5279 vdd.n2877 gnd 0.00713f
C5280 vdd.n2878 gnd 0.00713f
C5281 vdd.n2879 gnd 0.00713f
C5282 vdd.n2880 gnd 0.00713f
C5283 vdd.n2881 gnd 0.00713f
C5284 vdd.n2882 gnd 0.00713f
C5285 vdd.n2883 gnd 0.00713f
C5286 vdd.n2884 gnd 0.00713f
C5287 vdd.n2885 gnd 0.00713f
C5288 vdd.n2886 gnd 0.00713f
C5289 vdd.n2887 gnd 0.00713f
C5290 vdd.n2888 gnd 0.00713f
C5291 vdd.n2889 gnd 0.00519f
C5292 vdd.n2890 gnd 0.010189f
C5293 vdd.n2891 gnd 0.005504f
C5294 vdd.n2892 gnd 0.00713f
C5295 vdd.n2893 gnd 0.00713f
C5296 vdd.n2894 gnd 0.00713f
C5297 vdd.n2895 gnd 0.016433f
C5298 vdd.n2896 gnd 0.016433f
C5299 vdd.n2897 gnd 0.015441f
C5300 vdd.n2898 gnd 0.00713f
C5301 vdd.n2899 gnd 0.00713f
C5302 vdd.n2900 gnd 0.00713f
C5303 vdd.n2901 gnd 0.00713f
C5304 vdd.n2902 gnd 0.00713f
C5305 vdd.n2903 gnd 0.00713f
C5306 vdd.n2904 gnd 0.00713f
C5307 vdd.n2905 gnd 0.00713f
C5308 vdd.n2906 gnd 0.00713f
C5309 vdd.n2907 gnd 0.00713f
C5310 vdd.n2908 gnd 0.00713f
C5311 vdd.n2909 gnd 0.00713f
C5312 vdd.n2910 gnd 0.00713f
C5313 vdd.n2911 gnd 0.00713f
C5314 vdd.n2912 gnd 0.00713f
C5315 vdd.n2913 gnd 0.00713f
C5316 vdd.n2914 gnd 0.00713f
C5317 vdd.n2915 gnd 0.00713f
C5318 vdd.n2916 gnd 0.00713f
C5319 vdd.n2917 gnd 0.00713f
C5320 vdd.n2918 gnd 0.00713f
C5321 vdd.n2919 gnd 0.00713f
C5322 vdd.n2920 gnd 0.00713f
C5323 vdd.n2921 gnd 0.00713f
C5324 vdd.n2922 gnd 0.00713f
C5325 vdd.n2923 gnd 0.00713f
C5326 vdd.n2924 gnd 0.00713f
C5327 vdd.n2925 gnd 0.00713f
C5328 vdd.n2926 gnd 0.00713f
C5329 vdd.n2927 gnd 0.00713f
C5330 vdd.n2928 gnd 0.00713f
C5331 vdd.n2929 gnd 0.00713f
C5332 vdd.n2930 gnd 0.00713f
C5333 vdd.n2931 gnd 0.00713f
C5334 vdd.n2932 gnd 0.00713f
C5335 vdd.n2933 gnd 0.00713f
C5336 vdd.n2934 gnd 0.00713f
C5337 vdd.n2935 gnd 0.00713f
C5338 vdd.n2936 gnd 0.00713f
C5339 vdd.n2937 gnd 0.00713f
C5340 vdd.n2938 gnd 0.00713f
C5341 vdd.n2939 gnd 0.00713f
C5342 vdd.n2940 gnd 0.00713f
C5343 vdd.n2941 gnd 0.00713f
C5344 vdd.n2942 gnd 0.00713f
C5345 vdd.n2943 gnd 0.00713f
C5346 vdd.n2944 gnd 0.00713f
C5347 vdd.n2945 gnd 0.00713f
C5348 vdd.n2946 gnd 0.00713f
C5349 vdd.n2947 gnd 0.00713f
C5350 vdd.n2948 gnd 0.00713f
C5351 vdd.n2949 gnd 0.00713f
C5352 vdd.n2950 gnd 0.00713f
C5353 vdd.n2951 gnd 0.00713f
C5354 vdd.n2952 gnd 0.00713f
C5355 vdd.n2953 gnd 0.00713f
C5356 vdd.n2954 gnd 0.00713f
C5357 vdd.n2955 gnd 0.00713f
C5358 vdd.n2956 gnd 0.00713f
C5359 vdd.n2957 gnd 0.00713f
C5360 vdd.n2958 gnd 0.00713f
C5361 vdd.n2959 gnd 0.00713f
C5362 vdd.n2960 gnd 0.00713f
C5363 vdd.n2961 gnd 0.00713f
C5364 vdd.n2962 gnd 0.00713f
C5365 vdd.n2963 gnd 0.00713f
C5366 vdd.n2964 gnd 0.00713f
C5367 vdd.n2965 gnd 0.00713f
C5368 vdd.n2966 gnd 0.00713f
C5369 vdd.n2967 gnd 0.00713f
C5370 vdd.n2968 gnd 0.00713f
C5371 vdd.n2969 gnd 0.00713f
C5372 vdd.n2970 gnd 0.00713f
C5373 vdd.n2971 gnd 0.00713f
C5374 vdd.n2972 gnd 0.00713f
C5375 vdd.n2973 gnd 0.00713f
C5376 vdd.n2974 gnd 0.00713f
C5377 vdd.n2975 gnd 0.00713f
C5378 vdd.n2976 gnd 0.00713f
C5379 vdd.n2977 gnd 0.230369f
C5380 vdd.n2978 gnd 0.00713f
C5381 vdd.n2979 gnd 0.00713f
C5382 vdd.n2980 gnd 0.00713f
C5383 vdd.n2981 gnd 0.00713f
C5384 vdd.n2982 gnd 0.00713f
C5385 vdd.n2983 gnd 0.00713f
C5386 vdd.n2984 gnd 0.00713f
C5387 vdd.n2985 gnd 0.00713f
C5388 vdd.n2986 gnd 0.00713f
C5389 vdd.n2987 gnd 0.00713f
C5390 vdd.n2988 gnd 0.00713f
C5391 vdd.n2989 gnd 0.658962f
C5392 vdd.n2990 gnd 0.00713f
C5393 vdd.n2991 gnd 0.00713f
C5394 vdd.n2992 gnd 0.00713f
C5395 vdd.n2993 gnd 0.00713f
C5396 vdd.n2994 gnd 0.00713f
C5397 vdd.n2995 gnd 0.00713f
C5398 vdd.n2996 gnd 0.00713f
C5399 vdd.n2997 gnd 0.00713f
C5400 vdd.n2998 gnd 0.00713f
C5401 vdd.n2999 gnd 0.00713f
C5402 vdd.n3000 gnd 0.00713f
C5403 vdd.n3001 gnd 0.433951f
C5404 vdd.n3002 gnd 0.00713f
C5405 vdd.n3003 gnd 0.00713f
C5406 vdd.n3004 gnd 0.00713f
C5407 vdd.n3005 gnd 0.00713f
C5408 vdd.n3006 gnd 0.00713f
C5409 vdd.n3007 gnd 0.015441f
C5410 vdd.n3008 gnd 0.016433f
C5411 vdd.n3009 gnd 0.016433f
C5412 vdd.n3010 gnd 0.889331f
C5413 vdd.n3012 gnd 0.00713f
C5414 vdd.n3013 gnd 0.00713f
C5415 vdd.n3014 gnd 0.016433f
C5416 vdd.n3015 gnd 0.015441f
C5417 vdd.n3016 gnd 0.015441f
C5418 vdd.n3017 gnd 0.846472f
C5419 vdd.n3018 gnd 0.015441f
C5420 vdd.n3019 gnd 0.015441f
C5421 vdd.n3020 gnd 0.00713f
C5422 vdd.n3021 gnd 0.00713f
C5423 vdd.n3022 gnd 0.00713f
C5424 vdd.n3023 gnd 0.45538f
C5425 vdd.n3024 gnd 0.00713f
C5426 vdd.n3025 gnd 0.00713f
C5427 vdd.n3026 gnd 0.00713f
C5428 vdd.n3027 gnd 0.00713f
C5429 vdd.n3028 gnd 0.00713f
C5430 vdd.n3029 gnd 0.525027f
C5431 vdd.n3030 gnd 0.00713f
C5432 vdd.n3031 gnd 0.00713f
C5433 vdd.n3032 gnd 0.00713f
C5434 vdd.n3033 gnd 0.00713f
C5435 vdd.n3034 gnd 0.00713f
C5436 vdd.n3035 gnd 0.728608f
C5437 vdd.n3036 gnd 0.00713f
C5438 vdd.n3037 gnd 0.00713f
C5439 vdd.n3038 gnd 0.00713f
C5440 vdd.n3039 gnd 0.00713f
C5441 vdd.n3040 gnd 0.00713f
C5442 vdd.n3041 gnd 0.230369f
C5443 vdd.n3042 gnd 0.00713f
C5444 vdd.n3043 gnd 0.00713f
C5445 vdd.n3044 gnd 0.00713f
C5446 vdd.n3045 gnd 0.00713f
C5447 vdd.n3046 gnd 0.00713f
C5448 vdd.n3047 gnd 0.230369f
C5449 vdd.n3048 gnd 0.00713f
C5450 vdd.n3049 gnd 0.00713f
C5451 vdd.n3050 gnd 0.00713f
C5452 vdd.n3051 gnd 0.00713f
C5453 vdd.n3052 gnd 0.00713f
C5454 vdd.n3053 gnd 0.460738f
C5455 vdd.n3054 gnd 0.00713f
C5456 vdd.n3055 gnd 0.00713f
C5457 vdd.n3056 gnd 0.00713f
C5458 vdd.n3057 gnd 0.00713f
C5459 vdd.n3058 gnd 0.00713f
C5460 vdd.n3059 gnd 0.62146f
C5461 vdd.n3060 gnd 0.00713f
C5462 vdd.n3061 gnd 0.00713f
C5463 vdd.n3062 gnd 0.00713f
C5464 vdd.n3063 gnd 0.00713f
C5465 vdd.n3064 gnd 0.00713f
C5466 vdd.n3065 gnd 0.605388f
C5467 vdd.n3066 gnd 0.00713f
C5468 vdd.n3067 gnd 0.00713f
C5469 vdd.n3068 gnd 0.00713f
C5470 vdd.n3069 gnd 0.00713f
C5471 vdd.n3070 gnd 0.00713f
C5472 vdd.n3071 gnd 0.444665f
C5473 vdd.n3072 gnd 0.00713f
C5474 vdd.n3073 gnd 0.00713f
C5475 vdd.n3074 gnd 0.00713f
C5476 vdd.n3075 gnd 0.00713f
C5477 vdd.n3076 gnd 0.00713f
C5478 vdd.n3077 gnd 0.444665f
C5479 vdd.n3078 gnd 0.00713f
C5480 vdd.n3079 gnd 0.004823f
C5481 vdd.n3080 gnd 0.020653f
C5482 vdd.n3081 gnd 0.005871f
C5483 vdd.n3082 gnd 0.00713f
C5484 vdd.n3083 gnd 0.00713f
C5485 vdd.n3084 gnd 0.605388f
C5486 vdd.n3085 gnd 0.00713f
C5487 vdd.n3086 gnd 0.00713f
C5488 vdd.n3087 gnd 0.00713f
C5489 vdd.n3088 gnd 0.00713f
C5490 vdd.n3089 gnd 0.00713f
C5491 vdd.n3090 gnd 0.728608f
C5492 vdd.n3091 gnd 0.00713f
C5493 vdd.n3092 gnd 0.00713f
C5494 vdd.n3093 gnd 0.00713f
C5495 vdd.n3094 gnd 0.00713f
C5496 vdd.n3095 gnd 0.00713f
C5497 vdd.n3096 gnd 0.691107f
C5498 vdd.n3097 gnd 0.00713f
C5499 vdd.n3098 gnd 0.00713f
C5500 vdd.n3099 gnd 0.00713f
C5501 vdd.n3100 gnd 0.00713f
C5502 vdd.n3101 gnd 0.00713f
C5503 vdd.n3102 gnd 0.530384f
C5504 vdd.n3103 gnd 0.00713f
C5505 vdd.n3104 gnd 0.00713f
C5506 vdd.n3105 gnd 0.00713f
C5507 vdd.n3106 gnd 0.00713f
C5508 vdd.n3107 gnd 0.00713f
C5509 vdd.n3108 gnd 0.369662f
C5510 vdd.n3109 gnd 0.00713f
C5511 vdd.n3110 gnd 0.00713f
C5512 vdd.n3111 gnd 0.00713f
C5513 vdd.n3112 gnd 0.00713f
C5514 vdd.n3113 gnd 0.00713f
C5515 vdd.n3114 gnd 0.728608f
C5516 vdd.n3115 gnd 0.00713f
C5517 vdd.n3116 gnd 0.00713f
C5518 vdd.n3117 gnd 0.00713f
C5519 vdd.n3118 gnd 0.00713f
C5520 vdd.n3119 gnd 0.00713f
C5521 vdd.n3120 gnd 0.00713f
C5522 vdd.n3122 gnd 0.00713f
C5523 vdd.n3123 gnd 0.00713f
C5524 vdd.n3125 gnd 0.00713f
C5525 vdd.n3126 gnd 0.00713f
C5526 vdd.n3129 gnd 0.00713f
C5527 vdd.n3130 gnd 0.00713f
C5528 vdd.n3131 gnd 0.00713f
C5529 vdd.n3132 gnd 0.00713f
C5530 vdd.n3134 gnd 0.00713f
C5531 vdd.n3135 gnd 0.00713f
C5532 vdd.n3136 gnd 0.00713f
C5533 vdd.n3137 gnd 0.00713f
C5534 vdd.n3138 gnd 0.00713f
C5535 vdd.n3139 gnd 0.00713f
C5536 vdd.n3141 gnd 0.00713f
C5537 vdd.n3142 gnd 0.00713f
C5538 vdd.n3143 gnd 0.00713f
C5539 vdd.n3144 gnd 0.00713f
C5540 vdd.n3145 gnd 0.00713f
C5541 vdd.n3146 gnd 0.00713f
C5542 vdd.n3148 gnd 0.00713f
C5543 vdd.n3149 gnd 0.00713f
C5544 vdd.n3150 gnd 0.00713f
C5545 vdd.n3151 gnd 0.00713f
C5546 vdd.n3152 gnd 0.00713f
C5547 vdd.n3153 gnd 0.00713f
C5548 vdd.n3155 gnd 0.00713f
C5549 vdd.n3156 gnd 0.016433f
C5550 vdd.n3157 gnd 0.016433f
C5551 vdd.n3158 gnd 0.015441f
C5552 vdd.n3159 gnd 0.00713f
C5553 vdd.n3160 gnd 0.00713f
C5554 vdd.n3161 gnd 0.00713f
C5555 vdd.n3162 gnd 0.00713f
C5556 vdd.n3163 gnd 0.00713f
C5557 vdd.n3164 gnd 0.00713f
C5558 vdd.n3165 gnd 0.728608f
C5559 vdd.n3166 gnd 0.00713f
C5560 vdd.n3167 gnd 0.00713f
C5561 vdd.n3168 gnd 0.00713f
C5562 vdd.n3169 gnd 0.00713f
C5563 vdd.n3170 gnd 0.00713f
C5564 vdd.n3171 gnd 0.49824f
C5565 vdd.n3172 gnd 0.00713f
C5566 vdd.n3173 gnd 0.00713f
C5567 vdd.n3174 gnd 0.00713f
C5568 vdd.n3175 gnd 0.016345f
C5569 vdd.n3176 gnd 0.015529f
C5570 vdd.n3177 gnd 0.016433f
C5571 vdd.n3179 gnd 0.00713f
C5572 vdd.n3180 gnd 0.00713f
C5573 vdd.n3181 gnd 0.005504f
C5574 vdd.n3182 gnd 0.010189f
C5575 vdd.n3183 gnd 0.00519f
C5576 vdd.n3184 gnd 0.00713f
C5577 vdd.n3185 gnd 0.00713f
C5578 vdd.n3187 gnd 0.00713f
C5579 vdd.n3188 gnd 0.00713f
C5580 vdd.n3189 gnd 0.00713f
C5581 vdd.n3190 gnd 0.00713f
C5582 vdd.n3191 gnd 0.00713f
C5583 vdd.n3192 gnd 0.00713f
C5584 vdd.n3194 gnd 0.00713f
C5585 vdd.n3195 gnd 0.00713f
C5586 vdd.n3196 gnd 0.00713f
C5587 vdd.n3197 gnd 0.00713f
C5588 vdd.n3198 gnd 0.00713f
C5589 vdd.n3199 gnd 0.00713f
C5590 vdd.n3201 gnd 0.00713f
C5591 vdd.n3202 gnd 0.00713f
C5592 vdd.n3203 gnd 0.00713f
C5593 vdd.n3204 gnd 0.00713f
C5594 vdd.n3205 gnd 0.00713f
C5595 vdd.n3206 gnd 0.00713f
C5596 vdd.n3208 gnd 0.00713f
C5597 vdd.n3209 gnd 0.00713f
C5598 vdd.n3210 gnd 0.00713f
C5599 vdd.n3212 gnd 0.00713f
C5600 vdd.n3213 gnd 0.00713f
C5601 vdd.n3214 gnd 0.00713f
C5602 vdd.n3215 gnd 0.00713f
C5603 vdd.n3216 gnd 0.00713f
C5604 vdd.n3217 gnd 0.00713f
C5605 vdd.n3219 gnd 0.00713f
C5606 vdd.n3220 gnd 0.00713f
C5607 vdd.n3221 gnd 0.00713f
C5608 vdd.n3222 gnd 0.00713f
C5609 vdd.n3223 gnd 0.00713f
C5610 vdd.n3224 gnd 0.00713f
C5611 vdd.n3226 gnd 0.00713f
C5612 vdd.n3227 gnd 0.00713f
C5613 vdd.n3228 gnd 0.00713f
C5614 vdd.n3229 gnd 0.00713f
C5615 vdd.n3230 gnd 0.00713f
C5616 vdd.n3231 gnd 0.00713f
C5617 vdd.n3233 gnd 0.00713f
C5618 vdd.n3234 gnd 0.00713f
C5619 vdd.n3236 gnd 0.00713f
C5620 vdd.n3237 gnd 0.00713f
C5621 vdd.n3238 gnd 0.016433f
C5622 vdd.n3239 gnd 0.015441f
C5623 vdd.n3240 gnd 0.015441f
C5624 vdd.n3241 gnd 1.00719f
C5625 vdd.n3242 gnd 0.015441f
C5626 vdd.n3243 gnd 0.016433f
C5627 vdd.n3244 gnd 0.015529f
C5628 vdd.n3245 gnd 0.00713f
C5629 vdd.n3246 gnd 0.005504f
C5630 vdd.n3247 gnd 0.00713f
C5631 vdd.n3249 gnd 0.00713f
C5632 vdd.n3250 gnd 0.00713f
C5633 vdd.n3251 gnd 0.00713f
C5634 vdd.n3252 gnd 0.00713f
C5635 vdd.n3253 gnd 0.00713f
C5636 vdd.n3254 gnd 0.00713f
C5637 vdd.n3256 gnd 0.00713f
C5638 vdd.n3257 gnd 0.00713f
C5639 vdd.n3258 gnd 0.00713f
C5640 vdd.n3259 gnd 0.00713f
C5641 vdd.n3260 gnd 0.00713f
C5642 vdd.n3261 gnd 0.00713f
C5643 vdd.n3263 gnd 0.00713f
C5644 vdd.n3264 gnd 0.00713f
C5645 vdd.n3265 gnd 0.00713f
C5646 vdd.n3266 gnd 0.00713f
C5647 vdd.n3267 gnd 0.00713f
C5648 vdd.n3268 gnd 0.00713f
C5649 vdd.n3270 gnd 0.00713f
C5650 vdd.n3271 gnd 0.00713f
C5651 vdd.n3273 gnd 0.00713f
C5652 vdd.n3274 gnd 0.033466f
C5653 vdd.n3275 gnd 0.957817f
C5654 vdd.n3277 gnd 0.00443f
C5655 vdd.n3278 gnd 0.008439f
C5656 vdd.n3279 gnd 0.010485f
C5657 vdd.n3280 gnd 0.010485f
C5658 vdd.n3281 gnd 0.008439f
C5659 vdd.n3282 gnd 0.008439f
C5660 vdd.n3283 gnd 0.010485f
C5661 vdd.n3284 gnd 0.010485f
C5662 vdd.n3285 gnd 0.008439f
C5663 vdd.n3286 gnd 0.008439f
C5664 vdd.n3287 gnd 0.010485f
C5665 vdd.n3288 gnd 0.010485f
C5666 vdd.n3289 gnd 0.008439f
C5667 vdd.n3290 gnd 0.008439f
C5668 vdd.n3291 gnd 0.010485f
C5669 vdd.n3292 gnd 0.010485f
C5670 vdd.n3293 gnd 0.008439f
C5671 vdd.n3294 gnd 0.008439f
C5672 vdd.n3295 gnd 0.010485f
C5673 vdd.n3296 gnd 0.010485f
C5674 vdd.n3297 gnd 0.008439f
C5675 vdd.n3298 gnd 0.008439f
C5676 vdd.n3299 gnd 0.010485f
C5677 vdd.n3300 gnd 0.010485f
C5678 vdd.n3301 gnd 0.008439f
C5679 vdd.n3302 gnd 0.008439f
C5680 vdd.n3303 gnd 0.010485f
C5681 vdd.n3304 gnd 0.010485f
C5682 vdd.n3305 gnd 0.008439f
C5683 vdd.n3306 gnd 0.008439f
C5684 vdd.n3307 gnd 0.010485f
C5685 vdd.n3308 gnd 0.010485f
C5686 vdd.n3309 gnd 0.008439f
C5687 vdd.n3310 gnd 0.008439f
C5688 vdd.n3311 gnd 0.010485f
C5689 vdd.n3312 gnd 0.010485f
C5690 vdd.n3313 gnd 0.008439f
C5691 vdd.n3314 gnd 0.010485f
C5692 vdd.n3315 gnd 0.010485f
C5693 vdd.n3316 gnd 0.008439f
C5694 vdd.n3317 gnd 0.010485f
C5695 vdd.n3318 gnd 0.010485f
C5696 vdd.n3319 gnd 0.010485f
C5697 vdd.n3320 gnd 0.017215f
C5698 vdd.n3321 gnd 0.010485f
C5699 vdd.n3322 gnd 0.010485f
C5700 vdd.n3323 gnd 0.005738f
C5701 vdd.n3324 gnd 0.008439f
C5702 vdd.n3325 gnd 0.010485f
C5703 vdd.n3326 gnd 0.010485f
C5704 vdd.n3327 gnd 0.008439f
C5705 vdd.n3328 gnd 0.008439f
C5706 vdd.n3329 gnd 0.010485f
C5707 vdd.n3330 gnd 0.010485f
C5708 vdd.n3331 gnd 0.008439f
C5709 vdd.n3332 gnd 0.008439f
C5710 vdd.n3333 gnd 0.010485f
C5711 vdd.n3334 gnd 0.010485f
C5712 vdd.n3335 gnd 0.008439f
C5713 vdd.n3336 gnd 0.008439f
C5714 vdd.n3337 gnd 0.010485f
C5715 vdd.n3338 gnd 0.010485f
C5716 vdd.n3339 gnd 0.008439f
C5717 vdd.n3340 gnd 0.008439f
C5718 vdd.n3341 gnd 0.010485f
C5719 vdd.n3342 gnd 0.010485f
C5720 vdd.n3343 gnd 0.008439f
C5721 vdd.n3344 gnd 0.008439f
C5722 vdd.n3345 gnd 0.010485f
C5723 vdd.n3346 gnd 0.010485f
C5724 vdd.n3347 gnd 0.008439f
C5725 vdd.n3348 gnd 0.008439f
C5726 vdd.n3349 gnd 0.010485f
C5727 vdd.n3350 gnd 0.010485f
C5728 vdd.n3351 gnd 0.008439f
C5729 vdd.n3352 gnd 0.008439f
C5730 vdd.n3353 gnd 0.010485f
C5731 vdd.n3354 gnd 0.010485f
C5732 vdd.n3355 gnd 0.008439f
C5733 vdd.n3356 gnd 0.008439f
C5734 vdd.n3357 gnd 0.010485f
C5735 vdd.n3358 gnd 0.010485f
C5736 vdd.n3359 gnd 0.008439f
C5737 vdd.n3360 gnd 0.010485f
C5738 vdd.n3361 gnd 0.010485f
C5739 vdd.n3362 gnd 0.008439f
C5740 vdd.n3363 gnd 0.010485f
C5741 vdd.n3364 gnd 0.010485f
C5742 vdd.n3365 gnd 0.010485f
C5743 vdd.t38 gnd 0.128989f
C5744 vdd.t39 gnd 0.137854f
C5745 vdd.t37 gnd 0.168458f
C5746 vdd.n3366 gnd 0.215939f
C5747 vdd.n3367 gnd 0.181428f
C5748 vdd.n3368 gnd 0.017215f
C5749 vdd.n3369 gnd 0.010485f
C5750 vdd.n3370 gnd 0.010485f
C5751 vdd.n3371 gnd 0.007046f
C5752 vdd.n3372 gnd 0.008439f
C5753 vdd.n3373 gnd 0.010485f
C5754 vdd.n3374 gnd 0.010485f
C5755 vdd.n3375 gnd 0.008439f
C5756 vdd.n3376 gnd 0.008439f
C5757 vdd.n3377 gnd 0.010485f
C5758 vdd.n3378 gnd 0.010485f
C5759 vdd.n3379 gnd 0.008439f
C5760 vdd.n3380 gnd 0.008439f
C5761 vdd.n3381 gnd 0.010485f
C5762 vdd.n3382 gnd 0.010485f
C5763 vdd.n3383 gnd 0.008439f
C5764 vdd.n3384 gnd 0.008439f
C5765 vdd.n3385 gnd 0.010485f
C5766 vdd.n3386 gnd 0.010485f
C5767 vdd.n3387 gnd 0.008439f
C5768 vdd.n3388 gnd 0.008439f
C5769 vdd.n3389 gnd 0.010485f
C5770 vdd.n3390 gnd 0.010485f
C5771 vdd.n3391 gnd 0.008439f
C5772 vdd.n3392 gnd 0.008439f
C5773 vdd.n3393 gnd 0.010485f
C5774 vdd.n3394 gnd 0.010485f
C5775 vdd.n3395 gnd 0.008439f
C5776 vdd.n3396 gnd 0.008439f
C5777 vdd.n3398 gnd 0.957817f
C5778 vdd.n3400 gnd 0.008439f
C5779 vdd.n3401 gnd 0.008439f
C5780 vdd.n3402 gnd 0.007004f
C5781 vdd.n3403 gnd 0.025907f
C5782 vdd.n3405 gnd 11.304099f
C5783 vdd.n3406 gnd 0.025907f
C5784 vdd.n3407 gnd 0.004008f
C5785 vdd.n3408 gnd 0.025907f
C5786 vdd.n3409 gnd 0.025363f
C5787 vdd.n3410 gnd 0.010485f
C5788 vdd.n3411 gnd 0.008439f
C5789 vdd.n3412 gnd 0.010485f
C5790 vdd.n3413 gnd 0.648247f
C5791 vdd.n3414 gnd 0.010485f
C5792 vdd.n3415 gnd 0.008439f
C5793 vdd.n3416 gnd 0.010485f
C5794 vdd.n3417 gnd 0.010485f
C5795 vdd.n3418 gnd 0.010485f
C5796 vdd.n3419 gnd 0.008439f
C5797 vdd.n3420 gnd 0.010485f
C5798 vdd.n3421 gnd 1.07148f
C5799 vdd.n3422 gnd 0.010485f
C5800 vdd.n3423 gnd 0.008439f
C5801 vdd.n3424 gnd 0.010485f
C5802 vdd.n3425 gnd 0.010485f
C5803 vdd.n3426 gnd 0.010485f
C5804 vdd.n3427 gnd 0.008439f
C5805 vdd.n3428 gnd 0.010485f
C5806 vdd.n3429 gnd 0.691107f
C5807 vdd.n3430 gnd 0.733966f
C5808 vdd.n3431 gnd 0.010485f
C5809 vdd.n3432 gnd 0.008439f
C5810 vdd.n3433 gnd 0.010485f
C5811 vdd.n3434 gnd 0.010485f
C5812 vdd.n3435 gnd 0.010485f
C5813 vdd.n3436 gnd 0.008439f
C5814 vdd.n3437 gnd 0.010485f
C5815 vdd.n3438 gnd 0.889331f
C5816 vdd.n3439 gnd 0.010485f
C5817 vdd.n3440 gnd 0.008439f
C5818 vdd.n3441 gnd 0.010485f
C5819 vdd.n3442 gnd 0.010485f
C5820 vdd.n3443 gnd 0.010485f
C5821 vdd.n3444 gnd 0.008439f
C5822 vdd.n3445 gnd 0.010485f
C5823 vdd.t163 gnd 0.535742f
C5824 vdd.n3446 gnd 0.862544f
C5825 vdd.n3447 gnd 0.010485f
C5826 vdd.n3448 gnd 0.008439f
C5827 vdd.n3449 gnd 0.010485f
C5828 vdd.n3450 gnd 0.010485f
C5829 vdd.n3451 gnd 0.010485f
C5830 vdd.n3452 gnd 0.008439f
C5831 vdd.n3453 gnd 0.010485f
C5832 vdd.n3454 gnd 0.680392f
C5833 vdd.n3455 gnd 0.010485f
C5834 vdd.n3456 gnd 0.008439f
C5835 vdd.n3457 gnd 0.010485f
C5836 vdd.n3458 gnd 0.010485f
C5837 vdd.n3459 gnd 0.010485f
C5838 vdd.n3460 gnd 0.008439f
C5839 vdd.n3461 gnd 0.010485f
C5840 vdd.n3462 gnd 0.851829f
C5841 vdd.n3463 gnd 0.573243f
C5842 vdd.n3464 gnd 0.010485f
C5843 vdd.n3465 gnd 0.008439f
C5844 vdd.n3466 gnd 0.010485f
C5845 vdd.n3467 gnd 0.010485f
C5846 vdd.n3468 gnd 0.010485f
C5847 vdd.n3469 gnd 0.008439f
C5848 vdd.n3470 gnd 0.010485f
C5849 vdd.n3471 gnd 0.755396f
C5850 vdd.n3472 gnd 0.010485f
C5851 vdd.n3473 gnd 0.008439f
C5852 vdd.n3474 gnd 0.010485f
C5853 vdd.n3475 gnd 0.010485f
C5854 vdd.n3476 gnd 0.010485f
C5855 vdd.n3477 gnd 0.010485f
C5856 vdd.n3478 gnd 0.010485f
C5857 vdd.n3479 gnd 0.008439f
C5858 vdd.n3480 gnd 0.008439f
C5859 vdd.n3481 gnd 0.010485f
C5860 vdd.t256 gnd 0.535742f
C5861 vdd.n3482 gnd 0.889331f
C5862 vdd.n3483 gnd 0.010485f
C5863 vdd.n3484 gnd 0.008439f
C5864 vdd.n3485 gnd 0.010485f
C5865 vdd.n3486 gnd 0.010485f
C5866 vdd.n3487 gnd 0.010485f
C5867 vdd.n3488 gnd 0.008439f
C5868 vdd.n3489 gnd 0.010485f
C5869 vdd.n3490 gnd 0.841114f
C5870 vdd.n3491 gnd 0.010485f
C5871 vdd.n3492 gnd 0.010485f
C5872 vdd.n3493 gnd 0.008439f
C5873 vdd.n3494 gnd 0.008439f
C5874 vdd.n3495 gnd 0.010485f
C5875 vdd.n3496 gnd 0.010485f
C5876 vdd.n3497 gnd 0.010485f
C5877 vdd.n3498 gnd 0.008439f
C5878 vdd.n3499 gnd 0.010485f
C5879 vdd.n3500 gnd 0.008439f
C5880 vdd.n3501 gnd 0.008439f
C5881 vdd.n3502 gnd 0.010485f
C5882 vdd.n3503 gnd 0.010485f
C5883 vdd.n3504 gnd 0.010485f
C5884 vdd.n3505 gnd 0.008439f
C5885 vdd.n3506 gnd 0.010485f
C5886 vdd.n3507 gnd 0.008439f
C5887 vdd.n3508 gnd 0.008439f
C5888 vdd.n3509 gnd 0.010485f
C5889 vdd.n3510 gnd 0.010485f
C5890 vdd.n3511 gnd 0.010485f
C5891 vdd.n3512 gnd 0.008439f
C5892 vdd.n3513 gnd 0.889331f
C5893 vdd.n3514 gnd 0.010485f
C5894 vdd.n3515 gnd 0.008439f
C5895 vdd.n3516 gnd 0.008439f
C5896 vdd.n3517 gnd 0.010485f
C5897 vdd.n3518 gnd 0.010485f
C5898 vdd.n3519 gnd 0.010485f
C5899 vdd.n3520 gnd 0.008439f
C5900 vdd.n3521 gnd 0.010485f
C5901 vdd.n3522 gnd 0.008439f
C5902 vdd.n3523 gnd 0.008439f
C5903 vdd.n3524 gnd 0.010485f
C5904 vdd.n3525 gnd 0.010485f
C5905 vdd.n3526 gnd 0.010485f
C5906 vdd.n3527 gnd 0.008439f
C5907 vdd.n3528 gnd 0.010485f
C5908 vdd.n3529 gnd 0.008439f
C5909 vdd.n3530 gnd 0.007004f
C5910 vdd.n3531 gnd 0.025363f
C5911 vdd.n3532 gnd 0.025907f
C5912 vdd.n3533 gnd 0.004008f
C5913 vdd.n3534 gnd 0.025907f
C5914 vdd.n3536 gnd 2.53941f
C5915 vdd.n3537 gnd 1.58044f
C5916 vdd.n3538 gnd 0.025363f
C5917 vdd.n3539 gnd 0.007004f
C5918 vdd.n3540 gnd 0.008439f
C5919 vdd.n3541 gnd 0.008439f
C5920 vdd.n3542 gnd 0.010485f
C5921 vdd.n3543 gnd 1.07148f
C5922 vdd.n3544 gnd 1.07148f
C5923 vdd.n3545 gnd 0.980407f
C5924 vdd.n3546 gnd 0.010485f
C5925 vdd.n3547 gnd 0.008439f
C5926 vdd.n3548 gnd 0.008439f
C5927 vdd.n3549 gnd 0.008439f
C5928 vdd.n3550 gnd 0.010485f
C5929 vdd.n3551 gnd 0.798255f
C5930 vdd.t280 gnd 0.535742f
C5931 vdd.n3552 gnd 0.80897f
C5932 vdd.n3553 gnd 0.616103f
C5933 vdd.n3554 gnd 0.010485f
C5934 vdd.n3555 gnd 0.008439f
C5935 vdd.n3556 gnd 0.008439f
C5936 vdd.n3557 gnd 0.008439f
C5937 vdd.n3558 gnd 0.010485f
C5938 vdd.n3559 gnd 0.637532f
C5939 vdd.n3560 gnd 0.78754f
C5940 vdd.t157 gnd 0.535742f
C5941 vdd.n3561 gnd 0.819685f
C5942 vdd.n3562 gnd 0.010485f
C5943 vdd.n3563 gnd 0.008439f
C5944 vdd.n3564 gnd 0.008439f
C5945 vdd.n3565 gnd 0.008439f
C5946 vdd.n3566 gnd 0.010485f
C5947 vdd.n3567 gnd 0.889331f
C5948 vdd.t198 gnd 0.535742f
C5949 vdd.n3568 gnd 0.648247f
C5950 vdd.n3569 gnd 0.776825f
C5951 vdd.n3570 gnd 0.010485f
C5952 vdd.n3571 gnd 0.008439f
C5953 vdd.n3572 gnd 0.008439f
C5954 vdd.n3573 gnd 0.008439f
C5955 vdd.n3574 gnd 0.010485f
C5956 vdd.n3575 gnd 0.594673f
C5957 vdd.t210 gnd 0.535742f
C5958 vdd.n3576 gnd 0.889331f
C5959 vdd.t225 gnd 0.535742f
C5960 vdd.n3577 gnd 0.658962f
C5961 vdd.n3578 gnd 0.010485f
C5962 vdd.n3579 gnd 0.008439f
C5963 vdd.n3580 gnd 0.008058f
C5964 vdd.n3581 gnd 0.618425f
C5965 vdd.n3582 gnd 2.93502f
C5966 a_n8964_8799.n0 gnd 0.875393f
C5967 a_n8964_8799.n1 gnd 3.59739f
C5968 a_n8964_8799.n2 gnd 3.33951f
C5969 a_n8964_8799.n3 gnd 1.65962f
C5970 a_n8964_8799.n4 gnd 0.207089f
C5971 a_n8964_8799.n5 gnd 0.28436f
C5972 a_n8964_8799.n6 gnd 0.207089f
C5973 a_n8964_8799.n7 gnd 0.207089f
C5974 a_n8964_8799.n8 gnd 0.207089f
C5975 a_n8964_8799.n9 gnd 0.207089f
C5976 a_n8964_8799.n10 gnd 0.207089f
C5977 a_n8964_8799.n11 gnd 0.215335f
C5978 a_n8964_8799.n12 gnd 0.207089f
C5979 a_n8964_8799.n13 gnd 0.28436f
C5980 a_n8964_8799.n14 gnd 0.207089f
C5981 a_n8964_8799.n15 gnd 0.207089f
C5982 a_n8964_8799.n16 gnd 0.207089f
C5983 a_n8964_8799.n17 gnd 0.207089f
C5984 a_n8964_8799.n18 gnd 0.207089f
C5985 a_n8964_8799.n19 gnd 0.215335f
C5986 a_n8964_8799.n20 gnd 0.207089f
C5987 a_n8964_8799.n21 gnd 0.448852f
C5988 a_n8964_8799.n22 gnd 0.207089f
C5989 a_n8964_8799.n23 gnd 0.207089f
C5990 a_n8964_8799.n24 gnd 0.207089f
C5991 a_n8964_8799.n25 gnd 0.207089f
C5992 a_n8964_8799.n26 gnd 0.207089f
C5993 a_n8964_8799.n27 gnd 0.215335f
C5994 a_n8964_8799.n28 gnd 0.207089f
C5995 a_n8964_8799.n29 gnd 0.31888f
C5996 a_n8964_8799.n30 gnd 0.207089f
C5997 a_n8964_8799.n31 gnd 0.207089f
C5998 a_n8964_8799.n32 gnd 0.207089f
C5999 a_n8964_8799.n33 gnd 0.207089f
C6000 a_n8964_8799.n34 gnd 0.207089f
C6001 a_n8964_8799.n35 gnd 0.180816f
C6002 a_n8964_8799.n36 gnd 0.207089f
C6003 a_n8964_8799.n37 gnd 0.31888f
C6004 a_n8964_8799.n38 gnd 0.207089f
C6005 a_n8964_8799.n39 gnd 0.207089f
C6006 a_n8964_8799.n40 gnd 0.207089f
C6007 a_n8964_8799.n41 gnd 0.207089f
C6008 a_n8964_8799.n42 gnd 0.207089f
C6009 a_n8964_8799.n43 gnd 0.180816f
C6010 a_n8964_8799.n44 gnd 0.207089f
C6011 a_n8964_8799.n45 gnd 0.31888f
C6012 a_n8964_8799.n46 gnd 0.207089f
C6013 a_n8964_8799.n47 gnd 0.207089f
C6014 a_n8964_8799.n48 gnd 0.207089f
C6015 a_n8964_8799.n49 gnd 0.207089f
C6016 a_n8964_8799.n50 gnd 0.207089f
C6017 a_n8964_8799.n51 gnd 0.345308f
C6018 a_n8964_8799.n52 gnd 1.5178f
C6019 a_n8964_8799.n53 gnd 3.95401f
C6020 a_n8964_8799.n54 gnd 2.74076f
C6021 a_n8964_8799.n55 gnd 1.51779f
C6022 a_n8964_8799.n56 gnd 0.249316f
C6023 a_n8964_8799.n57 gnd 0.003645f
C6024 a_n8964_8799.n58 gnd 0.009608f
C6025 a_n8964_8799.n59 gnd 0.010498f
C6026 a_n8964_8799.n60 gnd 0.005547f
C6027 a_n8964_8799.n62 gnd 0.004654f
C6028 a_n8964_8799.n63 gnd 0.010066f
C6029 a_n8964_8799.n64 gnd 0.010066f
C6030 a_n8964_8799.n65 gnd 0.004654f
C6031 a_n8964_8799.n67 gnd 0.005547f
C6032 a_n8964_8799.n68 gnd 0.010498f
C6033 a_n8964_8799.n69 gnd 0.009608f
C6034 a_n8964_8799.n70 gnd 0.003645f
C6035 a_n8964_8799.n71 gnd 0.249316f
C6036 a_n8964_8799.n72 gnd 0.003645f
C6037 a_n8964_8799.n73 gnd 0.009608f
C6038 a_n8964_8799.n74 gnd 0.010498f
C6039 a_n8964_8799.n75 gnd 0.005547f
C6040 a_n8964_8799.n77 gnd 0.004654f
C6041 a_n8964_8799.n78 gnd 0.010066f
C6042 a_n8964_8799.n79 gnd 0.010066f
C6043 a_n8964_8799.n80 gnd 0.004654f
C6044 a_n8964_8799.n82 gnd 0.005547f
C6045 a_n8964_8799.n83 gnd 0.010498f
C6046 a_n8964_8799.n84 gnd 0.009608f
C6047 a_n8964_8799.n85 gnd 0.003645f
C6048 a_n8964_8799.n86 gnd 0.249316f
C6049 a_n8964_8799.n87 gnd 0.003645f
C6050 a_n8964_8799.n88 gnd 0.009608f
C6051 a_n8964_8799.n89 gnd 0.010498f
C6052 a_n8964_8799.n90 gnd 0.005547f
C6053 a_n8964_8799.n92 gnd 0.004654f
C6054 a_n8964_8799.n93 gnd 0.010066f
C6055 a_n8964_8799.n94 gnd 0.010066f
C6056 a_n8964_8799.n95 gnd 0.004654f
C6057 a_n8964_8799.n97 gnd 0.005547f
C6058 a_n8964_8799.n98 gnd 0.010498f
C6059 a_n8964_8799.n99 gnd 0.009608f
C6060 a_n8964_8799.n100 gnd 0.003645f
C6061 a_n8964_8799.n101 gnd 0.003645f
C6062 a_n8964_8799.n102 gnd 0.009608f
C6063 a_n8964_8799.n103 gnd 0.010498f
C6064 a_n8964_8799.n104 gnd 0.005547f
C6065 a_n8964_8799.n106 gnd 0.004654f
C6066 a_n8964_8799.n107 gnd 0.010066f
C6067 a_n8964_8799.n108 gnd 0.010066f
C6068 a_n8964_8799.n109 gnd 0.004654f
C6069 a_n8964_8799.n111 gnd 0.005547f
C6070 a_n8964_8799.n112 gnd 0.010498f
C6071 a_n8964_8799.n113 gnd 0.009608f
C6072 a_n8964_8799.n114 gnd 0.003645f
C6073 a_n8964_8799.n115 gnd 0.249316f
C6074 a_n8964_8799.n116 gnd 0.003645f
C6075 a_n8964_8799.n117 gnd 0.009608f
C6076 a_n8964_8799.n118 gnd 0.010498f
C6077 a_n8964_8799.n119 gnd 0.005547f
C6078 a_n8964_8799.n121 gnd 0.004654f
C6079 a_n8964_8799.n122 gnd 0.010066f
C6080 a_n8964_8799.n123 gnd 0.010066f
C6081 a_n8964_8799.n124 gnd 0.004654f
C6082 a_n8964_8799.n126 gnd 0.005547f
C6083 a_n8964_8799.n127 gnd 0.010498f
C6084 a_n8964_8799.n128 gnd 0.009608f
C6085 a_n8964_8799.n129 gnd 0.003645f
C6086 a_n8964_8799.n130 gnd 0.249316f
C6087 a_n8964_8799.n131 gnd 0.003645f
C6088 a_n8964_8799.n132 gnd 0.009608f
C6089 a_n8964_8799.n133 gnd 0.010498f
C6090 a_n8964_8799.n134 gnd 0.005547f
C6091 a_n8964_8799.n136 gnd 0.004654f
C6092 a_n8964_8799.n137 gnd 0.010066f
C6093 a_n8964_8799.n138 gnd 0.010066f
C6094 a_n8964_8799.n139 gnd 0.004654f
C6095 a_n8964_8799.n141 gnd 0.005547f
C6096 a_n8964_8799.n142 gnd 0.010498f
C6097 a_n8964_8799.n143 gnd 0.009608f
C6098 a_n8964_8799.n144 gnd 0.003645f
C6099 a_n8964_8799.n145 gnd 0.249316f
C6100 a_n8964_8799.t8 gnd 0.143639f
C6101 a_n8964_8799.t4 gnd 0.143639f
C6102 a_n8964_8799.t29 gnd 0.143639f
C6103 a_n8964_8799.n146 gnd 1.1329f
C6104 a_n8964_8799.t21 gnd 0.143639f
C6105 a_n8964_8799.t7 gnd 0.143639f
C6106 a_n8964_8799.n147 gnd 1.13104f
C6107 a_n8964_8799.t1 gnd 0.143639f
C6108 a_n8964_8799.t2 gnd 0.143639f
C6109 a_n8964_8799.n148 gnd 1.13104f
C6110 a_n8964_8799.t34 gnd 0.143639f
C6111 a_n8964_8799.t24 gnd 0.143639f
C6112 a_n8964_8799.n149 gnd 1.13104f
C6113 a_n8964_8799.t16 gnd 0.143639f
C6114 a_n8964_8799.t22 gnd 0.143639f
C6115 a_n8964_8799.n150 gnd 1.13104f
C6116 a_n8964_8799.t20 gnd 0.111719f
C6117 a_n8964_8799.t26 gnd 0.111719f
C6118 a_n8964_8799.n151 gnd 0.990103f
C6119 a_n8964_8799.t15 gnd 0.111719f
C6120 a_n8964_8799.t18 gnd 0.111719f
C6121 a_n8964_8799.n152 gnd 0.987192f
C6122 a_n8964_8799.t3 gnd 0.111719f
C6123 a_n8964_8799.t37 gnd 0.111719f
C6124 a_n8964_8799.n153 gnd 0.987192f
C6125 a_n8964_8799.t36 gnd 0.111719f
C6126 a_n8964_8799.t33 gnd 0.111719f
C6127 a_n8964_8799.n154 gnd 0.990102f
C6128 a_n8964_8799.t6 gnd 0.111719f
C6129 a_n8964_8799.t12 gnd 0.111719f
C6130 a_n8964_8799.n155 gnd 0.987191f
C6131 a_n8964_8799.t14 gnd 0.111719f
C6132 a_n8964_8799.t23 gnd 0.111719f
C6133 a_n8964_8799.n156 gnd 0.987191f
C6134 a_n8964_8799.t32 gnd 0.111719f
C6135 a_n8964_8799.t9 gnd 0.111719f
C6136 a_n8964_8799.n157 gnd 0.990102f
C6137 a_n8964_8799.t11 gnd 0.111719f
C6138 a_n8964_8799.t13 gnd 0.111719f
C6139 a_n8964_8799.n158 gnd 0.987191f
C6140 a_n8964_8799.t39 gnd 0.111719f
C6141 a_n8964_8799.t10 gnd 0.111719f
C6142 a_n8964_8799.n159 gnd 0.987192f
C6143 a_n8964_8799.t19 gnd 0.111719f
C6144 a_n8964_8799.t30 gnd 0.111719f
C6145 a_n8964_8799.n160 gnd 0.987192f
C6146 a_n8964_8799.t73 gnd 0.595595f
C6147 a_n8964_8799.n161 gnd 0.268145f
C6148 a_n8964_8799.t118 gnd 0.595595f
C6149 a_n8964_8799.t141 gnd 0.595595f
C6150 a_n8964_8799.n162 gnd 0.270066f
C6151 a_n8964_8799.t86 gnd 0.595595f
C6152 a_n8964_8799.t89 gnd 0.595595f
C6153 a_n8964_8799.n163 gnd 0.263291f
C6154 a_n8964_8799.t142 gnd 0.595595f
C6155 a_n8964_8799.t147 gnd 0.595595f
C6156 a_n8964_8799.n164 gnd 0.267255f
C6157 a_n8964_8799.t72 gnd 0.595595f
C6158 a_n8964_8799.t117 gnd 0.595595f
C6159 a_n8964_8799.t87 gnd 0.606868f
C6160 a_n8964_8799.n165 gnd 0.249678f
C6161 a_n8964_8799.n166 gnd 0.270437f
C6162 a_n8964_8799.t44 gnd 0.595595f
C6163 a_n8964_8799.n167 gnd 0.268145f
C6164 a_n8964_8799.n168 gnd 0.263929f
C6165 a_n8964_8799.t110 gnd 0.595595f
C6166 a_n8964_8799.n169 gnd 0.262653f
C6167 a_n8964_8799.t70 gnd 0.595595f
C6168 a_n8964_8799.n170 gnd 0.269811f
C6169 a_n8964_8799.t105 gnd 0.595595f
C6170 a_n8964_8799.n171 gnd 0.270066f
C6171 a_n8964_8799.n172 gnd 0.267686f
C6172 a_n8964_8799.t143 gnd 0.595595f
C6173 a_n8964_8799.n173 gnd 0.263291f
C6174 a_n8964_8799.t121 gnd 0.595595f
C6175 a_n8964_8799.n174 gnd 0.267686f
C6176 a_n8964_8799.n175 gnd 0.269811f
C6177 a_n8964_8799.t88 gnd 0.595595f
C6178 a_n8964_8799.n176 gnd 0.267255f
C6179 a_n8964_8799.n177 gnd 0.262653f
C6180 a_n8964_8799.t71 gnd 0.595595f
C6181 a_n8964_8799.n178 gnd 0.263929f
C6182 a_n8964_8799.t114 gnd 0.595595f
C6183 a_n8964_8799.n179 gnd 0.270437f
C6184 a_n8964_8799.t40 gnd 0.606858f
C6185 a_n8964_8799.t84 gnd 0.595595f
C6186 a_n8964_8799.n180 gnd 0.268145f
C6187 a_n8964_8799.t135 gnd 0.595595f
C6188 a_n8964_8799.t154 gnd 0.595595f
C6189 a_n8964_8799.n181 gnd 0.270066f
C6190 a_n8964_8799.t96 gnd 0.595595f
C6191 a_n8964_8799.t101 gnd 0.595595f
C6192 a_n8964_8799.n182 gnd 0.263291f
C6193 a_n8964_8799.t156 gnd 0.595595f
C6194 a_n8964_8799.t159 gnd 0.595595f
C6195 a_n8964_8799.n183 gnd 0.267255f
C6196 a_n8964_8799.t83 gnd 0.595595f
C6197 a_n8964_8799.t134 gnd 0.595595f
C6198 a_n8964_8799.t97 gnd 0.606868f
C6199 a_n8964_8799.n184 gnd 0.249678f
C6200 a_n8964_8799.n185 gnd 0.270437f
C6201 a_n8964_8799.t56 gnd 0.595595f
C6202 a_n8964_8799.n186 gnd 0.268145f
C6203 a_n8964_8799.n187 gnd 0.263929f
C6204 a_n8964_8799.t125 gnd 0.595595f
C6205 a_n8964_8799.n188 gnd 0.262653f
C6206 a_n8964_8799.t79 gnd 0.595595f
C6207 a_n8964_8799.n189 gnd 0.269811f
C6208 a_n8964_8799.t119 gnd 0.595595f
C6209 a_n8964_8799.n190 gnd 0.270066f
C6210 a_n8964_8799.n191 gnd 0.267686f
C6211 a_n8964_8799.t158 gnd 0.595595f
C6212 a_n8964_8799.n192 gnd 0.263291f
C6213 a_n8964_8799.t138 gnd 0.595595f
C6214 a_n8964_8799.n193 gnd 0.267686f
C6215 a_n8964_8799.n194 gnd 0.269811f
C6216 a_n8964_8799.t98 gnd 0.595595f
C6217 a_n8964_8799.n195 gnd 0.267255f
C6218 a_n8964_8799.n196 gnd 0.262653f
C6219 a_n8964_8799.t82 gnd 0.595595f
C6220 a_n8964_8799.n197 gnd 0.263929f
C6221 a_n8964_8799.t132 gnd 0.595595f
C6222 a_n8964_8799.n198 gnd 0.270437f
C6223 a_n8964_8799.t52 gnd 0.606858f
C6224 a_n8964_8799.n199 gnd 0.895395f
C6225 a_n8964_8799.t120 gnd 0.595595f
C6226 a_n8964_8799.n200 gnd 0.268145f
C6227 a_n8964_8799.t102 gnd 0.595595f
C6228 a_n8964_8799.t144 gnd 0.595595f
C6229 a_n8964_8799.n201 gnd 0.270066f
C6230 a_n8964_8799.t62 gnd 0.595595f
C6231 a_n8964_8799.t137 gnd 0.595595f
C6232 a_n8964_8799.n202 gnd 0.263291f
C6233 a_n8964_8799.t115 gnd 0.595595f
C6234 a_n8964_8799.t75 gnd 0.595595f
C6235 a_n8964_8799.n203 gnd 0.267255f
C6236 a_n8964_8799.t60 gnd 0.595595f
C6237 a_n8964_8799.t45 gnd 0.595595f
C6238 a_n8964_8799.t90 gnd 0.606868f
C6239 a_n8964_8799.n204 gnd 0.249678f
C6240 a_n8964_8799.n205 gnd 0.270437f
C6241 a_n8964_8799.t106 gnd 0.595595f
C6242 a_n8964_8799.n206 gnd 0.268145f
C6243 a_n8964_8799.n207 gnd 0.263929f
C6244 a_n8964_8799.t127 gnd 0.595595f
C6245 a_n8964_8799.n208 gnd 0.262653f
C6246 a_n8964_8799.t99 gnd 0.595595f
C6247 a_n8964_8799.n209 gnd 0.269811f
C6248 a_n8964_8799.t53 gnd 0.595595f
C6249 a_n8964_8799.n210 gnd 0.270066f
C6250 a_n8964_8799.n211 gnd 0.267686f
C6251 a_n8964_8799.t94 gnd 0.595595f
C6252 a_n8964_8799.n212 gnd 0.263291f
C6253 a_n8964_8799.t80 gnd 0.595595f
C6254 a_n8964_8799.n213 gnd 0.267686f
C6255 a_n8964_8799.n214 gnd 0.269811f
C6256 a_n8964_8799.t41 gnd 0.595595f
C6257 a_n8964_8799.n215 gnd 0.267255f
C6258 a_n8964_8799.n216 gnd 0.262653f
C6259 a_n8964_8799.t146 gnd 0.595595f
C6260 a_n8964_8799.n217 gnd 0.263929f
C6261 a_n8964_8799.t153 gnd 0.595595f
C6262 a_n8964_8799.n218 gnd 0.270437f
C6263 a_n8964_8799.t95 gnd 0.606858f
C6264 a_n8964_8799.n219 gnd 1.74676f
C6265 a_n8964_8799.t107 gnd 0.606858f
C6266 a_n8964_8799.t43 gnd 0.595595f
C6267 a_n8964_8799.t113 gnd 0.595595f
C6268 a_n8964_8799.n220 gnd 0.268145f
C6269 a_n8964_8799.t111 gnd 0.595595f
C6270 a_n8964_8799.t49 gnd 0.595595f
C6271 a_n8964_8799.t47 gnd 0.595595f
C6272 a_n8964_8799.n221 gnd 0.267255f
C6273 a_n8964_8799.t133 gnd 0.595595f
C6274 a_n8964_8799.t65 gnd 0.595595f
C6275 a_n8964_8799.t51 gnd 0.595595f
C6276 a_n8964_8799.n222 gnd 0.267686f
C6277 a_n8964_8799.t139 gnd 0.595595f
C6278 a_n8964_8799.t91 gnd 0.595595f
C6279 a_n8964_8799.t66 gnd 0.595595f
C6280 a_n8964_8799.n223 gnd 0.267686f
C6281 a_n8964_8799.t157 gnd 0.595595f
C6282 a_n8964_8799.t109 gnd 0.595595f
C6283 a_n8964_8799.t68 gnd 0.595595f
C6284 a_n8964_8799.n224 gnd 0.267255f
C6285 a_n8964_8799.t151 gnd 0.595595f
C6286 a_n8964_8799.t112 gnd 0.595595f
C6287 a_n8964_8799.t85 gnd 0.595595f
C6288 a_n8964_8799.n225 gnd 0.268145f
C6289 a_n8964_8799.t136 gnd 0.606868f
C6290 a_n8964_8799.n226 gnd 0.249678f
C6291 a_n8964_8799.t48 gnd 0.595595f
C6292 a_n8964_8799.n227 gnd 0.270437f
C6293 a_n8964_8799.n228 gnd 0.263929f
C6294 a_n8964_8799.n229 gnd 0.262653f
C6295 a_n8964_8799.n230 gnd 0.269811f
C6296 a_n8964_8799.n231 gnd 0.270066f
C6297 a_n8964_8799.n232 gnd 0.263291f
C6298 a_n8964_8799.n233 gnd 0.263291f
C6299 a_n8964_8799.n234 gnd 0.270066f
C6300 a_n8964_8799.n235 gnd 0.269811f
C6301 a_n8964_8799.n236 gnd 0.262653f
C6302 a_n8964_8799.n237 gnd 0.263929f
C6303 a_n8964_8799.n238 gnd 0.270437f
C6304 a_n8964_8799.t123 gnd 0.606858f
C6305 a_n8964_8799.t55 gnd 0.595595f
C6306 a_n8964_8799.t131 gnd 0.595595f
C6307 a_n8964_8799.n239 gnd 0.268145f
C6308 a_n8964_8799.t129 gnd 0.595595f
C6309 a_n8964_8799.t58 gnd 0.595595f
C6310 a_n8964_8799.t57 gnd 0.595595f
C6311 a_n8964_8799.n240 gnd 0.267255f
C6312 a_n8964_8799.t149 gnd 0.595595f
C6313 a_n8964_8799.t74 gnd 0.595595f
C6314 a_n8964_8799.t64 gnd 0.595595f
C6315 a_n8964_8799.n241 gnd 0.267686f
C6316 a_n8964_8799.t152 gnd 0.595595f
C6317 a_n8964_8799.t104 gnd 0.595595f
C6318 a_n8964_8799.t77 gnd 0.595595f
C6319 a_n8964_8799.n242 gnd 0.267686f
C6320 a_n8964_8799.t50 gnd 0.595595f
C6321 a_n8964_8799.t124 gnd 0.595595f
C6322 a_n8964_8799.t78 gnd 0.595595f
C6323 a_n8964_8799.n243 gnd 0.267255f
C6324 a_n8964_8799.t42 gnd 0.595595f
C6325 a_n8964_8799.t130 gnd 0.595595f
C6326 a_n8964_8799.t93 gnd 0.595595f
C6327 a_n8964_8799.n244 gnd 0.268145f
C6328 a_n8964_8799.t150 gnd 0.606868f
C6329 a_n8964_8799.n245 gnd 0.249678f
C6330 a_n8964_8799.t59 gnd 0.595595f
C6331 a_n8964_8799.n246 gnd 0.270437f
C6332 a_n8964_8799.n247 gnd 0.263929f
C6333 a_n8964_8799.n248 gnd 0.262653f
C6334 a_n8964_8799.n249 gnd 0.269811f
C6335 a_n8964_8799.n250 gnd 0.270066f
C6336 a_n8964_8799.n251 gnd 0.263291f
C6337 a_n8964_8799.n252 gnd 0.263291f
C6338 a_n8964_8799.n253 gnd 0.270066f
C6339 a_n8964_8799.n254 gnd 0.269811f
C6340 a_n8964_8799.n255 gnd 0.262653f
C6341 a_n8964_8799.n256 gnd 0.263929f
C6342 a_n8964_8799.n257 gnd 0.270437f
C6343 a_n8964_8799.n258 gnd 0.895395f
C6344 a_n8964_8799.t69 gnd 0.606858f
C6345 a_n8964_8799.t155 gnd 0.595595f
C6346 a_n8964_8799.t122 gnd 0.595595f
C6347 a_n8964_8799.n259 gnd 0.268145f
C6348 a_n8964_8799.t148 gnd 0.595595f
C6349 a_n8964_8799.t103 gnd 0.595595f
C6350 a_n8964_8799.t128 gnd 0.595595f
C6351 a_n8964_8799.n260 gnd 0.267255f
C6352 a_n8964_8799.t63 gnd 0.595595f
C6353 a_n8964_8799.t145 gnd 0.595595f
C6354 a_n8964_8799.t81 gnd 0.595595f
C6355 a_n8964_8799.n261 gnd 0.267686f
C6356 a_n8964_8799.t140 gnd 0.595595f
C6357 a_n8964_8799.t67 gnd 0.595595f
C6358 a_n8964_8799.t116 gnd 0.595595f
C6359 a_n8964_8799.n262 gnd 0.267686f
C6360 a_n8964_8799.t54 gnd 0.595595f
C6361 a_n8964_8799.t100 gnd 0.595595f
C6362 a_n8964_8799.t76 gnd 0.595595f
C6363 a_n8964_8799.n263 gnd 0.267255f
C6364 a_n8964_8799.t126 gnd 0.595595f
C6365 a_n8964_8799.t61 gnd 0.595595f
C6366 a_n8964_8799.t108 gnd 0.595595f
C6367 a_n8964_8799.n264 gnd 0.268145f
C6368 a_n8964_8799.t92 gnd 0.606868f
C6369 a_n8964_8799.n265 gnd 0.249678f
C6370 a_n8964_8799.t46 gnd 0.595595f
C6371 a_n8964_8799.n266 gnd 0.270437f
C6372 a_n8964_8799.n267 gnd 0.263929f
C6373 a_n8964_8799.n268 gnd 0.262653f
C6374 a_n8964_8799.n269 gnd 0.269811f
C6375 a_n8964_8799.n270 gnd 0.270066f
C6376 a_n8964_8799.n271 gnd 0.263291f
C6377 a_n8964_8799.n272 gnd 0.263291f
C6378 a_n8964_8799.n273 gnd 0.270066f
C6379 a_n8964_8799.n274 gnd 0.269811f
C6380 a_n8964_8799.n275 gnd 0.262653f
C6381 a_n8964_8799.n276 gnd 0.263929f
C6382 a_n8964_8799.n277 gnd 0.270437f
C6383 a_n8964_8799.n278 gnd 1.27195f
C6384 a_n8964_8799.n279 gnd 15.6153f
C6385 a_n8964_8799.n280 gnd 4.35889f
C6386 a_n8964_8799.n281 gnd 6.96179f
C6387 a_n8964_8799.t38 gnd 0.143639f
C6388 a_n8964_8799.t25 gnd 0.143639f
C6389 a_n8964_8799.n282 gnd 1.13104f
C6390 a_n8964_8799.t31 gnd 0.143639f
C6391 a_n8964_8799.t28 gnd 0.143639f
C6392 a_n8964_8799.n283 gnd 1.13104f
C6393 a_n8964_8799.t5 gnd 0.143639f
C6394 a_n8964_8799.t35 gnd 0.143639f
C6395 a_n8964_8799.n284 gnd 1.13104f
C6396 a_n8964_8799.t27 gnd 0.143639f
C6397 a_n8964_8799.t17 gnd 0.143639f
C6398 a_n8964_8799.n285 gnd 1.13104f
C6399 a_n8964_8799.n286 gnd 1.13291f
C6400 a_n8964_8799.t0 gnd 0.143639f
.ends

