* NGSPICE file created from opamp375.ext - technology: sky130A

.subckt opamp375 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd.t269 commonsourceibias.t48 CSoutput.t151 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 gnd.t134 gnd.t132 gnd.t133 gnd.t116 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X2 commonsourceibias.t47 commonsourceibias.t46 gnd.t268 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X3 a_n2804_13878.t7 a_n2982_13878.t64 vdd.t291 vdd.t290 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 a_n2804_13878.t31 a_n2982_13878.t21 a_n2982_13878.t22 vdd.t278 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 vdd.t68 a_n9628_8799.t40 CSoutput.t30 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 vdd.t23 CSoutput.t168 output.t16 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X7 a_n9628_8799.t1 plus.t5 a_n2903_n3924.t18 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X8 CSoutput.t31 a_n9628_8799.t41 vdd.t69 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 gnd.t267 commonsourceibias.t49 CSoutput.t150 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 gnd.t266 commonsourceibias.t8 commonsourceibias.t9 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 minus.t4 gnd.t129 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X12 vdd.t219 a_n9628_8799.t42 CSoutput.t88 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 gnd.t265 commonsourceibias.t50 CSoutput.t110 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 a_n2982_8322.t29 a_n2982_13878.t65 a_n9628_8799.t26 vdd.t288 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 CSoutput.t89 a_n9628_8799.t43 vdd.t220 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 vdd.t234 a_n9628_8799.t44 CSoutput.t102 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X17 CSoutput.t103 a_n9628_8799.t45 vdd.t235 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 vdd.t65 a_n9628_8799.t46 CSoutput.t28 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X19 vdd.t67 a_n9628_8799.t47 CSoutput.t29 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 CSoutput.t86 a_n9628_8799.t48 vdd.t217 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 a_n2982_13878.t7 minus.t5 a_n2903_n3924.t25 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X22 gnd.t264 commonsourceibias.t6 commonsourceibias.t7 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 a_n9628_8799.t15 plus.t6 a_n2903_n3924.t17 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X24 a_n9628_8799.t33 a_n2982_13878.t66 a_n2982_8322.t28 vdd.t274 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 a_n2982_13878.t11 minus.t6 a_n2903_n3924.t30 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 vdd.t218 a_n9628_8799.t49 CSoutput.t87 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X27 vdd.t232 a_n9628_8799.t50 CSoutput.t100 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 CSoutput.t101 a_n9628_8799.t51 vdd.t233 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 a_n9628_8799.t27 a_n2982_13878.t67 a_n2982_8322.t27 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X30 outputibias.t7 outputibias.t6 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X31 CSoutput.t109 commonsourceibias.t51 gnd.t263 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 gnd.t262 commonsourceibias.t4 commonsourceibias.t5 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 output.t15 CSoutput.t169 vdd.t16 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X34 a_n2903_n3924.t16 plus.t7 a_n9628_8799.t11 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X35 outputibias.t5 outputibias.t4 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X36 CSoutput.t108 commonsourceibias.t52 gnd.t261 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 CSoutput.t76 a_n9628_8799.t52 vdd.t206 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 a_n2903_n3924.t21 diffpairibias.t16 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X39 a_n2903_n3924.t29 minus.t7 a_n2982_13878.t10 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X40 CSoutput.t77 a_n9628_8799.t53 vdd.t208 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X41 vdd.t230 a_n9628_8799.t54 CSoutput.t98 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X42 vdd.t231 a_n9628_8799.t55 CSoutput.t99 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 CSoutput.t170 a_n2982_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X44 CSoutput.t107 commonsourceibias.t53 gnd.t260 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 vdd.t158 vdd.t156 vdd.t157 vdd.t147 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X46 outputibias.t3 outputibias.t2 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X47 vdd.t204 a_n9628_8799.t56 CSoutput.t74 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 a_n2804_13878.t30 a_n2982_13878.t19 a_n2982_13878.t20 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X49 CSoutput.t106 commonsourceibias.t54 gnd.t259 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X50 vdd.t155 vdd.t153 vdd.t154 vdd.t147 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X51 a_n2982_13878.t26 a_n2982_13878.t25 a_n2804_13878.t29 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X52 gnd.t128 gnd.t126 plus.t4 gnd.t127 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X53 CSoutput.t75 a_n9628_8799.t57 vdd.t205 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 gnd.t125 gnd.t122 gnd.t124 gnd.t123 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X55 vdd.t152 vdd.t150 vdd.t151 vdd.t129 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X56 a_n2903_n3924.t15 plus.t8 a_n9628_8799.t14 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X57 vdd.t81 a_n9628_8799.t58 CSoutput.t38 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X58 vdd.t82 a_n9628_8799.t59 CSoutput.t39 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 diffpairibias.t15 diffpairibias.t14 gnd.t271 gnd.t270 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X60 CSoutput.t96 a_n9628_8799.t60 vdd.t228 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 gnd.t121 gnd.t119 gnd.t120 gnd.t116 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X62 a_n2982_13878.t24 a_n2982_13878.t23 a_n2804_13878.t28 vdd.t273 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X63 CSoutput.t97 a_n9628_8799.t61 vdd.t229 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 vdd.t292 a_n9628_8799.t62 CSoutput.t152 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 a_n9628_8799.t29 a_n2982_13878.t68 a_n2982_8322.t26 vdd.t268 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X66 CSoutput.t153 a_n9628_8799.t63 vdd.t293 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 CSoutput.t171 a_n2982_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X68 a_n2982_13878.t18 a_n2982_13878.t17 a_n2804_13878.t27 vdd.t289 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X69 vdd.t294 a_n9628_8799.t64 CSoutput.t154 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 vdd.t295 a_n9628_8799.t65 CSoutput.t155 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 a_n9628_8799.t38 a_n2982_13878.t69 a_n2982_8322.t25 vdd.t266 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X72 CSoutput.t20 a_n9628_8799.t66 vdd.t53 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 gnd.t258 commonsourceibias.t55 CSoutput.t105 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 diffpairibias.t13 diffpairibias.t12 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X75 gnd.t257 commonsourceibias.t56 CSoutput.t104 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 CSoutput.t21 a_n9628_8799.t67 vdd.t55 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 commonsourceibias.t3 commonsourceibias.t2 gnd.t256 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 a_n9628_8799.t16 a_n2982_13878.t70 a_n2982_8322.t24 vdd.t281 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X79 gnd.t251 commonsourceibias.t57 CSoutput.t116 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 a_n2982_8322.t23 a_n2982_13878.t71 a_n9628_8799.t20 vdd.t289 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X81 CSoutput.t36 a_n9628_8799.t68 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 a_n2903_n3924.t23 minus.t8 a_n2982_13878.t5 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X83 a_n2903_n3924.t14 plus.t9 a_n9628_8799.t6 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X84 commonsourceibias.t1 commonsourceibias.t0 gnd.t255 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 gnd.t254 commonsourceibias.t58 CSoutput.t117 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 vdd.t149 vdd.t146 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X87 gnd.t253 commonsourceibias.t18 commonsourceibias.t19 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 a_n2903_n3924.t20 diffpairibias.t17 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X89 CSoutput.t37 a_n9628_8799.t69 vdd.t80 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 vdd.t226 a_n9628_8799.t70 CSoutput.t94 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X91 a_n2982_13878.t16 a_n2982_13878.t15 a_n2804_13878.t26 vdd.t288 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X92 vdd.t227 a_n9628_8799.t71 CSoutput.t95 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 a_n2903_n3924.t13 plus.t10 a_n9628_8799.t3 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X94 vdd.t224 a_n9628_8799.t72 CSoutput.t92 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 a_n9628_8799.t17 a_n2982_13878.t72 a_n2982_8322.t22 vdd.t277 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X96 a_n2982_13878.t58 a_n2982_13878.t57 a_n2804_13878.t25 vdd.t242 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X97 gnd.t252 commonsourceibias.t16 commonsourceibias.t17 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X98 commonsourceibias.t15 commonsourceibias.t14 gnd.t250 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 CSoutput.t115 commonsourceibias.t59 gnd.t249 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 output.t14 CSoutput.t172 vdd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X101 vdd.t225 a_n9628_8799.t73 CSoutput.t93 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X102 CSoutput.t72 a_n9628_8799.t74 vdd.t201 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 CSoutput.t73 a_n9628_8799.t75 vdd.t202 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X104 vdd.t145 vdd.t143 vdd.t144 vdd.t136 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X105 CSoutput.t114 commonsourceibias.t60 gnd.t248 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 CSoutput.t34 a_n9628_8799.t76 vdd.t74 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 vdd.t142 vdd.t139 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X108 gnd.t243 commonsourceibias.t61 CSoutput.t112 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X109 commonsourceibias.t13 commonsourceibias.t12 gnd.t247 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X110 gnd.t118 gnd.t115 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X111 CSoutput.t113 commonsourceibias.t62 gnd.t246 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X112 CSoutput.t35 a_n9628_8799.t77 vdd.t76 vdd.t75 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 a_n2804_13878.t24 a_n2982_13878.t55 a_n2982_13878.t56 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X114 vdd.t199 a_n9628_8799.t78 CSoutput.t70 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 vdd.t287 a_n2982_13878.t73 a_n2982_8322.t37 vdd.t286 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X116 a_n2982_13878.t62 a_n2982_13878.t61 a_n2804_13878.t23 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X117 gnd.t114 gnd.t112 minus.t3 gnd.t113 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X118 a_n2982_8322.t36 a_n2982_13878.t74 vdd.t285 vdd.t284 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X119 a_n2903_n3924.t31 diffpairibias.t18 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X120 CSoutput.t71 a_n9628_8799.t79 vdd.t200 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 commonsourceibias.t11 commonsourceibias.t10 gnd.t244 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 gnd.t111 gnd.t109 gnd.t110 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X123 vdd.t283 a_n2982_13878.t75 a_n2804_13878.t6 vdd.t282 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X124 vdd.t138 vdd.t135 vdd.t137 vdd.t136 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X125 a_n2804_13878.t22 a_n2982_13878.t59 a_n2982_13878.t60 vdd.t281 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 vdd.t71 a_n9628_8799.t80 CSoutput.t32 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X127 vdd.t73 a_n9628_8799.t81 CSoutput.t33 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 gnd.t242 commonsourceibias.t63 CSoutput.t111 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X129 a_n2982_8322.t21 a_n2982_13878.t76 a_n9628_8799.t37 vdd.t267 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 gnd.t241 commonsourceibias.t44 commonsourceibias.t45 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 a_n9628_8799.t7 plus.t11 a_n2903_n3924.t12 gnd.t142 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X132 vdd.t17 CSoutput.t173 output.t13 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X133 vdd.t134 vdd.t132 vdd.t133 vdd.t109 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X134 vdd.t131 vdd.t128 vdd.t130 vdd.t129 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X135 a_n2982_8322.t35 a_n2982_13878.t77 vdd.t280 vdd.t279 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X136 gnd.t239 commonsourceibias.t64 CSoutput.t149 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X137 output.t12 CSoutput.t174 vdd.t19 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X138 gnd.t238 commonsourceibias.t65 CSoutput.t148 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 a_n9628_8799.t39 a_n2982_13878.t78 a_n2982_8322.t20 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X140 a_n9628_8799.t2 plus.t12 a_n2903_n3924.t11 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X141 CSoutput.t90 a_n9628_8799.t82 vdd.t221 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 diffpairibias.t11 diffpairibias.t10 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X143 vdd.t223 a_n9628_8799.t83 CSoutput.t91 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X144 a_n2982_13878.t54 a_n2982_13878.t53 a_n2804_13878.t21 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X145 a_n9628_8799.t32 a_n2982_13878.t79 a_n2982_8322.t19 vdd.t278 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X146 CSoutput.t18 a_n9628_8799.t84 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X147 CSoutput.t19 a_n9628_8799.t85 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 gnd.t236 commonsourceibias.t66 CSoutput.t147 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 a_n2804_13878.t20 a_n2982_13878.t51 a_n2982_13878.t52 vdd.t277 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X150 gnd.t108 gnd.t106 gnd.t107 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X151 gnd.t235 commonsourceibias.t67 CSoutput.t146 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X152 vdd.t127 vdd.t125 vdd.t126 vdd.t88 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X153 CSoutput.t158 a_n9628_8799.t86 vdd.t298 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 vdd.t276 a_n2982_13878.t80 a_n2982_8322.t34 vdd.t275 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X155 CSoutput.t145 commonsourceibias.t68 gnd.t233 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 a_n2804_13878.t19 a_n2982_13878.t49 a_n2982_13878.t50 vdd.t274 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 vdd.t299 a_n9628_8799.t87 CSoutput.t159 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 vdd.t36 a_n9628_8799.t88 CSoutput.t10 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 a_n2982_13878.t8 minus.t9 a_n2903_n3924.t26 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X160 a_n2903_n3924.t10 plus.t13 a_n9628_8799.t0 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X161 a_n2982_13878.t48 a_n2982_13878.t47 a_n2804_13878.t18 vdd.t246 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 outputibias.t1 outputibias.t0 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X163 plus.t3 gnd.t103 gnd.t105 gnd.t104 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X164 vdd.t38 a_n9628_8799.t89 CSoutput.t11 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X165 vdd.t215 a_n9628_8799.t90 CSoutput.t84 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X166 CSoutput.t85 a_n9628_8799.t91 vdd.t216 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X167 a_n2903_n3924.t27 diffpairibias.t19 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X168 gnd.t102 gnd.t100 minus.t2 gnd.t101 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X169 gnd.t99 gnd.t96 gnd.t98 gnd.t97 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X170 vdd.t124 vdd.t122 vdd.t123 vdd.t96 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X171 a_n2903_n3924.t39 diffpairibias.t20 gnd.t281 gnd.t280 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X172 output.t11 CSoutput.t175 vdd.t8 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X173 a_n9628_8799.t13 plus.t14 a_n2903_n3924.t9 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X174 vdd.t5 a_n9628_8799.t92 CSoutput.t2 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 vdd.t15 CSoutput.t176 output.t10 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X176 CSoutput.t144 commonsourceibias.t69 gnd.t232 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 CSoutput.t143 commonsourceibias.t70 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 CSoutput.t3 a_n9628_8799.t93 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X179 vdd.t172 a_n9628_8799.t94 CSoutput.t48 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X180 gnd.t229 commonsourceibias.t71 CSoutput.t142 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X181 output.t0 outputibias.t8 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X182 vdd.t121 vdd.t119 vdd.t120 vdd.t109 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X183 CSoutput.t126 commonsourceibias.t72 gnd.t227 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 a_n9628_8799.t8 plus.t15 a_n2903_n3924.t8 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X185 a_n2804_13878.t17 a_n2982_13878.t45 a_n2982_13878.t46 vdd.t251 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X186 a_n2982_8322.t18 a_n2982_13878.t81 a_n9628_8799.t19 vdd.t273 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X187 CSoutput.t49 a_n9628_8799.t95 vdd.t173 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 CSoutput.t64 a_n9628_8799.t96 vdd.t192 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 output.t17 outputibias.t9 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X190 gnd.t95 gnd.t93 gnd.t94 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X191 CSoutput.t177 a_n2982_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X192 diffpairibias.t9 diffpairibias.t8 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X193 a_n2804_13878.t5 a_n2982_13878.t82 vdd.t272 vdd.t271 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X194 a_n2982_13878.t6 minus.t10 a_n2903_n3924.t24 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X195 vdd.t270 a_n2982_13878.t83 a_n2804_13878.t4 vdd.t269 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X196 CSoutput.t65 a_n9628_8799.t97 vdd.t194 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 CSoutput.t178 a_n2982_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X198 a_n2903_n3924.t7 plus.t16 a_n9628_8799.t10 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X199 vdd.t10 CSoutput.t179 output.t9 gnd.t14 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X200 vdd.t182 a_n9628_8799.t98 CSoutput.t56 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X201 vdd.t183 a_n9628_8799.t99 CSoutput.t57 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 vdd.t169 a_n9628_8799.t100 CSoutput.t46 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 gnd.t226 commonsourceibias.t73 CSoutput.t125 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 CSoutput.t124 commonsourceibias.t74 gnd.t225 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X205 CSoutput.t47 a_n9628_8799.t101 vdd.t171 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 a_n2804_13878.t16 a_n2982_13878.t43 a_n2982_13878.t44 vdd.t268 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 gnd.t224 commonsourceibias.t24 commonsourceibias.t25 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 gnd.t223 commonsourceibias.t75 CSoutput.t123 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X209 vdd.t60 a_n9628_8799.t102 CSoutput.t24 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X210 vdd.t61 a_n9628_8799.t103 CSoutput.t25 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 vdd.t18 CSoutput.t180 output.t8 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X212 CSoutput.t16 a_n9628_8799.t104 vdd.t46 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 output.t7 CSoutput.t181 vdd.t21 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X214 a_n2903_n3924.t32 minus.t11 a_n2982_13878.t12 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X215 gnd.t222 commonsourceibias.t76 CSoutput.t122 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 a_n2982_8322.t17 a_n2982_13878.t84 a_n9628_8799.t18 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X217 CSoutput.t17 a_n9628_8799.t105 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X218 a_n2982_13878.t34 a_n2982_13878.t33 a_n2804_13878.t15 vdd.t267 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X219 diffpairibias.t7 diffpairibias.t6 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X220 vdd.t32 a_n9628_8799.t106 CSoutput.t8 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X221 a_n2804_13878.t14 a_n2982_13878.t31 a_n2982_13878.t32 vdd.t266 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X222 vdd.t265 a_n2982_13878.t85 a_n2982_8322.t33 vdd.t264 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X223 gnd.t221 commonsourceibias.t22 commonsourceibias.t23 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X224 vdd.t34 a_n9628_8799.t107 CSoutput.t9 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 gnd.t92 gnd.t89 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X226 gnd.t88 gnd.t86 gnd.t87 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X227 gnd.t85 gnd.t83 gnd.t84 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X228 CSoutput.t121 commonsourceibias.t77 gnd.t219 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 plus.t2 gnd.t80 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X230 gnd.t79 gnd.t77 minus.t1 gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X231 CSoutput.t120 commonsourceibias.t78 gnd.t218 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X232 CSoutput.t164 a_n9628_8799.t108 vdd.t304 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 a_n2804_13878.t3 a_n2982_13878.t86 vdd.t263 vdd.t262 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X234 vdd.t305 a_n9628_8799.t109 CSoutput.t165 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 CSoutput.t62 a_n9628_8799.t110 vdd.t190 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X236 CSoutput.t63 a_n9628_8799.t111 vdd.t191 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 gnd.t217 commonsourceibias.t20 commonsourceibias.t21 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 gnd.t76 gnd.t73 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X239 vdd.t118 vdd.t116 vdd.t117 vdd.t92 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X240 vdd.t180 a_n9628_8799.t112 CSoutput.t54 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 a_n2903_n3924.t35 diffpairibias.t21 gnd.t273 gnd.t272 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X242 CSoutput.t119 commonsourceibias.t79 gnd.t216 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 vdd.t261 a_n2982_13878.t87 a_n2982_8322.t32 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X244 a_n2982_8322.t16 a_n2982_13878.t88 a_n9628_8799.t34 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X245 a_n9628_8799.t12 plus.t17 a_n2903_n3924.t6 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X246 a_n2982_13878.t1 minus.t12 a_n2903_n3924.t1 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X247 CSoutput.t118 commonsourceibias.t80 gnd.t215 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 a_n2903_n3924.t2 minus.t13 a_n2982_13878.t2 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X249 vdd.t181 a_n9628_8799.t113 CSoutput.t55 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 output.t6 CSoutput.t182 vdd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X251 vdd.t11 CSoutput.t183 output.t5 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X252 CSoutput.t134 commonsourceibias.t81 gnd.t214 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 gnd.t213 commonsourceibias.t82 CSoutput.t133 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 vdd.t115 vdd.t112 vdd.t114 vdd.t113 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X255 vdd.t166 a_n9628_8799.t114 CSoutput.t44 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 a_n2903_n3924.t28 minus.t14 a_n2982_13878.t9 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X257 gnd.t72 gnd.t70 gnd.t71 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X258 vdd.t168 a_n9628_8799.t115 CSoutput.t45 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X259 CSoutput.t0 a_n9628_8799.t116 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X260 vdd.t3 a_n9628_8799.t117 CSoutput.t1 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 CSoutput.t162 a_n9628_8799.t118 vdd.t302 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 a_n2903_n3924.t0 minus.t15 a_n2982_13878.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X263 a_n2804_13878.t13 a_n2982_13878.t37 a_n2982_13878.t38 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X264 CSoutput.t163 a_n9628_8799.t119 vdd.t303 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 CSoutput.t80 a_n9628_8799.t120 vdd.t211 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X266 gnd.t69 gnd.t67 gnd.t68 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X267 vdd.t22 CSoutput.t184 output.t4 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X268 a_n2982_8322.t15 a_n2982_13878.t89 a_n9628_8799.t21 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X269 diffpairibias.t5 diffpairibias.t4 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X270 CSoutput.t81 a_n9628_8799.t121 vdd.t212 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 CSoutput.t22 a_n9628_8799.t122 vdd.t57 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 vdd.t111 vdd.t108 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X273 gnd.t212 commonsourceibias.t83 CSoutput.t132 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 output.t19 outputibias.t10 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X275 CSoutput.t131 commonsourceibias.t84 gnd.t210 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X276 vdd.t59 a_n9628_8799.t123 CSoutput.t23 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 CSoutput.t185 a_n2982_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X278 a_n2982_8322.t31 a_n2982_13878.t90 vdd.t257 vdd.t256 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X279 output.t3 CSoutput.t186 vdd.t14 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X280 gnd.t209 commonsourceibias.t26 commonsourceibias.t27 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X281 gnd.t207 commonsourceibias.t85 CSoutput.t130 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 CSoutput.t160 a_n9628_8799.t124 vdd.t300 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 a_n2903_n3924.t19 minus.t16 a_n2982_13878.t3 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X284 vdd.t301 a_n9628_8799.t125 CSoutput.t161 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 CSoutput.t60 a_n9628_8799.t126 vdd.t188 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 vdd.t255 a_n2982_13878.t91 a_n2804_13878.t2 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X287 vdd.t189 a_n9628_8799.t127 CSoutput.t61 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 CSoutput.t6 a_n9628_8799.t128 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 output.t18 outputibias.t11 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X290 output.t2 CSoutput.t187 vdd.t9 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X291 gnd.t66 gnd.t63 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X292 vdd.t30 a_n9628_8799.t129 CSoutput.t7 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 CSoutput.t129 commonsourceibias.t86 gnd.t206 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 CSoutput.t128 commonsourceibias.t87 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 gnd.t62 gnd.t60 gnd.t61 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X296 gnd.t59 gnd.t56 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X297 gnd.t55 gnd.t53 plus.t1 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X298 a_n2982_8322.t14 a_n2982_13878.t92 a_n9628_8799.t31 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X299 a_n9628_8799.t30 a_n2982_13878.t93 a_n2982_8322.t13 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X300 a_n2804_13878.t1 a_n2982_13878.t94 vdd.t241 vdd.t240 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X301 vdd.t177 a_n9628_8799.t130 CSoutput.t52 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 vdd.t107 vdd.t105 vdd.t106 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X303 vdd.t104 vdd.t102 vdd.t103 vdd.t96 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X304 vdd.t178 a_n9628_8799.t131 CSoutput.t53 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 CSoutput.t42 a_n9628_8799.t132 vdd.t164 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 CSoutput.t43 a_n9628_8799.t133 vdd.t165 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X307 a_n2982_13878.t36 a_n2982_13878.t35 a_n2804_13878.t12 vdd.t243 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X308 CSoutput.t14 a_n9628_8799.t134 vdd.t42 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 a_n9628_8799.t22 a_n2982_13878.t95 a_n2982_8322.t12 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X310 a_n2903_n3924.t5 plus.t18 a_n9628_8799.t4 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X311 a_n2982_13878.t63 minus.t17 a_n2903_n3924.t37 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X312 a_n9628_8799.t35 a_n2982_13878.t96 a_n2982_8322.t11 vdd.t251 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X313 CSoutput.t127 commonsourceibias.t88 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 a_n2982_8322.t10 a_n2982_13878.t97 a_n9628_8799.t28 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X315 vdd.t44 a_n9628_8799.t135 CSoutput.t15 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 CSoutput.t78 a_n9628_8799.t136 vdd.t209 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 CSoutput.t79 a_n9628_8799.t137 vdd.t210 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X318 CSoutput.t4 a_n9628_8799.t138 vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 CSoutput.t5 a_n9628_8799.t139 vdd.t26 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 a_n2804_13878.t11 a_n2982_13878.t29 a_n2982_13878.t30 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X321 vdd.t296 a_n9628_8799.t140 CSoutput.t156 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 vdd.t297 a_n9628_8799.t141 CSoutput.t157 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 commonsourceibias.t33 commonsourceibias.t32 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 gnd.t199 commonsourceibias.t89 CSoutput.t139 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 vdd.t306 a_n9628_8799.t142 CSoutput.t166 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 gnd.t52 gnd.t49 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X327 gnd.t198 commonsourceibias.t90 CSoutput.t138 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 vdd.t13 CSoutput.t188 output.t1 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X329 a_n2903_n3924.t33 minus.t18 a_n2982_13878.t13 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X330 a_n2903_n3924.t36 diffpairibias.t22 gnd.t275 gnd.t274 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X331 vdd.t307 a_n9628_8799.t143 CSoutput.t167 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 gnd.t48 gnd.t45 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X333 gnd.t196 commonsourceibias.t91 CSoutput.t137 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 CSoutput.t82 a_n9628_8799.t144 vdd.t213 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 a_n2982_13878.t28 a_n2982_13878.t27 a_n2804_13878.t10 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X336 commonsourceibias.t31 commonsourceibias.t30 gnd.t194 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 a_n9628_8799.t24 a_n2982_13878.t98 a_n2982_8322.t9 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X338 vdd.t214 a_n9628_8799.t145 CSoutput.t83 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 CSoutput.t189 a_n2982_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X340 CSoutput.t68 a_n9628_8799.t146 vdd.t197 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 vdd.t101 vdd.t99 vdd.t100 vdd.t92 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X342 diffpairibias.t3 diffpairibias.t2 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X343 CSoutput.t69 a_n9628_8799.t147 vdd.t198 vdd.t75 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X344 gnd.t44 gnd.t42 plus.t0 gnd.t43 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X345 minus.t0 gnd.t39 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X346 gnd.t38 gnd.t35 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X347 a_n2982_8322.t8 a_n2982_13878.t99 a_n9628_8799.t25 vdd.t246 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X348 a_n2982_13878.t14 minus.t19 a_n2903_n3924.t34 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X349 commonsourceibias.t29 commonsourceibias.t28 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 vdd.t63 a_n9628_8799.t148 CSoutput.t26 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 vdd.t98 vdd.t95 vdd.t97 vdd.t96 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X352 gnd.t191 commonsourceibias.t92 CSoutput.t136 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 CSoutput.t27 a_n9628_8799.t149 vdd.t64 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 diffpairibias.t1 diffpairibias.t0 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X355 CSoutput.t12 a_n9628_8799.t150 vdd.t40 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X356 CSoutput.t135 commonsourceibias.t93 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 vdd.t245 a_n2982_13878.t100 a_n2804_13878.t0 vdd.t244 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X358 CSoutput.t13 a_n9628_8799.t151 vdd.t41 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 CSoutput.t58 a_n9628_8799.t152 vdd.t185 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X360 CSoutput.t141 commonsourceibias.t94 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X361 gnd.t34 gnd.t31 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X362 vdd.t187 a_n9628_8799.t153 CSoutput.t59 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 commonsourceibias.t43 commonsourceibias.t42 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 vdd.t175 a_n9628_8799.t154 CSoutput.t50 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X365 a_n9628_8799.t9 plus.t19 a_n2903_n3924.t4 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X366 a_n2982_8322.t7 a_n2982_13878.t101 a_n9628_8799.t23 vdd.t243 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X367 a_n2982_13878.t4 minus.t20 a_n2903_n3924.t22 gnd.t142 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X368 CSoutput.t140 commonsourceibias.t95 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 a_n2982_8322.t6 a_n2982_13878.t102 a_n9628_8799.t36 vdd.t242 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X370 gnd.t183 commonsourceibias.t40 commonsourceibias.t41 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 vdd.t176 a_n9628_8799.t155 CSoutput.t51 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 vdd.t160 a_n9628_8799.t156 CSoutput.t40 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X373 CSoutput.t41 a_n9628_8799.t157 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 commonsourceibias.t39 commonsourceibias.t38 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X375 vdd.t94 vdd.t91 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X376 a_n2982_8322.t30 a_n2982_13878.t103 vdd.t239 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X377 gnd.t30 gnd.t27 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X378 a_n2804_13878.t9 a_n2982_13878.t41 a_n2982_13878.t42 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X379 commonsourceibias.t37 commonsourceibias.t36 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X380 vdd.t90 vdd.t87 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X381 a_n2903_n3924.t3 plus.t20 a_n9628_8799.t5 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X382 a_n2903_n3924.t38 diffpairibias.t23 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X383 vdd.t86 vdd.t83 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X384 vdd.t195 a_n9628_8799.t158 CSoutput.t66 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X385 CSoutput.t67 a_n9628_8799.t159 vdd.t196 vdd.t75 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 gnd.t175 commonsourceibias.t34 commonsourceibias.t35 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 a_n2982_13878.t40 a_n2982_13878.t39 a_n2804_13878.t8 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 commonsourceibias.n25 commonsourceibias.t46 230.006
R1 commonsourceibias.n91 commonsourceibias.t62 230.006
R2 commonsourceibias.n154 commonsourceibias.t54 230.006
R3 commonsourceibias.n258 commonsourceibias.t26 230.006
R4 commonsourceibias.n217 commonsourceibias.t75 230.006
R5 commonsourceibias.n355 commonsourceibias.t64 230.006
R6 commonsourceibias.n70 commonsourceibias.t16 207.983
R7 commonsourceibias.n136 commonsourceibias.t71 207.983
R8 commonsourceibias.n199 commonsourceibias.t61 207.983
R9 commonsourceibias.n304 commonsourceibias.t36 207.983
R10 commonsourceibias.n338 commonsourceibias.t84 207.983
R11 commonsourceibias.n401 commonsourceibias.t74 207.983
R12 commonsourceibias.n10 commonsourceibias.t32 168.701
R13 commonsourceibias.n63 commonsourceibias.t44 168.701
R14 commonsourceibias.n57 commonsourceibias.t14 168.701
R15 commonsourceibias.n16 commonsourceibias.t22 168.701
R16 commonsourceibias.n49 commonsourceibias.t0 168.701
R17 commonsourceibias.n43 commonsourceibias.t8 168.701
R18 commonsourceibias.n19 commonsourceibias.t10 168.701
R19 commonsourceibias.n21 commonsourceibias.t18 168.701
R20 commonsourceibias.n23 commonsourceibias.t28 168.701
R21 commonsourceibias.n26 commonsourceibias.t4 168.701
R22 commonsourceibias.n1 commonsourceibias.t81 168.701
R23 commonsourceibias.n129 commonsourceibias.t55 168.701
R24 commonsourceibias.n123 commonsourceibias.t53 168.701
R25 commonsourceibias.n7 commonsourceibias.t76 168.701
R26 commonsourceibias.n115 commonsourceibias.t87 168.701
R27 commonsourceibias.n109 commonsourceibias.t50 168.701
R28 commonsourceibias.n85 commonsourceibias.t70 168.701
R29 commonsourceibias.n87 commonsourceibias.t67 168.701
R30 commonsourceibias.n89 commonsourceibias.t78 168.701
R31 commonsourceibias.n92 commonsourceibias.t65 168.701
R32 commonsourceibias.n155 commonsourceibias.t57 168.701
R33 commonsourceibias.n152 commonsourceibias.t68 168.701
R34 commonsourceibias.n150 commonsourceibias.t58 168.701
R35 commonsourceibias.n148 commonsourceibias.t60 168.701
R36 commonsourceibias.n172 commonsourceibias.t91 168.701
R37 commonsourceibias.n178 commonsourceibias.t77 168.701
R38 commonsourceibias.n145 commonsourceibias.t66 168.701
R39 commonsourceibias.n186 commonsourceibias.t95 168.701
R40 commonsourceibias.n192 commonsourceibias.t49 168.701
R41 commonsourceibias.n139 commonsourceibias.t72 168.701
R42 commonsourceibias.n259 commonsourceibias.t42 168.701
R43 commonsourceibias.n256 commonsourceibias.t20 168.701
R44 commonsourceibias.n254 commonsourceibias.t38 168.701
R45 commonsourceibias.n252 commonsourceibias.t6 168.701
R46 commonsourceibias.n276 commonsourceibias.t30 168.701
R47 commonsourceibias.n282 commonsourceibias.t40 168.701
R48 commonsourceibias.n284 commonsourceibias.t12 168.701
R49 commonsourceibias.n291 commonsourceibias.t34 168.701
R50 commonsourceibias.n297 commonsourceibias.t2 168.701
R51 commonsourceibias.n244 commonsourceibias.t24 168.701
R52 commonsourceibias.n203 commonsourceibias.t92 168.701
R53 commonsourceibias.n331 commonsourceibias.t51 168.701
R54 commonsourceibias.n325 commonsourceibias.t63 168.701
R55 commonsourceibias.n318 commonsourceibias.t88 168.701
R56 commonsourceibias.n316 commonsourceibias.t48 168.701
R57 commonsourceibias.n218 commonsourceibias.t59 168.701
R58 commonsourceibias.n215 commonsourceibias.t90 168.701
R59 commonsourceibias.n213 commonsourceibias.t80 168.701
R60 commonsourceibias.n211 commonsourceibias.t83 168.701
R61 commonsourceibias.n235 commonsourceibias.t94 168.701
R62 commonsourceibias.n356 commonsourceibias.t52 168.701
R63 commonsourceibias.n353 commonsourceibias.t82 168.701
R64 commonsourceibias.n351 commonsourceibias.t69 168.701
R65 commonsourceibias.n349 commonsourceibias.t73 168.701
R66 commonsourceibias.n373 commonsourceibias.t86 168.701
R67 commonsourceibias.n379 commonsourceibias.t89 168.701
R68 commonsourceibias.n381 commonsourceibias.t79 168.701
R69 commonsourceibias.n388 commonsourceibias.t56 168.701
R70 commonsourceibias.n394 commonsourceibias.t93 168.701
R71 commonsourceibias.n341 commonsourceibias.t85 168.701
R72 commonsourceibias.n27 commonsourceibias.n24 161.3
R73 commonsourceibias.n29 commonsourceibias.n28 161.3
R74 commonsourceibias.n31 commonsourceibias.n30 161.3
R75 commonsourceibias.n32 commonsourceibias.n22 161.3
R76 commonsourceibias.n34 commonsourceibias.n33 161.3
R77 commonsourceibias.n36 commonsourceibias.n35 161.3
R78 commonsourceibias.n37 commonsourceibias.n20 161.3
R79 commonsourceibias.n39 commonsourceibias.n38 161.3
R80 commonsourceibias.n41 commonsourceibias.n40 161.3
R81 commonsourceibias.n42 commonsourceibias.n18 161.3
R82 commonsourceibias.n45 commonsourceibias.n44 161.3
R83 commonsourceibias.n46 commonsourceibias.n17 161.3
R84 commonsourceibias.n48 commonsourceibias.n47 161.3
R85 commonsourceibias.n50 commonsourceibias.n15 161.3
R86 commonsourceibias.n52 commonsourceibias.n51 161.3
R87 commonsourceibias.n53 commonsourceibias.n14 161.3
R88 commonsourceibias.n55 commonsourceibias.n54 161.3
R89 commonsourceibias.n56 commonsourceibias.n13 161.3
R90 commonsourceibias.n59 commonsourceibias.n58 161.3
R91 commonsourceibias.n60 commonsourceibias.n12 161.3
R92 commonsourceibias.n62 commonsourceibias.n61 161.3
R93 commonsourceibias.n64 commonsourceibias.n11 161.3
R94 commonsourceibias.n66 commonsourceibias.n65 161.3
R95 commonsourceibias.n68 commonsourceibias.n67 161.3
R96 commonsourceibias.n69 commonsourceibias.n9 161.3
R97 commonsourceibias.n93 commonsourceibias.n90 161.3
R98 commonsourceibias.n95 commonsourceibias.n94 161.3
R99 commonsourceibias.n97 commonsourceibias.n96 161.3
R100 commonsourceibias.n98 commonsourceibias.n88 161.3
R101 commonsourceibias.n100 commonsourceibias.n99 161.3
R102 commonsourceibias.n102 commonsourceibias.n101 161.3
R103 commonsourceibias.n103 commonsourceibias.n86 161.3
R104 commonsourceibias.n105 commonsourceibias.n104 161.3
R105 commonsourceibias.n107 commonsourceibias.n106 161.3
R106 commonsourceibias.n108 commonsourceibias.n84 161.3
R107 commonsourceibias.n111 commonsourceibias.n110 161.3
R108 commonsourceibias.n112 commonsourceibias.n8 161.3
R109 commonsourceibias.n114 commonsourceibias.n113 161.3
R110 commonsourceibias.n116 commonsourceibias.n6 161.3
R111 commonsourceibias.n118 commonsourceibias.n117 161.3
R112 commonsourceibias.n119 commonsourceibias.n5 161.3
R113 commonsourceibias.n121 commonsourceibias.n120 161.3
R114 commonsourceibias.n122 commonsourceibias.n4 161.3
R115 commonsourceibias.n125 commonsourceibias.n124 161.3
R116 commonsourceibias.n126 commonsourceibias.n3 161.3
R117 commonsourceibias.n128 commonsourceibias.n127 161.3
R118 commonsourceibias.n130 commonsourceibias.n2 161.3
R119 commonsourceibias.n132 commonsourceibias.n131 161.3
R120 commonsourceibias.n134 commonsourceibias.n133 161.3
R121 commonsourceibias.n135 commonsourceibias.n0 161.3
R122 commonsourceibias.n198 commonsourceibias.n138 161.3
R123 commonsourceibias.n197 commonsourceibias.n196 161.3
R124 commonsourceibias.n195 commonsourceibias.n194 161.3
R125 commonsourceibias.n193 commonsourceibias.n140 161.3
R126 commonsourceibias.n191 commonsourceibias.n190 161.3
R127 commonsourceibias.n189 commonsourceibias.n141 161.3
R128 commonsourceibias.n188 commonsourceibias.n187 161.3
R129 commonsourceibias.n185 commonsourceibias.n142 161.3
R130 commonsourceibias.n184 commonsourceibias.n183 161.3
R131 commonsourceibias.n182 commonsourceibias.n143 161.3
R132 commonsourceibias.n181 commonsourceibias.n180 161.3
R133 commonsourceibias.n179 commonsourceibias.n144 161.3
R134 commonsourceibias.n177 commonsourceibias.n176 161.3
R135 commonsourceibias.n175 commonsourceibias.n146 161.3
R136 commonsourceibias.n174 commonsourceibias.n173 161.3
R137 commonsourceibias.n171 commonsourceibias.n147 161.3
R138 commonsourceibias.n170 commonsourceibias.n169 161.3
R139 commonsourceibias.n168 commonsourceibias.n167 161.3
R140 commonsourceibias.n166 commonsourceibias.n149 161.3
R141 commonsourceibias.n165 commonsourceibias.n164 161.3
R142 commonsourceibias.n163 commonsourceibias.n162 161.3
R143 commonsourceibias.n161 commonsourceibias.n151 161.3
R144 commonsourceibias.n160 commonsourceibias.n159 161.3
R145 commonsourceibias.n158 commonsourceibias.n157 161.3
R146 commonsourceibias.n156 commonsourceibias.n153 161.3
R147 commonsourceibias.n303 commonsourceibias.n243 161.3
R148 commonsourceibias.n302 commonsourceibias.n301 161.3
R149 commonsourceibias.n300 commonsourceibias.n299 161.3
R150 commonsourceibias.n298 commonsourceibias.n245 161.3
R151 commonsourceibias.n296 commonsourceibias.n295 161.3
R152 commonsourceibias.n294 commonsourceibias.n246 161.3
R153 commonsourceibias.n293 commonsourceibias.n292 161.3
R154 commonsourceibias.n290 commonsourceibias.n247 161.3
R155 commonsourceibias.n289 commonsourceibias.n288 161.3
R156 commonsourceibias.n287 commonsourceibias.n248 161.3
R157 commonsourceibias.n286 commonsourceibias.n285 161.3
R158 commonsourceibias.n283 commonsourceibias.n249 161.3
R159 commonsourceibias.n281 commonsourceibias.n280 161.3
R160 commonsourceibias.n279 commonsourceibias.n250 161.3
R161 commonsourceibias.n278 commonsourceibias.n277 161.3
R162 commonsourceibias.n275 commonsourceibias.n251 161.3
R163 commonsourceibias.n274 commonsourceibias.n273 161.3
R164 commonsourceibias.n272 commonsourceibias.n271 161.3
R165 commonsourceibias.n270 commonsourceibias.n253 161.3
R166 commonsourceibias.n269 commonsourceibias.n268 161.3
R167 commonsourceibias.n267 commonsourceibias.n266 161.3
R168 commonsourceibias.n265 commonsourceibias.n255 161.3
R169 commonsourceibias.n264 commonsourceibias.n263 161.3
R170 commonsourceibias.n262 commonsourceibias.n261 161.3
R171 commonsourceibias.n260 commonsourceibias.n257 161.3
R172 commonsourceibias.n237 commonsourceibias.n236 161.3
R173 commonsourceibias.n234 commonsourceibias.n210 161.3
R174 commonsourceibias.n233 commonsourceibias.n232 161.3
R175 commonsourceibias.n231 commonsourceibias.n230 161.3
R176 commonsourceibias.n229 commonsourceibias.n212 161.3
R177 commonsourceibias.n228 commonsourceibias.n227 161.3
R178 commonsourceibias.n226 commonsourceibias.n225 161.3
R179 commonsourceibias.n224 commonsourceibias.n214 161.3
R180 commonsourceibias.n223 commonsourceibias.n222 161.3
R181 commonsourceibias.n221 commonsourceibias.n220 161.3
R182 commonsourceibias.n219 commonsourceibias.n216 161.3
R183 commonsourceibias.n313 commonsourceibias.n209 161.3
R184 commonsourceibias.n337 commonsourceibias.n202 161.3
R185 commonsourceibias.n336 commonsourceibias.n335 161.3
R186 commonsourceibias.n334 commonsourceibias.n333 161.3
R187 commonsourceibias.n332 commonsourceibias.n204 161.3
R188 commonsourceibias.n330 commonsourceibias.n329 161.3
R189 commonsourceibias.n328 commonsourceibias.n205 161.3
R190 commonsourceibias.n327 commonsourceibias.n326 161.3
R191 commonsourceibias.n324 commonsourceibias.n206 161.3
R192 commonsourceibias.n323 commonsourceibias.n322 161.3
R193 commonsourceibias.n321 commonsourceibias.n207 161.3
R194 commonsourceibias.n320 commonsourceibias.n319 161.3
R195 commonsourceibias.n317 commonsourceibias.n208 161.3
R196 commonsourceibias.n315 commonsourceibias.n314 161.3
R197 commonsourceibias.n400 commonsourceibias.n340 161.3
R198 commonsourceibias.n399 commonsourceibias.n398 161.3
R199 commonsourceibias.n397 commonsourceibias.n396 161.3
R200 commonsourceibias.n395 commonsourceibias.n342 161.3
R201 commonsourceibias.n393 commonsourceibias.n392 161.3
R202 commonsourceibias.n391 commonsourceibias.n343 161.3
R203 commonsourceibias.n390 commonsourceibias.n389 161.3
R204 commonsourceibias.n387 commonsourceibias.n344 161.3
R205 commonsourceibias.n386 commonsourceibias.n385 161.3
R206 commonsourceibias.n384 commonsourceibias.n345 161.3
R207 commonsourceibias.n383 commonsourceibias.n382 161.3
R208 commonsourceibias.n380 commonsourceibias.n346 161.3
R209 commonsourceibias.n378 commonsourceibias.n377 161.3
R210 commonsourceibias.n376 commonsourceibias.n347 161.3
R211 commonsourceibias.n375 commonsourceibias.n374 161.3
R212 commonsourceibias.n372 commonsourceibias.n348 161.3
R213 commonsourceibias.n371 commonsourceibias.n370 161.3
R214 commonsourceibias.n369 commonsourceibias.n368 161.3
R215 commonsourceibias.n367 commonsourceibias.n350 161.3
R216 commonsourceibias.n366 commonsourceibias.n365 161.3
R217 commonsourceibias.n364 commonsourceibias.n363 161.3
R218 commonsourceibias.n362 commonsourceibias.n352 161.3
R219 commonsourceibias.n361 commonsourceibias.n360 161.3
R220 commonsourceibias.n359 commonsourceibias.n358 161.3
R221 commonsourceibias.n357 commonsourceibias.n354 161.3
R222 commonsourceibias.n80 commonsourceibias.n78 81.5057
R223 commonsourceibias.n240 commonsourceibias.n238 81.5057
R224 commonsourceibias.n80 commonsourceibias.n79 80.9324
R225 commonsourceibias.n82 commonsourceibias.n81 80.9324
R226 commonsourceibias.n77 commonsourceibias.n76 80.9324
R227 commonsourceibias.n75 commonsourceibias.n74 80.9324
R228 commonsourceibias.n73 commonsourceibias.n72 80.9324
R229 commonsourceibias.n307 commonsourceibias.n306 80.9324
R230 commonsourceibias.n309 commonsourceibias.n308 80.9324
R231 commonsourceibias.n311 commonsourceibias.n310 80.9324
R232 commonsourceibias.n242 commonsourceibias.n241 80.9324
R233 commonsourceibias.n240 commonsourceibias.n239 80.9324
R234 commonsourceibias.n71 commonsourceibias.n70 80.6037
R235 commonsourceibias.n137 commonsourceibias.n136 80.6037
R236 commonsourceibias.n200 commonsourceibias.n199 80.6037
R237 commonsourceibias.n305 commonsourceibias.n304 80.6037
R238 commonsourceibias.n339 commonsourceibias.n338 80.6037
R239 commonsourceibias.n402 commonsourceibias.n401 80.6037
R240 commonsourceibias.n65 commonsourceibias.n64 56.5617
R241 commonsourceibias.n51 commonsourceibias.n50 56.5617
R242 commonsourceibias.n42 commonsourceibias.n41 56.5617
R243 commonsourceibias.n28 commonsourceibias.n27 56.5617
R244 commonsourceibias.n131 commonsourceibias.n130 56.5617
R245 commonsourceibias.n117 commonsourceibias.n116 56.5617
R246 commonsourceibias.n108 commonsourceibias.n107 56.5617
R247 commonsourceibias.n94 commonsourceibias.n93 56.5617
R248 commonsourceibias.n157 commonsourceibias.n156 56.5617
R249 commonsourceibias.n171 commonsourceibias.n170 56.5617
R250 commonsourceibias.n180 commonsourceibias.n179 56.5617
R251 commonsourceibias.n194 commonsourceibias.n193 56.5617
R252 commonsourceibias.n261 commonsourceibias.n260 56.5617
R253 commonsourceibias.n275 commonsourceibias.n274 56.5617
R254 commonsourceibias.n285 commonsourceibias.n283 56.5617
R255 commonsourceibias.n299 commonsourceibias.n298 56.5617
R256 commonsourceibias.n333 commonsourceibias.n332 56.5617
R257 commonsourceibias.n319 commonsourceibias.n317 56.5617
R258 commonsourceibias.n220 commonsourceibias.n219 56.5617
R259 commonsourceibias.n234 commonsourceibias.n233 56.5617
R260 commonsourceibias.n358 commonsourceibias.n357 56.5617
R261 commonsourceibias.n372 commonsourceibias.n371 56.5617
R262 commonsourceibias.n382 commonsourceibias.n380 56.5617
R263 commonsourceibias.n396 commonsourceibias.n395 56.5617
R264 commonsourceibias.n56 commonsourceibias.n55 56.0773
R265 commonsourceibias.n37 commonsourceibias.n36 56.0773
R266 commonsourceibias.n122 commonsourceibias.n121 56.0773
R267 commonsourceibias.n103 commonsourceibias.n102 56.0773
R268 commonsourceibias.n166 commonsourceibias.n165 56.0773
R269 commonsourceibias.n185 commonsourceibias.n184 56.0773
R270 commonsourceibias.n270 commonsourceibias.n269 56.0773
R271 commonsourceibias.n290 commonsourceibias.n289 56.0773
R272 commonsourceibias.n324 commonsourceibias.n323 56.0773
R273 commonsourceibias.n229 commonsourceibias.n228 56.0773
R274 commonsourceibias.n367 commonsourceibias.n366 56.0773
R275 commonsourceibias.n387 commonsourceibias.n386 56.0773
R276 commonsourceibias.n70 commonsourceibias.n69 46.0096
R277 commonsourceibias.n136 commonsourceibias.n135 46.0096
R278 commonsourceibias.n199 commonsourceibias.n198 46.0096
R279 commonsourceibias.n304 commonsourceibias.n303 46.0096
R280 commonsourceibias.n338 commonsourceibias.n337 46.0096
R281 commonsourceibias.n401 commonsourceibias.n400 46.0096
R282 commonsourceibias.n58 commonsourceibias.n12 41.5458
R283 commonsourceibias.n33 commonsourceibias.n32 41.5458
R284 commonsourceibias.n124 commonsourceibias.n3 41.5458
R285 commonsourceibias.n99 commonsourceibias.n98 41.5458
R286 commonsourceibias.n162 commonsourceibias.n161 41.5458
R287 commonsourceibias.n187 commonsourceibias.n141 41.5458
R288 commonsourceibias.n266 commonsourceibias.n265 41.5458
R289 commonsourceibias.n292 commonsourceibias.n246 41.5458
R290 commonsourceibias.n326 commonsourceibias.n205 41.5458
R291 commonsourceibias.n225 commonsourceibias.n224 41.5458
R292 commonsourceibias.n363 commonsourceibias.n362 41.5458
R293 commonsourceibias.n389 commonsourceibias.n343 41.5458
R294 commonsourceibias.n48 commonsourceibias.n17 40.577
R295 commonsourceibias.n44 commonsourceibias.n17 40.577
R296 commonsourceibias.n114 commonsourceibias.n8 40.577
R297 commonsourceibias.n110 commonsourceibias.n8 40.577
R298 commonsourceibias.n173 commonsourceibias.n146 40.577
R299 commonsourceibias.n177 commonsourceibias.n146 40.577
R300 commonsourceibias.n277 commonsourceibias.n250 40.577
R301 commonsourceibias.n281 commonsourceibias.n250 40.577
R302 commonsourceibias.n315 commonsourceibias.n209 40.577
R303 commonsourceibias.n236 commonsourceibias.n209 40.577
R304 commonsourceibias.n374 commonsourceibias.n347 40.577
R305 commonsourceibias.n378 commonsourceibias.n347 40.577
R306 commonsourceibias.n62 commonsourceibias.n12 39.6083
R307 commonsourceibias.n32 commonsourceibias.n31 39.6083
R308 commonsourceibias.n128 commonsourceibias.n3 39.6083
R309 commonsourceibias.n98 commonsourceibias.n97 39.6083
R310 commonsourceibias.n161 commonsourceibias.n160 39.6083
R311 commonsourceibias.n191 commonsourceibias.n141 39.6083
R312 commonsourceibias.n265 commonsourceibias.n264 39.6083
R313 commonsourceibias.n296 commonsourceibias.n246 39.6083
R314 commonsourceibias.n330 commonsourceibias.n205 39.6083
R315 commonsourceibias.n224 commonsourceibias.n223 39.6083
R316 commonsourceibias.n362 commonsourceibias.n361 39.6083
R317 commonsourceibias.n393 commonsourceibias.n343 39.6083
R318 commonsourceibias.n26 commonsourceibias.n25 33.0515
R319 commonsourceibias.n92 commonsourceibias.n91 33.0515
R320 commonsourceibias.n155 commonsourceibias.n154 33.0515
R321 commonsourceibias.n259 commonsourceibias.n258 33.0515
R322 commonsourceibias.n218 commonsourceibias.n217 33.0515
R323 commonsourceibias.n356 commonsourceibias.n355 33.0515
R324 commonsourceibias.n25 commonsourceibias.n24 28.5514
R325 commonsourceibias.n91 commonsourceibias.n90 28.5514
R326 commonsourceibias.n154 commonsourceibias.n153 28.5514
R327 commonsourceibias.n258 commonsourceibias.n257 28.5514
R328 commonsourceibias.n217 commonsourceibias.n216 28.5514
R329 commonsourceibias.n355 commonsourceibias.n354 28.5514
R330 commonsourceibias.n69 commonsourceibias.n68 26.0455
R331 commonsourceibias.n135 commonsourceibias.n134 26.0455
R332 commonsourceibias.n198 commonsourceibias.n197 26.0455
R333 commonsourceibias.n303 commonsourceibias.n302 26.0455
R334 commonsourceibias.n337 commonsourceibias.n336 26.0455
R335 commonsourceibias.n400 commonsourceibias.n399 26.0455
R336 commonsourceibias.n55 commonsourceibias.n14 25.0767
R337 commonsourceibias.n38 commonsourceibias.n37 25.0767
R338 commonsourceibias.n121 commonsourceibias.n5 25.0767
R339 commonsourceibias.n104 commonsourceibias.n103 25.0767
R340 commonsourceibias.n167 commonsourceibias.n166 25.0767
R341 commonsourceibias.n184 commonsourceibias.n143 25.0767
R342 commonsourceibias.n271 commonsourceibias.n270 25.0767
R343 commonsourceibias.n289 commonsourceibias.n248 25.0767
R344 commonsourceibias.n323 commonsourceibias.n207 25.0767
R345 commonsourceibias.n230 commonsourceibias.n229 25.0767
R346 commonsourceibias.n368 commonsourceibias.n367 25.0767
R347 commonsourceibias.n386 commonsourceibias.n345 25.0767
R348 commonsourceibias.n51 commonsourceibias.n16 24.3464
R349 commonsourceibias.n41 commonsourceibias.n19 24.3464
R350 commonsourceibias.n117 commonsourceibias.n7 24.3464
R351 commonsourceibias.n107 commonsourceibias.n85 24.3464
R352 commonsourceibias.n170 commonsourceibias.n148 24.3464
R353 commonsourceibias.n180 commonsourceibias.n145 24.3464
R354 commonsourceibias.n274 commonsourceibias.n252 24.3464
R355 commonsourceibias.n285 commonsourceibias.n284 24.3464
R356 commonsourceibias.n319 commonsourceibias.n318 24.3464
R357 commonsourceibias.n233 commonsourceibias.n211 24.3464
R358 commonsourceibias.n371 commonsourceibias.n349 24.3464
R359 commonsourceibias.n382 commonsourceibias.n381 24.3464
R360 commonsourceibias.n65 commonsourceibias.n10 23.8546
R361 commonsourceibias.n27 commonsourceibias.n26 23.8546
R362 commonsourceibias.n131 commonsourceibias.n1 23.8546
R363 commonsourceibias.n93 commonsourceibias.n92 23.8546
R364 commonsourceibias.n156 commonsourceibias.n155 23.8546
R365 commonsourceibias.n194 commonsourceibias.n139 23.8546
R366 commonsourceibias.n260 commonsourceibias.n259 23.8546
R367 commonsourceibias.n299 commonsourceibias.n244 23.8546
R368 commonsourceibias.n333 commonsourceibias.n203 23.8546
R369 commonsourceibias.n219 commonsourceibias.n218 23.8546
R370 commonsourceibias.n357 commonsourceibias.n356 23.8546
R371 commonsourceibias.n396 commonsourceibias.n341 23.8546
R372 commonsourceibias.n64 commonsourceibias.n63 16.9689
R373 commonsourceibias.n28 commonsourceibias.n23 16.9689
R374 commonsourceibias.n130 commonsourceibias.n129 16.9689
R375 commonsourceibias.n94 commonsourceibias.n89 16.9689
R376 commonsourceibias.n157 commonsourceibias.n152 16.9689
R377 commonsourceibias.n193 commonsourceibias.n192 16.9689
R378 commonsourceibias.n261 commonsourceibias.n256 16.9689
R379 commonsourceibias.n298 commonsourceibias.n297 16.9689
R380 commonsourceibias.n332 commonsourceibias.n331 16.9689
R381 commonsourceibias.n220 commonsourceibias.n215 16.9689
R382 commonsourceibias.n358 commonsourceibias.n353 16.9689
R383 commonsourceibias.n395 commonsourceibias.n394 16.9689
R384 commonsourceibias.n50 commonsourceibias.n49 16.477
R385 commonsourceibias.n43 commonsourceibias.n42 16.477
R386 commonsourceibias.n116 commonsourceibias.n115 16.477
R387 commonsourceibias.n109 commonsourceibias.n108 16.477
R388 commonsourceibias.n172 commonsourceibias.n171 16.477
R389 commonsourceibias.n179 commonsourceibias.n178 16.477
R390 commonsourceibias.n276 commonsourceibias.n275 16.477
R391 commonsourceibias.n283 commonsourceibias.n282 16.477
R392 commonsourceibias.n317 commonsourceibias.n316 16.477
R393 commonsourceibias.n235 commonsourceibias.n234 16.477
R394 commonsourceibias.n373 commonsourceibias.n372 16.477
R395 commonsourceibias.n380 commonsourceibias.n379 16.477
R396 commonsourceibias.n57 commonsourceibias.n56 15.9852
R397 commonsourceibias.n36 commonsourceibias.n21 15.9852
R398 commonsourceibias.n123 commonsourceibias.n122 15.9852
R399 commonsourceibias.n102 commonsourceibias.n87 15.9852
R400 commonsourceibias.n165 commonsourceibias.n150 15.9852
R401 commonsourceibias.n186 commonsourceibias.n185 15.9852
R402 commonsourceibias.n269 commonsourceibias.n254 15.9852
R403 commonsourceibias.n291 commonsourceibias.n290 15.9852
R404 commonsourceibias.n325 commonsourceibias.n324 15.9852
R405 commonsourceibias.n228 commonsourceibias.n213 15.9852
R406 commonsourceibias.n366 commonsourceibias.n351 15.9852
R407 commonsourceibias.n388 commonsourceibias.n387 15.9852
R408 commonsourceibias.n73 commonsourceibias.n71 13.2057
R409 commonsourceibias.n307 commonsourceibias.n305 13.2057
R410 commonsourceibias.n404 commonsourceibias.n201 11.9876
R411 commonsourceibias.n404 commonsourceibias.n403 10.3347
R412 commonsourceibias.n112 commonsourceibias.n83 9.50363
R413 commonsourceibias.n313 commonsourceibias.n312 9.50363
R414 commonsourceibias.n201 commonsourceibias.n137 8.732
R415 commonsourceibias.n403 commonsourceibias.n339 8.732
R416 commonsourceibias.n58 commonsourceibias.n57 8.60764
R417 commonsourceibias.n33 commonsourceibias.n21 8.60764
R418 commonsourceibias.n124 commonsourceibias.n123 8.60764
R419 commonsourceibias.n99 commonsourceibias.n87 8.60764
R420 commonsourceibias.n162 commonsourceibias.n150 8.60764
R421 commonsourceibias.n187 commonsourceibias.n186 8.60764
R422 commonsourceibias.n266 commonsourceibias.n254 8.60764
R423 commonsourceibias.n292 commonsourceibias.n291 8.60764
R424 commonsourceibias.n326 commonsourceibias.n325 8.60764
R425 commonsourceibias.n225 commonsourceibias.n213 8.60764
R426 commonsourceibias.n363 commonsourceibias.n351 8.60764
R427 commonsourceibias.n389 commonsourceibias.n388 8.60764
R428 commonsourceibias.n49 commonsourceibias.n48 8.11581
R429 commonsourceibias.n44 commonsourceibias.n43 8.11581
R430 commonsourceibias.n115 commonsourceibias.n114 8.11581
R431 commonsourceibias.n110 commonsourceibias.n109 8.11581
R432 commonsourceibias.n173 commonsourceibias.n172 8.11581
R433 commonsourceibias.n178 commonsourceibias.n177 8.11581
R434 commonsourceibias.n277 commonsourceibias.n276 8.11581
R435 commonsourceibias.n282 commonsourceibias.n281 8.11581
R436 commonsourceibias.n316 commonsourceibias.n315 8.11581
R437 commonsourceibias.n236 commonsourceibias.n235 8.11581
R438 commonsourceibias.n374 commonsourceibias.n373 8.11581
R439 commonsourceibias.n379 commonsourceibias.n378 8.11581
R440 commonsourceibias.n63 commonsourceibias.n62 7.62397
R441 commonsourceibias.n31 commonsourceibias.n23 7.62397
R442 commonsourceibias.n129 commonsourceibias.n128 7.62397
R443 commonsourceibias.n97 commonsourceibias.n89 7.62397
R444 commonsourceibias.n160 commonsourceibias.n152 7.62397
R445 commonsourceibias.n192 commonsourceibias.n191 7.62397
R446 commonsourceibias.n264 commonsourceibias.n256 7.62397
R447 commonsourceibias.n297 commonsourceibias.n296 7.62397
R448 commonsourceibias.n331 commonsourceibias.n330 7.62397
R449 commonsourceibias.n223 commonsourceibias.n215 7.62397
R450 commonsourceibias.n361 commonsourceibias.n353 7.62397
R451 commonsourceibias.n394 commonsourceibias.n393 7.62397
R452 commonsourceibias.n201 commonsourceibias.n200 5.00473
R453 commonsourceibias.n403 commonsourceibias.n402 5.00473
R454 commonsourceibias commonsourceibias.n404 4.08303
R455 commonsourceibias.n78 commonsourceibias.t5 2.82907
R456 commonsourceibias.n78 commonsourceibias.t47 2.82907
R457 commonsourceibias.n79 commonsourceibias.t19 2.82907
R458 commonsourceibias.n79 commonsourceibias.t29 2.82907
R459 commonsourceibias.n81 commonsourceibias.t9 2.82907
R460 commonsourceibias.n81 commonsourceibias.t11 2.82907
R461 commonsourceibias.n76 commonsourceibias.t23 2.82907
R462 commonsourceibias.n76 commonsourceibias.t1 2.82907
R463 commonsourceibias.n74 commonsourceibias.t45 2.82907
R464 commonsourceibias.n74 commonsourceibias.t15 2.82907
R465 commonsourceibias.n72 commonsourceibias.t17 2.82907
R466 commonsourceibias.n72 commonsourceibias.t33 2.82907
R467 commonsourceibias.n306 commonsourceibias.t25 2.82907
R468 commonsourceibias.n306 commonsourceibias.t37 2.82907
R469 commonsourceibias.n308 commonsourceibias.t35 2.82907
R470 commonsourceibias.n308 commonsourceibias.t3 2.82907
R471 commonsourceibias.n310 commonsourceibias.t41 2.82907
R472 commonsourceibias.n310 commonsourceibias.t13 2.82907
R473 commonsourceibias.n241 commonsourceibias.t7 2.82907
R474 commonsourceibias.n241 commonsourceibias.t31 2.82907
R475 commonsourceibias.n239 commonsourceibias.t21 2.82907
R476 commonsourceibias.n239 commonsourceibias.t39 2.82907
R477 commonsourceibias.n238 commonsourceibias.t27 2.82907
R478 commonsourceibias.n238 commonsourceibias.t43 2.82907
R479 commonsourceibias.n68 commonsourceibias.n10 0.738255
R480 commonsourceibias.n134 commonsourceibias.n1 0.738255
R481 commonsourceibias.n197 commonsourceibias.n139 0.738255
R482 commonsourceibias.n302 commonsourceibias.n244 0.738255
R483 commonsourceibias.n336 commonsourceibias.n203 0.738255
R484 commonsourceibias.n399 commonsourceibias.n341 0.738255
R485 commonsourceibias.n75 commonsourceibias.n73 0.573776
R486 commonsourceibias.n77 commonsourceibias.n75 0.573776
R487 commonsourceibias.n82 commonsourceibias.n80 0.573776
R488 commonsourceibias.n242 commonsourceibias.n240 0.573776
R489 commonsourceibias.n311 commonsourceibias.n309 0.573776
R490 commonsourceibias.n309 commonsourceibias.n307 0.573776
R491 commonsourceibias.n83 commonsourceibias.n77 0.287138
R492 commonsourceibias.n83 commonsourceibias.n82 0.287138
R493 commonsourceibias.n312 commonsourceibias.n242 0.287138
R494 commonsourceibias.n312 commonsourceibias.n311 0.287138
R495 commonsourceibias.n71 commonsourceibias.n9 0.285035
R496 commonsourceibias.n137 commonsourceibias.n0 0.285035
R497 commonsourceibias.n200 commonsourceibias.n138 0.285035
R498 commonsourceibias.n305 commonsourceibias.n243 0.285035
R499 commonsourceibias.n339 commonsourceibias.n202 0.285035
R500 commonsourceibias.n402 commonsourceibias.n340 0.285035
R501 commonsourceibias.n16 commonsourceibias.n14 0.246418
R502 commonsourceibias.n38 commonsourceibias.n19 0.246418
R503 commonsourceibias.n7 commonsourceibias.n5 0.246418
R504 commonsourceibias.n104 commonsourceibias.n85 0.246418
R505 commonsourceibias.n167 commonsourceibias.n148 0.246418
R506 commonsourceibias.n145 commonsourceibias.n143 0.246418
R507 commonsourceibias.n271 commonsourceibias.n252 0.246418
R508 commonsourceibias.n284 commonsourceibias.n248 0.246418
R509 commonsourceibias.n318 commonsourceibias.n207 0.246418
R510 commonsourceibias.n230 commonsourceibias.n211 0.246418
R511 commonsourceibias.n368 commonsourceibias.n349 0.246418
R512 commonsourceibias.n381 commonsourceibias.n345 0.246418
R513 commonsourceibias.n67 commonsourceibias.n9 0.189894
R514 commonsourceibias.n67 commonsourceibias.n66 0.189894
R515 commonsourceibias.n66 commonsourceibias.n11 0.189894
R516 commonsourceibias.n61 commonsourceibias.n11 0.189894
R517 commonsourceibias.n61 commonsourceibias.n60 0.189894
R518 commonsourceibias.n60 commonsourceibias.n59 0.189894
R519 commonsourceibias.n59 commonsourceibias.n13 0.189894
R520 commonsourceibias.n54 commonsourceibias.n13 0.189894
R521 commonsourceibias.n54 commonsourceibias.n53 0.189894
R522 commonsourceibias.n53 commonsourceibias.n52 0.189894
R523 commonsourceibias.n52 commonsourceibias.n15 0.189894
R524 commonsourceibias.n47 commonsourceibias.n15 0.189894
R525 commonsourceibias.n47 commonsourceibias.n46 0.189894
R526 commonsourceibias.n46 commonsourceibias.n45 0.189894
R527 commonsourceibias.n45 commonsourceibias.n18 0.189894
R528 commonsourceibias.n40 commonsourceibias.n18 0.189894
R529 commonsourceibias.n40 commonsourceibias.n39 0.189894
R530 commonsourceibias.n39 commonsourceibias.n20 0.189894
R531 commonsourceibias.n35 commonsourceibias.n20 0.189894
R532 commonsourceibias.n35 commonsourceibias.n34 0.189894
R533 commonsourceibias.n34 commonsourceibias.n22 0.189894
R534 commonsourceibias.n30 commonsourceibias.n22 0.189894
R535 commonsourceibias.n30 commonsourceibias.n29 0.189894
R536 commonsourceibias.n29 commonsourceibias.n24 0.189894
R537 commonsourceibias.n111 commonsourceibias.n84 0.189894
R538 commonsourceibias.n106 commonsourceibias.n84 0.189894
R539 commonsourceibias.n106 commonsourceibias.n105 0.189894
R540 commonsourceibias.n105 commonsourceibias.n86 0.189894
R541 commonsourceibias.n101 commonsourceibias.n86 0.189894
R542 commonsourceibias.n101 commonsourceibias.n100 0.189894
R543 commonsourceibias.n100 commonsourceibias.n88 0.189894
R544 commonsourceibias.n96 commonsourceibias.n88 0.189894
R545 commonsourceibias.n96 commonsourceibias.n95 0.189894
R546 commonsourceibias.n95 commonsourceibias.n90 0.189894
R547 commonsourceibias.n133 commonsourceibias.n0 0.189894
R548 commonsourceibias.n133 commonsourceibias.n132 0.189894
R549 commonsourceibias.n132 commonsourceibias.n2 0.189894
R550 commonsourceibias.n127 commonsourceibias.n2 0.189894
R551 commonsourceibias.n127 commonsourceibias.n126 0.189894
R552 commonsourceibias.n126 commonsourceibias.n125 0.189894
R553 commonsourceibias.n125 commonsourceibias.n4 0.189894
R554 commonsourceibias.n120 commonsourceibias.n4 0.189894
R555 commonsourceibias.n120 commonsourceibias.n119 0.189894
R556 commonsourceibias.n119 commonsourceibias.n118 0.189894
R557 commonsourceibias.n118 commonsourceibias.n6 0.189894
R558 commonsourceibias.n113 commonsourceibias.n6 0.189894
R559 commonsourceibias.n196 commonsourceibias.n138 0.189894
R560 commonsourceibias.n196 commonsourceibias.n195 0.189894
R561 commonsourceibias.n195 commonsourceibias.n140 0.189894
R562 commonsourceibias.n190 commonsourceibias.n140 0.189894
R563 commonsourceibias.n190 commonsourceibias.n189 0.189894
R564 commonsourceibias.n189 commonsourceibias.n188 0.189894
R565 commonsourceibias.n188 commonsourceibias.n142 0.189894
R566 commonsourceibias.n183 commonsourceibias.n142 0.189894
R567 commonsourceibias.n183 commonsourceibias.n182 0.189894
R568 commonsourceibias.n182 commonsourceibias.n181 0.189894
R569 commonsourceibias.n181 commonsourceibias.n144 0.189894
R570 commonsourceibias.n176 commonsourceibias.n144 0.189894
R571 commonsourceibias.n176 commonsourceibias.n175 0.189894
R572 commonsourceibias.n175 commonsourceibias.n174 0.189894
R573 commonsourceibias.n174 commonsourceibias.n147 0.189894
R574 commonsourceibias.n169 commonsourceibias.n147 0.189894
R575 commonsourceibias.n169 commonsourceibias.n168 0.189894
R576 commonsourceibias.n168 commonsourceibias.n149 0.189894
R577 commonsourceibias.n164 commonsourceibias.n149 0.189894
R578 commonsourceibias.n164 commonsourceibias.n163 0.189894
R579 commonsourceibias.n163 commonsourceibias.n151 0.189894
R580 commonsourceibias.n159 commonsourceibias.n151 0.189894
R581 commonsourceibias.n159 commonsourceibias.n158 0.189894
R582 commonsourceibias.n158 commonsourceibias.n153 0.189894
R583 commonsourceibias.n262 commonsourceibias.n257 0.189894
R584 commonsourceibias.n263 commonsourceibias.n262 0.189894
R585 commonsourceibias.n263 commonsourceibias.n255 0.189894
R586 commonsourceibias.n267 commonsourceibias.n255 0.189894
R587 commonsourceibias.n268 commonsourceibias.n267 0.189894
R588 commonsourceibias.n268 commonsourceibias.n253 0.189894
R589 commonsourceibias.n272 commonsourceibias.n253 0.189894
R590 commonsourceibias.n273 commonsourceibias.n272 0.189894
R591 commonsourceibias.n273 commonsourceibias.n251 0.189894
R592 commonsourceibias.n278 commonsourceibias.n251 0.189894
R593 commonsourceibias.n279 commonsourceibias.n278 0.189894
R594 commonsourceibias.n280 commonsourceibias.n279 0.189894
R595 commonsourceibias.n280 commonsourceibias.n249 0.189894
R596 commonsourceibias.n286 commonsourceibias.n249 0.189894
R597 commonsourceibias.n287 commonsourceibias.n286 0.189894
R598 commonsourceibias.n288 commonsourceibias.n287 0.189894
R599 commonsourceibias.n288 commonsourceibias.n247 0.189894
R600 commonsourceibias.n293 commonsourceibias.n247 0.189894
R601 commonsourceibias.n294 commonsourceibias.n293 0.189894
R602 commonsourceibias.n295 commonsourceibias.n294 0.189894
R603 commonsourceibias.n295 commonsourceibias.n245 0.189894
R604 commonsourceibias.n300 commonsourceibias.n245 0.189894
R605 commonsourceibias.n301 commonsourceibias.n300 0.189894
R606 commonsourceibias.n301 commonsourceibias.n243 0.189894
R607 commonsourceibias.n221 commonsourceibias.n216 0.189894
R608 commonsourceibias.n222 commonsourceibias.n221 0.189894
R609 commonsourceibias.n222 commonsourceibias.n214 0.189894
R610 commonsourceibias.n226 commonsourceibias.n214 0.189894
R611 commonsourceibias.n227 commonsourceibias.n226 0.189894
R612 commonsourceibias.n227 commonsourceibias.n212 0.189894
R613 commonsourceibias.n231 commonsourceibias.n212 0.189894
R614 commonsourceibias.n232 commonsourceibias.n231 0.189894
R615 commonsourceibias.n232 commonsourceibias.n210 0.189894
R616 commonsourceibias.n237 commonsourceibias.n210 0.189894
R617 commonsourceibias.n314 commonsourceibias.n208 0.189894
R618 commonsourceibias.n320 commonsourceibias.n208 0.189894
R619 commonsourceibias.n321 commonsourceibias.n320 0.189894
R620 commonsourceibias.n322 commonsourceibias.n321 0.189894
R621 commonsourceibias.n322 commonsourceibias.n206 0.189894
R622 commonsourceibias.n327 commonsourceibias.n206 0.189894
R623 commonsourceibias.n328 commonsourceibias.n327 0.189894
R624 commonsourceibias.n329 commonsourceibias.n328 0.189894
R625 commonsourceibias.n329 commonsourceibias.n204 0.189894
R626 commonsourceibias.n334 commonsourceibias.n204 0.189894
R627 commonsourceibias.n335 commonsourceibias.n334 0.189894
R628 commonsourceibias.n335 commonsourceibias.n202 0.189894
R629 commonsourceibias.n359 commonsourceibias.n354 0.189894
R630 commonsourceibias.n360 commonsourceibias.n359 0.189894
R631 commonsourceibias.n360 commonsourceibias.n352 0.189894
R632 commonsourceibias.n364 commonsourceibias.n352 0.189894
R633 commonsourceibias.n365 commonsourceibias.n364 0.189894
R634 commonsourceibias.n365 commonsourceibias.n350 0.189894
R635 commonsourceibias.n369 commonsourceibias.n350 0.189894
R636 commonsourceibias.n370 commonsourceibias.n369 0.189894
R637 commonsourceibias.n370 commonsourceibias.n348 0.189894
R638 commonsourceibias.n375 commonsourceibias.n348 0.189894
R639 commonsourceibias.n376 commonsourceibias.n375 0.189894
R640 commonsourceibias.n377 commonsourceibias.n376 0.189894
R641 commonsourceibias.n377 commonsourceibias.n346 0.189894
R642 commonsourceibias.n383 commonsourceibias.n346 0.189894
R643 commonsourceibias.n384 commonsourceibias.n383 0.189894
R644 commonsourceibias.n385 commonsourceibias.n384 0.189894
R645 commonsourceibias.n385 commonsourceibias.n344 0.189894
R646 commonsourceibias.n390 commonsourceibias.n344 0.189894
R647 commonsourceibias.n391 commonsourceibias.n390 0.189894
R648 commonsourceibias.n392 commonsourceibias.n391 0.189894
R649 commonsourceibias.n392 commonsourceibias.n342 0.189894
R650 commonsourceibias.n397 commonsourceibias.n342 0.189894
R651 commonsourceibias.n398 commonsourceibias.n397 0.189894
R652 commonsourceibias.n398 commonsourceibias.n340 0.189894
R653 commonsourceibias.n112 commonsourceibias.n111 0.170955
R654 commonsourceibias.n113 commonsourceibias.n112 0.170955
R655 commonsourceibias.n313 commonsourceibias.n237 0.170955
R656 commonsourceibias.n314 commonsourceibias.n313 0.170955
R657 CSoutput.n19 CSoutput.t175 184.661
R658 CSoutput.n78 CSoutput.n77 165.8
R659 CSoutput.n76 CSoutput.n0 165.8
R660 CSoutput.n75 CSoutput.n74 165.8
R661 CSoutput.n73 CSoutput.n72 165.8
R662 CSoutput.n71 CSoutput.n2 165.8
R663 CSoutput.n69 CSoutput.n68 165.8
R664 CSoutput.n67 CSoutput.n3 165.8
R665 CSoutput.n66 CSoutput.n65 165.8
R666 CSoutput.n63 CSoutput.n4 165.8
R667 CSoutput.n61 CSoutput.n60 165.8
R668 CSoutput.n59 CSoutput.n5 165.8
R669 CSoutput.n58 CSoutput.n57 165.8
R670 CSoutput.n55 CSoutput.n6 165.8
R671 CSoutput.n54 CSoutput.n53 165.8
R672 CSoutput.n52 CSoutput.n51 165.8
R673 CSoutput.n50 CSoutput.n8 165.8
R674 CSoutput.n48 CSoutput.n47 165.8
R675 CSoutput.n46 CSoutput.n9 165.8
R676 CSoutput.n45 CSoutput.n44 165.8
R677 CSoutput.n42 CSoutput.n10 165.8
R678 CSoutput.n41 CSoutput.n40 165.8
R679 CSoutput.n39 CSoutput.n38 165.8
R680 CSoutput.n37 CSoutput.n12 165.8
R681 CSoutput.n35 CSoutput.n34 165.8
R682 CSoutput.n33 CSoutput.n13 165.8
R683 CSoutput.n32 CSoutput.n31 165.8
R684 CSoutput.n29 CSoutput.n14 165.8
R685 CSoutput.n28 CSoutput.n27 165.8
R686 CSoutput.n26 CSoutput.n25 165.8
R687 CSoutput.n24 CSoutput.n16 165.8
R688 CSoutput.n22 CSoutput.n21 165.8
R689 CSoutput.n20 CSoutput.n17 165.8
R690 CSoutput.n77 CSoutput.t179 162.194
R691 CSoutput.n18 CSoutput.t184 120.501
R692 CSoutput.n23 CSoutput.t187 120.501
R693 CSoutput.n15 CSoutput.t180 120.501
R694 CSoutput.n30 CSoutput.t174 120.501
R695 CSoutput.n36 CSoutput.t188 120.501
R696 CSoutput.n11 CSoutput.t182 120.501
R697 CSoutput.n43 CSoutput.t176 120.501
R698 CSoutput.n49 CSoutput.t172 120.501
R699 CSoutput.n7 CSoutput.t168 120.501
R700 CSoutput.n56 CSoutput.t181 120.501
R701 CSoutput.n62 CSoutput.t173 120.501
R702 CSoutput.n64 CSoutput.t169 120.501
R703 CSoutput.n70 CSoutput.t183 120.501
R704 CSoutput.n1 CSoutput.t186 120.501
R705 CSoutput.n330 CSoutput.n328 103.469
R706 CSoutput.n310 CSoutput.n308 103.469
R707 CSoutput.n291 CSoutput.n289 103.469
R708 CSoutput.n120 CSoutput.n118 103.469
R709 CSoutput.n100 CSoutput.n98 103.469
R710 CSoutput.n81 CSoutput.n79 103.469
R711 CSoutput.n344 CSoutput.n343 103.111
R712 CSoutput.n342 CSoutput.n341 103.111
R713 CSoutput.n340 CSoutput.n339 103.111
R714 CSoutput.n338 CSoutput.n337 103.111
R715 CSoutput.n336 CSoutput.n335 103.111
R716 CSoutput.n334 CSoutput.n333 103.111
R717 CSoutput.n332 CSoutput.n331 103.111
R718 CSoutput.n330 CSoutput.n329 103.111
R719 CSoutput.n326 CSoutput.n325 103.111
R720 CSoutput.n324 CSoutput.n323 103.111
R721 CSoutput.n322 CSoutput.n321 103.111
R722 CSoutput.n320 CSoutput.n319 103.111
R723 CSoutput.n318 CSoutput.n317 103.111
R724 CSoutput.n316 CSoutput.n315 103.111
R725 CSoutput.n314 CSoutput.n313 103.111
R726 CSoutput.n312 CSoutput.n311 103.111
R727 CSoutput.n310 CSoutput.n309 103.111
R728 CSoutput.n307 CSoutput.n306 103.111
R729 CSoutput.n305 CSoutput.n304 103.111
R730 CSoutput.n303 CSoutput.n302 103.111
R731 CSoutput.n301 CSoutput.n300 103.111
R732 CSoutput.n299 CSoutput.n298 103.111
R733 CSoutput.n297 CSoutput.n296 103.111
R734 CSoutput.n295 CSoutput.n294 103.111
R735 CSoutput.n293 CSoutput.n292 103.111
R736 CSoutput.n291 CSoutput.n290 103.111
R737 CSoutput.n120 CSoutput.n119 103.111
R738 CSoutput.n122 CSoutput.n121 103.111
R739 CSoutput.n124 CSoutput.n123 103.111
R740 CSoutput.n126 CSoutput.n125 103.111
R741 CSoutput.n128 CSoutput.n127 103.111
R742 CSoutput.n130 CSoutput.n129 103.111
R743 CSoutput.n132 CSoutput.n131 103.111
R744 CSoutput.n134 CSoutput.n133 103.111
R745 CSoutput.n136 CSoutput.n135 103.111
R746 CSoutput.n100 CSoutput.n99 103.111
R747 CSoutput.n102 CSoutput.n101 103.111
R748 CSoutput.n104 CSoutput.n103 103.111
R749 CSoutput.n106 CSoutput.n105 103.111
R750 CSoutput.n108 CSoutput.n107 103.111
R751 CSoutput.n110 CSoutput.n109 103.111
R752 CSoutput.n112 CSoutput.n111 103.111
R753 CSoutput.n114 CSoutput.n113 103.111
R754 CSoutput.n116 CSoutput.n115 103.111
R755 CSoutput.n81 CSoutput.n80 103.111
R756 CSoutput.n83 CSoutput.n82 103.111
R757 CSoutput.n85 CSoutput.n84 103.111
R758 CSoutput.n87 CSoutput.n86 103.111
R759 CSoutput.n89 CSoutput.n88 103.111
R760 CSoutput.n91 CSoutput.n90 103.111
R761 CSoutput.n93 CSoutput.n92 103.111
R762 CSoutput.n95 CSoutput.n94 103.111
R763 CSoutput.n97 CSoutput.n96 103.111
R764 CSoutput.n346 CSoutput.n345 103.111
R765 CSoutput.n362 CSoutput.n360 81.5057
R766 CSoutput.n351 CSoutput.n349 81.5057
R767 CSoutput.n386 CSoutput.n384 81.5057
R768 CSoutput.n375 CSoutput.n373 81.5057
R769 CSoutput.n370 CSoutput.n369 80.9324
R770 CSoutput.n368 CSoutput.n367 80.9324
R771 CSoutput.n366 CSoutput.n365 80.9324
R772 CSoutput.n364 CSoutput.n363 80.9324
R773 CSoutput.n362 CSoutput.n361 80.9324
R774 CSoutput.n359 CSoutput.n358 80.9324
R775 CSoutput.n357 CSoutput.n356 80.9324
R776 CSoutput.n355 CSoutput.n354 80.9324
R777 CSoutput.n353 CSoutput.n352 80.9324
R778 CSoutput.n351 CSoutput.n350 80.9324
R779 CSoutput.n386 CSoutput.n385 80.9324
R780 CSoutput.n388 CSoutput.n387 80.9324
R781 CSoutput.n390 CSoutput.n389 80.9324
R782 CSoutput.n392 CSoutput.n391 80.9324
R783 CSoutput.n394 CSoutput.n393 80.9324
R784 CSoutput.n375 CSoutput.n374 80.9324
R785 CSoutput.n377 CSoutput.n376 80.9324
R786 CSoutput.n379 CSoutput.n378 80.9324
R787 CSoutput.n381 CSoutput.n380 80.9324
R788 CSoutput.n383 CSoutput.n382 80.9324
R789 CSoutput.n25 CSoutput.n24 48.1486
R790 CSoutput.n69 CSoutput.n3 48.1486
R791 CSoutput.n38 CSoutput.n37 48.1486
R792 CSoutput.n42 CSoutput.n41 48.1486
R793 CSoutput.n51 CSoutput.n50 48.1486
R794 CSoutput.n55 CSoutput.n54 48.1486
R795 CSoutput.n22 CSoutput.n17 46.462
R796 CSoutput.n72 CSoutput.n71 46.462
R797 CSoutput.n20 CSoutput.n19 44.9055
R798 CSoutput.n29 CSoutput.n28 43.7635
R799 CSoutput.n65 CSoutput.n63 43.7635
R800 CSoutput.n35 CSoutput.n13 41.7396
R801 CSoutput.n57 CSoutput.n5 41.7396
R802 CSoutput.n44 CSoutput.n9 37.0171
R803 CSoutput.n48 CSoutput.n9 37.0171
R804 CSoutput.n76 CSoutput.n75 34.9932
R805 CSoutput.n31 CSoutput.n13 32.2947
R806 CSoutput.n61 CSoutput.n5 32.2947
R807 CSoutput.n30 CSoutput.n29 29.6014
R808 CSoutput.n63 CSoutput.n62 29.6014
R809 CSoutput.n19 CSoutput.n18 28.4085
R810 CSoutput.n18 CSoutput.n17 25.1176
R811 CSoutput.n72 CSoutput.n1 25.1176
R812 CSoutput.n43 CSoutput.n42 22.0922
R813 CSoutput.n50 CSoutput.n49 22.0922
R814 CSoutput.n77 CSoutput.n76 21.8586
R815 CSoutput.n37 CSoutput.n36 18.9681
R816 CSoutput.n56 CSoutput.n55 18.9681
R817 CSoutput.n25 CSoutput.n15 17.6292
R818 CSoutput.n64 CSoutput.n3 17.6292
R819 CSoutput.n24 CSoutput.n23 15.844
R820 CSoutput.n70 CSoutput.n69 15.844
R821 CSoutput.n38 CSoutput.n11 14.5051
R822 CSoutput.n54 CSoutput.n7 14.5051
R823 CSoutput.n397 CSoutput.n78 11.6125
R824 CSoutput.n41 CSoutput.n11 11.3811
R825 CSoutput.n51 CSoutput.n7 11.3811
R826 CSoutput.n23 CSoutput.n22 10.0422
R827 CSoutput.n71 CSoutput.n70 10.0422
R828 CSoutput.n327 CSoutput.n307 9.25285
R829 CSoutput.n117 CSoutput.n97 9.25285
R830 CSoutput.n371 CSoutput.n359 8.97993
R831 CSoutput.n395 CSoutput.n383 8.97993
R832 CSoutput.n372 CSoutput.n348 8.71742
R833 CSoutput.n28 CSoutput.n15 8.25698
R834 CSoutput.n65 CSoutput.n64 8.25698
R835 CSoutput.n372 CSoutput.n371 7.89345
R836 CSoutput.n396 CSoutput.n395 7.89345
R837 CSoutput.n348 CSoutput.n347 7.12641
R838 CSoutput.n138 CSoutput.n137 7.12641
R839 CSoutput.n36 CSoutput.n35 6.91809
R840 CSoutput.n57 CSoutput.n56 6.91809
R841 CSoutput.n371 CSoutput.n370 5.25266
R842 CSoutput.n395 CSoutput.n394 5.25266
R843 CSoutput.n347 CSoutput.n346 5.1449
R844 CSoutput.n327 CSoutput.n326 5.1449
R845 CSoutput.n137 CSoutput.n136 5.1449
R846 CSoutput.n117 CSoutput.n116 5.1449
R847 CSoutput.n397 CSoutput.n138 4.91834
R848 CSoutput.n229 CSoutput.n182 4.5005
R849 CSoutput.n198 CSoutput.n182 4.5005
R850 CSoutput.n193 CSoutput.n177 4.5005
R851 CSoutput.n193 CSoutput.n179 4.5005
R852 CSoutput.n193 CSoutput.n176 4.5005
R853 CSoutput.n193 CSoutput.n180 4.5005
R854 CSoutput.n193 CSoutput.n175 4.5005
R855 CSoutput.n193 CSoutput.t171 4.5005
R856 CSoutput.n193 CSoutput.n174 4.5005
R857 CSoutput.n193 CSoutput.n181 4.5005
R858 CSoutput.n193 CSoutput.n182 4.5005
R859 CSoutput.n191 CSoutput.n177 4.5005
R860 CSoutput.n191 CSoutput.n179 4.5005
R861 CSoutput.n191 CSoutput.n176 4.5005
R862 CSoutput.n191 CSoutput.n180 4.5005
R863 CSoutput.n191 CSoutput.n175 4.5005
R864 CSoutput.n191 CSoutput.t171 4.5005
R865 CSoutput.n191 CSoutput.n174 4.5005
R866 CSoutput.n191 CSoutput.n181 4.5005
R867 CSoutput.n191 CSoutput.n182 4.5005
R868 CSoutput.n190 CSoutput.n177 4.5005
R869 CSoutput.n190 CSoutput.n179 4.5005
R870 CSoutput.n190 CSoutput.n176 4.5005
R871 CSoutput.n190 CSoutput.n180 4.5005
R872 CSoutput.n190 CSoutput.n175 4.5005
R873 CSoutput.n190 CSoutput.t171 4.5005
R874 CSoutput.n190 CSoutput.n174 4.5005
R875 CSoutput.n190 CSoutput.n181 4.5005
R876 CSoutput.n190 CSoutput.n182 4.5005
R877 CSoutput.n275 CSoutput.n177 4.5005
R878 CSoutput.n275 CSoutput.n179 4.5005
R879 CSoutput.n275 CSoutput.n176 4.5005
R880 CSoutput.n275 CSoutput.n180 4.5005
R881 CSoutput.n275 CSoutput.n175 4.5005
R882 CSoutput.n275 CSoutput.t171 4.5005
R883 CSoutput.n275 CSoutput.n174 4.5005
R884 CSoutput.n275 CSoutput.n181 4.5005
R885 CSoutput.n275 CSoutput.n182 4.5005
R886 CSoutput.n273 CSoutput.n177 4.5005
R887 CSoutput.n273 CSoutput.n179 4.5005
R888 CSoutput.n273 CSoutput.n176 4.5005
R889 CSoutput.n273 CSoutput.n180 4.5005
R890 CSoutput.n273 CSoutput.n175 4.5005
R891 CSoutput.n273 CSoutput.t171 4.5005
R892 CSoutput.n273 CSoutput.n174 4.5005
R893 CSoutput.n273 CSoutput.n181 4.5005
R894 CSoutput.n271 CSoutput.n177 4.5005
R895 CSoutput.n271 CSoutput.n179 4.5005
R896 CSoutput.n271 CSoutput.n176 4.5005
R897 CSoutput.n271 CSoutput.n180 4.5005
R898 CSoutput.n271 CSoutput.n175 4.5005
R899 CSoutput.n271 CSoutput.t171 4.5005
R900 CSoutput.n271 CSoutput.n174 4.5005
R901 CSoutput.n271 CSoutput.n181 4.5005
R902 CSoutput.n201 CSoutput.n177 4.5005
R903 CSoutput.n201 CSoutput.n179 4.5005
R904 CSoutput.n201 CSoutput.n176 4.5005
R905 CSoutput.n201 CSoutput.n180 4.5005
R906 CSoutput.n201 CSoutput.n175 4.5005
R907 CSoutput.n201 CSoutput.t171 4.5005
R908 CSoutput.n201 CSoutput.n174 4.5005
R909 CSoutput.n201 CSoutput.n181 4.5005
R910 CSoutput.n201 CSoutput.n182 4.5005
R911 CSoutput.n200 CSoutput.n177 4.5005
R912 CSoutput.n200 CSoutput.n179 4.5005
R913 CSoutput.n200 CSoutput.n176 4.5005
R914 CSoutput.n200 CSoutput.n180 4.5005
R915 CSoutput.n200 CSoutput.n175 4.5005
R916 CSoutput.n200 CSoutput.t171 4.5005
R917 CSoutput.n200 CSoutput.n174 4.5005
R918 CSoutput.n200 CSoutput.n181 4.5005
R919 CSoutput.n200 CSoutput.n182 4.5005
R920 CSoutput.n204 CSoutput.n177 4.5005
R921 CSoutput.n204 CSoutput.n179 4.5005
R922 CSoutput.n204 CSoutput.n176 4.5005
R923 CSoutput.n204 CSoutput.n180 4.5005
R924 CSoutput.n204 CSoutput.n175 4.5005
R925 CSoutput.n204 CSoutput.t171 4.5005
R926 CSoutput.n204 CSoutput.n174 4.5005
R927 CSoutput.n204 CSoutput.n181 4.5005
R928 CSoutput.n204 CSoutput.n182 4.5005
R929 CSoutput.n203 CSoutput.n177 4.5005
R930 CSoutput.n203 CSoutput.n179 4.5005
R931 CSoutput.n203 CSoutput.n176 4.5005
R932 CSoutput.n203 CSoutput.n180 4.5005
R933 CSoutput.n203 CSoutput.n175 4.5005
R934 CSoutput.n203 CSoutput.t171 4.5005
R935 CSoutput.n203 CSoutput.n174 4.5005
R936 CSoutput.n203 CSoutput.n181 4.5005
R937 CSoutput.n203 CSoutput.n182 4.5005
R938 CSoutput.n186 CSoutput.n177 4.5005
R939 CSoutput.n186 CSoutput.n179 4.5005
R940 CSoutput.n186 CSoutput.n176 4.5005
R941 CSoutput.n186 CSoutput.n180 4.5005
R942 CSoutput.n186 CSoutput.n175 4.5005
R943 CSoutput.n186 CSoutput.t171 4.5005
R944 CSoutput.n186 CSoutput.n174 4.5005
R945 CSoutput.n186 CSoutput.n181 4.5005
R946 CSoutput.n186 CSoutput.n182 4.5005
R947 CSoutput.n278 CSoutput.n177 4.5005
R948 CSoutput.n278 CSoutput.n179 4.5005
R949 CSoutput.n278 CSoutput.n176 4.5005
R950 CSoutput.n278 CSoutput.n180 4.5005
R951 CSoutput.n278 CSoutput.n175 4.5005
R952 CSoutput.n278 CSoutput.t171 4.5005
R953 CSoutput.n278 CSoutput.n174 4.5005
R954 CSoutput.n278 CSoutput.n181 4.5005
R955 CSoutput.n278 CSoutput.n182 4.5005
R956 CSoutput.n265 CSoutput.n236 4.5005
R957 CSoutput.n265 CSoutput.n242 4.5005
R958 CSoutput.n223 CSoutput.n212 4.5005
R959 CSoutput.n223 CSoutput.n214 4.5005
R960 CSoutput.n223 CSoutput.n211 4.5005
R961 CSoutput.n223 CSoutput.n215 4.5005
R962 CSoutput.n223 CSoutput.n210 4.5005
R963 CSoutput.n223 CSoutput.t178 4.5005
R964 CSoutput.n223 CSoutput.n209 4.5005
R965 CSoutput.n223 CSoutput.n216 4.5005
R966 CSoutput.n265 CSoutput.n223 4.5005
R967 CSoutput.n244 CSoutput.n212 4.5005
R968 CSoutput.n244 CSoutput.n214 4.5005
R969 CSoutput.n244 CSoutput.n211 4.5005
R970 CSoutput.n244 CSoutput.n215 4.5005
R971 CSoutput.n244 CSoutput.n210 4.5005
R972 CSoutput.n244 CSoutput.t178 4.5005
R973 CSoutput.n244 CSoutput.n209 4.5005
R974 CSoutput.n244 CSoutput.n216 4.5005
R975 CSoutput.n265 CSoutput.n244 4.5005
R976 CSoutput.n222 CSoutput.n212 4.5005
R977 CSoutput.n222 CSoutput.n214 4.5005
R978 CSoutput.n222 CSoutput.n211 4.5005
R979 CSoutput.n222 CSoutput.n215 4.5005
R980 CSoutput.n222 CSoutput.n210 4.5005
R981 CSoutput.n222 CSoutput.t178 4.5005
R982 CSoutput.n222 CSoutput.n209 4.5005
R983 CSoutput.n222 CSoutput.n216 4.5005
R984 CSoutput.n265 CSoutput.n222 4.5005
R985 CSoutput.n246 CSoutput.n212 4.5005
R986 CSoutput.n246 CSoutput.n214 4.5005
R987 CSoutput.n246 CSoutput.n211 4.5005
R988 CSoutput.n246 CSoutput.n215 4.5005
R989 CSoutput.n246 CSoutput.n210 4.5005
R990 CSoutput.n246 CSoutput.t178 4.5005
R991 CSoutput.n246 CSoutput.n209 4.5005
R992 CSoutput.n246 CSoutput.n216 4.5005
R993 CSoutput.n265 CSoutput.n246 4.5005
R994 CSoutput.n212 CSoutput.n207 4.5005
R995 CSoutput.n214 CSoutput.n207 4.5005
R996 CSoutput.n211 CSoutput.n207 4.5005
R997 CSoutput.n215 CSoutput.n207 4.5005
R998 CSoutput.n210 CSoutput.n207 4.5005
R999 CSoutput.t178 CSoutput.n207 4.5005
R1000 CSoutput.n209 CSoutput.n207 4.5005
R1001 CSoutput.n216 CSoutput.n207 4.5005
R1002 CSoutput.n268 CSoutput.n212 4.5005
R1003 CSoutput.n268 CSoutput.n214 4.5005
R1004 CSoutput.n268 CSoutput.n211 4.5005
R1005 CSoutput.n268 CSoutput.n215 4.5005
R1006 CSoutput.n268 CSoutput.n210 4.5005
R1007 CSoutput.n268 CSoutput.t178 4.5005
R1008 CSoutput.n268 CSoutput.n209 4.5005
R1009 CSoutput.n268 CSoutput.n216 4.5005
R1010 CSoutput.n266 CSoutput.n212 4.5005
R1011 CSoutput.n266 CSoutput.n214 4.5005
R1012 CSoutput.n266 CSoutput.n211 4.5005
R1013 CSoutput.n266 CSoutput.n215 4.5005
R1014 CSoutput.n266 CSoutput.n210 4.5005
R1015 CSoutput.n266 CSoutput.t178 4.5005
R1016 CSoutput.n266 CSoutput.n209 4.5005
R1017 CSoutput.n266 CSoutput.n216 4.5005
R1018 CSoutput.n266 CSoutput.n265 4.5005
R1019 CSoutput.n248 CSoutput.n212 4.5005
R1020 CSoutput.n248 CSoutput.n214 4.5005
R1021 CSoutput.n248 CSoutput.n211 4.5005
R1022 CSoutput.n248 CSoutput.n215 4.5005
R1023 CSoutput.n248 CSoutput.n210 4.5005
R1024 CSoutput.n248 CSoutput.t178 4.5005
R1025 CSoutput.n248 CSoutput.n209 4.5005
R1026 CSoutput.n248 CSoutput.n216 4.5005
R1027 CSoutput.n265 CSoutput.n248 4.5005
R1028 CSoutput.n220 CSoutput.n212 4.5005
R1029 CSoutput.n220 CSoutput.n214 4.5005
R1030 CSoutput.n220 CSoutput.n211 4.5005
R1031 CSoutput.n220 CSoutput.n215 4.5005
R1032 CSoutput.n220 CSoutput.n210 4.5005
R1033 CSoutput.n220 CSoutput.t178 4.5005
R1034 CSoutput.n220 CSoutput.n209 4.5005
R1035 CSoutput.n220 CSoutput.n216 4.5005
R1036 CSoutput.n265 CSoutput.n220 4.5005
R1037 CSoutput.n250 CSoutput.n212 4.5005
R1038 CSoutput.n250 CSoutput.n214 4.5005
R1039 CSoutput.n250 CSoutput.n211 4.5005
R1040 CSoutput.n250 CSoutput.n215 4.5005
R1041 CSoutput.n250 CSoutput.n210 4.5005
R1042 CSoutput.n250 CSoutput.t178 4.5005
R1043 CSoutput.n250 CSoutput.n209 4.5005
R1044 CSoutput.n250 CSoutput.n216 4.5005
R1045 CSoutput.n265 CSoutput.n250 4.5005
R1046 CSoutput.n219 CSoutput.n212 4.5005
R1047 CSoutput.n219 CSoutput.n214 4.5005
R1048 CSoutput.n219 CSoutput.n211 4.5005
R1049 CSoutput.n219 CSoutput.n215 4.5005
R1050 CSoutput.n219 CSoutput.n210 4.5005
R1051 CSoutput.n219 CSoutput.t178 4.5005
R1052 CSoutput.n219 CSoutput.n209 4.5005
R1053 CSoutput.n219 CSoutput.n216 4.5005
R1054 CSoutput.n265 CSoutput.n219 4.5005
R1055 CSoutput.n264 CSoutput.n212 4.5005
R1056 CSoutput.n264 CSoutput.n214 4.5005
R1057 CSoutput.n264 CSoutput.n211 4.5005
R1058 CSoutput.n264 CSoutput.n215 4.5005
R1059 CSoutput.n264 CSoutput.n210 4.5005
R1060 CSoutput.n264 CSoutput.t178 4.5005
R1061 CSoutput.n264 CSoutput.n209 4.5005
R1062 CSoutput.n264 CSoutput.n216 4.5005
R1063 CSoutput.n265 CSoutput.n264 4.5005
R1064 CSoutput.n263 CSoutput.n148 4.5005
R1065 CSoutput.n164 CSoutput.n148 4.5005
R1066 CSoutput.n159 CSoutput.n143 4.5005
R1067 CSoutput.n159 CSoutput.n145 4.5005
R1068 CSoutput.n159 CSoutput.n142 4.5005
R1069 CSoutput.n159 CSoutput.n146 4.5005
R1070 CSoutput.n159 CSoutput.n141 4.5005
R1071 CSoutput.n159 CSoutput.t185 4.5005
R1072 CSoutput.n159 CSoutput.n140 4.5005
R1073 CSoutput.n159 CSoutput.n147 4.5005
R1074 CSoutput.n159 CSoutput.n148 4.5005
R1075 CSoutput.n157 CSoutput.n143 4.5005
R1076 CSoutput.n157 CSoutput.n145 4.5005
R1077 CSoutput.n157 CSoutput.n142 4.5005
R1078 CSoutput.n157 CSoutput.n146 4.5005
R1079 CSoutput.n157 CSoutput.n141 4.5005
R1080 CSoutput.n157 CSoutput.t185 4.5005
R1081 CSoutput.n157 CSoutput.n140 4.5005
R1082 CSoutput.n157 CSoutput.n147 4.5005
R1083 CSoutput.n157 CSoutput.n148 4.5005
R1084 CSoutput.n156 CSoutput.n143 4.5005
R1085 CSoutput.n156 CSoutput.n145 4.5005
R1086 CSoutput.n156 CSoutput.n142 4.5005
R1087 CSoutput.n156 CSoutput.n146 4.5005
R1088 CSoutput.n156 CSoutput.n141 4.5005
R1089 CSoutput.n156 CSoutput.t185 4.5005
R1090 CSoutput.n156 CSoutput.n140 4.5005
R1091 CSoutput.n156 CSoutput.n147 4.5005
R1092 CSoutput.n156 CSoutput.n148 4.5005
R1093 CSoutput.n285 CSoutput.n143 4.5005
R1094 CSoutput.n285 CSoutput.n145 4.5005
R1095 CSoutput.n285 CSoutput.n142 4.5005
R1096 CSoutput.n285 CSoutput.n146 4.5005
R1097 CSoutput.n285 CSoutput.n141 4.5005
R1098 CSoutput.n285 CSoutput.t185 4.5005
R1099 CSoutput.n285 CSoutput.n140 4.5005
R1100 CSoutput.n285 CSoutput.n147 4.5005
R1101 CSoutput.n285 CSoutput.n148 4.5005
R1102 CSoutput.n283 CSoutput.n143 4.5005
R1103 CSoutput.n283 CSoutput.n145 4.5005
R1104 CSoutput.n283 CSoutput.n142 4.5005
R1105 CSoutput.n283 CSoutput.n146 4.5005
R1106 CSoutput.n283 CSoutput.n141 4.5005
R1107 CSoutput.n283 CSoutput.t185 4.5005
R1108 CSoutput.n283 CSoutput.n140 4.5005
R1109 CSoutput.n283 CSoutput.n147 4.5005
R1110 CSoutput.n281 CSoutput.n143 4.5005
R1111 CSoutput.n281 CSoutput.n145 4.5005
R1112 CSoutput.n281 CSoutput.n142 4.5005
R1113 CSoutput.n281 CSoutput.n146 4.5005
R1114 CSoutput.n281 CSoutput.n141 4.5005
R1115 CSoutput.n281 CSoutput.t185 4.5005
R1116 CSoutput.n281 CSoutput.n140 4.5005
R1117 CSoutput.n281 CSoutput.n147 4.5005
R1118 CSoutput.n167 CSoutput.n143 4.5005
R1119 CSoutput.n167 CSoutput.n145 4.5005
R1120 CSoutput.n167 CSoutput.n142 4.5005
R1121 CSoutput.n167 CSoutput.n146 4.5005
R1122 CSoutput.n167 CSoutput.n141 4.5005
R1123 CSoutput.n167 CSoutput.t185 4.5005
R1124 CSoutput.n167 CSoutput.n140 4.5005
R1125 CSoutput.n167 CSoutput.n147 4.5005
R1126 CSoutput.n167 CSoutput.n148 4.5005
R1127 CSoutput.n166 CSoutput.n143 4.5005
R1128 CSoutput.n166 CSoutput.n145 4.5005
R1129 CSoutput.n166 CSoutput.n142 4.5005
R1130 CSoutput.n166 CSoutput.n146 4.5005
R1131 CSoutput.n166 CSoutput.n141 4.5005
R1132 CSoutput.n166 CSoutput.t185 4.5005
R1133 CSoutput.n166 CSoutput.n140 4.5005
R1134 CSoutput.n166 CSoutput.n147 4.5005
R1135 CSoutput.n166 CSoutput.n148 4.5005
R1136 CSoutput.n170 CSoutput.n143 4.5005
R1137 CSoutput.n170 CSoutput.n145 4.5005
R1138 CSoutput.n170 CSoutput.n142 4.5005
R1139 CSoutput.n170 CSoutput.n146 4.5005
R1140 CSoutput.n170 CSoutput.n141 4.5005
R1141 CSoutput.n170 CSoutput.t185 4.5005
R1142 CSoutput.n170 CSoutput.n140 4.5005
R1143 CSoutput.n170 CSoutput.n147 4.5005
R1144 CSoutput.n170 CSoutput.n148 4.5005
R1145 CSoutput.n169 CSoutput.n143 4.5005
R1146 CSoutput.n169 CSoutput.n145 4.5005
R1147 CSoutput.n169 CSoutput.n142 4.5005
R1148 CSoutput.n169 CSoutput.n146 4.5005
R1149 CSoutput.n169 CSoutput.n141 4.5005
R1150 CSoutput.n169 CSoutput.t185 4.5005
R1151 CSoutput.n169 CSoutput.n140 4.5005
R1152 CSoutput.n169 CSoutput.n147 4.5005
R1153 CSoutput.n169 CSoutput.n148 4.5005
R1154 CSoutput.n152 CSoutput.n143 4.5005
R1155 CSoutput.n152 CSoutput.n145 4.5005
R1156 CSoutput.n152 CSoutput.n142 4.5005
R1157 CSoutput.n152 CSoutput.n146 4.5005
R1158 CSoutput.n152 CSoutput.n141 4.5005
R1159 CSoutput.n152 CSoutput.t185 4.5005
R1160 CSoutput.n152 CSoutput.n140 4.5005
R1161 CSoutput.n152 CSoutput.n147 4.5005
R1162 CSoutput.n152 CSoutput.n148 4.5005
R1163 CSoutput.n288 CSoutput.n143 4.5005
R1164 CSoutput.n288 CSoutput.n145 4.5005
R1165 CSoutput.n288 CSoutput.n142 4.5005
R1166 CSoutput.n288 CSoutput.n146 4.5005
R1167 CSoutput.n288 CSoutput.n141 4.5005
R1168 CSoutput.n288 CSoutput.t185 4.5005
R1169 CSoutput.n288 CSoutput.n140 4.5005
R1170 CSoutput.n288 CSoutput.n147 4.5005
R1171 CSoutput.n288 CSoutput.n148 4.5005
R1172 CSoutput.n347 CSoutput.n327 4.10845
R1173 CSoutput.n137 CSoutput.n117 4.10845
R1174 CSoutput.n345 CSoutput.t157 4.06363
R1175 CSoutput.n345 CSoutput.t79 4.06363
R1176 CSoutput.n343 CSoutput.t1 4.06363
R1177 CSoutput.n343 CSoutput.t101 4.06363
R1178 CSoutput.n341 CSoutput.t29 4.06363
R1179 CSoutput.n341 CSoutput.t14 4.06363
R1180 CSoutput.n339 CSoutput.t55 4.06363
R1181 CSoutput.n339 CSoutput.t19 4.06363
R1182 CSoutput.n337 CSoutput.t95 4.06363
R1183 CSoutput.n337 CSoutput.t12 4.06363
R1184 CSoutput.n335 CSoutput.t40 4.06363
R1185 CSoutput.n335 CSoutput.t63 4.06363
R1186 CSoutput.n333 CSoutput.t48 4.06363
R1187 CSoutput.n333 CSoutput.t36 4.06363
R1188 CSoutput.n331 CSoutput.t100 4.06363
R1189 CSoutput.n331 CSoutput.t5 4.06363
R1190 CSoutput.n329 CSoutput.t53 4.06363
R1191 CSoutput.n329 CSoutput.t21 4.06363
R1192 CSoutput.n328 CSoutput.t28 4.06363
R1193 CSoutput.n328 CSoutput.t103 4.06363
R1194 CSoutput.n325 CSoutput.t59 4.06363
R1195 CSoutput.n325 CSoutput.t58 4.06363
R1196 CSoutput.n323 CSoutput.t52 4.06363
R1197 CSoutput.n323 CSoutput.t20 4.06363
R1198 CSoutput.n321 CSoutput.t39 4.06363
R1199 CSoutput.n321 CSoutput.t27 4.06363
R1200 CSoutput.n319 CSoutput.t7 4.06363
R1201 CSoutput.n319 CSoutput.t49 4.06363
R1202 CSoutput.n317 CSoutput.t32 4.06363
R1203 CSoutput.n317 CSoutput.t31 4.06363
R1204 CSoutput.n315 CSoutput.t87 4.06363
R1205 CSoutput.n315 CSoutput.t160 4.06363
R1206 CSoutput.n313 CSoutput.t9 4.06363
R1207 CSoutput.n313 CSoutput.t71 4.06363
R1208 CSoutput.n311 CSoutput.t155 4.06363
R1209 CSoutput.n311 CSoutput.t13 4.06363
R1210 CSoutput.n309 CSoutput.t26 4.06363
R1211 CSoutput.n309 CSoutput.t34 4.06363
R1212 CSoutput.n308 CSoutput.t38 4.06363
R1213 CSoutput.n308 CSoutput.t75 4.06363
R1214 CSoutput.n306 CSoutput.t98 4.06363
R1215 CSoutput.n306 CSoutput.t73 4.06363
R1216 CSoutput.n304 CSoutput.t66 4.06363
R1217 CSoutput.n304 CSoutput.t0 4.06363
R1218 CSoutput.n302 CSoutput.t102 4.06363
R1219 CSoutput.n302 CSoutput.t3 4.06363
R1220 CSoutput.n300 CSoutput.t152 4.06363
R1221 CSoutput.n300 CSoutput.t62 4.06363
R1222 CSoutput.n298 CSoutput.t70 4.06363
R1223 CSoutput.n298 CSoutput.t60 4.06363
R1224 CSoutput.n296 CSoutput.t99 4.06363
R1225 CSoutput.n296 CSoutput.t47 4.06363
R1226 CSoutput.n294 CSoutput.t94 4.06363
R1227 CSoutput.n294 CSoutput.t162 4.06363
R1228 CSoutput.n292 CSoutput.t91 4.06363
R1229 CSoutput.n292 CSoutput.t4 4.06363
R1230 CSoutput.n290 CSoutput.t154 4.06363
R1231 CSoutput.n290 CSoutput.t68 4.06363
R1232 CSoutput.n289 CSoutput.t8 4.06363
R1233 CSoutput.n289 CSoutput.t6 4.06363
R1234 CSoutput.n118 CSoutput.t10 4.06363
R1235 CSoutput.n118 CSoutput.t80 4.06363
R1236 CSoutput.n119 CSoutput.t166 4.06363
R1237 CSoutput.n119 CSoutput.t158 4.06363
R1238 CSoutput.n121 CSoutput.t84 4.06363
R1239 CSoutput.n121 CSoutput.t22 4.06363
R1240 CSoutput.n123 CSoutput.t167 4.06363
R1241 CSoutput.n123 CSoutput.t82 4.06363
R1242 CSoutput.n125 CSoutput.t92 4.06363
R1243 CSoutput.n125 CSoutput.t164 4.06363
R1244 CSoutput.n127 CSoutput.t54 4.06363
R1245 CSoutput.n127 CSoutput.t69 4.06363
R1246 CSoutput.n129 CSoutput.t88 4.06363
R1247 CSoutput.n129 CSoutput.t72 4.06363
R1248 CSoutput.n131 CSoutput.t159 4.06363
R1249 CSoutput.n131 CSoutput.t163 4.06363
R1250 CSoutput.n133 CSoutput.t23 4.06363
R1251 CSoutput.n133 CSoutput.t86 4.06363
R1252 CSoutput.n135 CSoutput.t11 4.06363
R1253 CSoutput.n135 CSoutput.t85 4.06363
R1254 CSoutput.n98 CSoutput.t57 4.06363
R1255 CSoutput.n98 CSoutput.t43 4.06363
R1256 CSoutput.n99 CSoutput.t50 4.06363
R1257 CSoutput.n99 CSoutput.t65 4.06363
R1258 CSoutput.n101 CSoutput.t25 4.06363
R1259 CSoutput.n101 CSoutput.t78 4.06363
R1260 CSoutput.n103 CSoutput.t51 4.06363
R1261 CSoutput.n103 CSoutput.t41 4.06363
R1262 CSoutput.n105 CSoutput.t33 4.06363
R1263 CSoutput.n105 CSoutput.t81 4.06363
R1264 CSoutput.n107 CSoutput.t161 4.06363
R1265 CSoutput.n107 CSoutput.t67 4.06363
R1266 CSoutput.n109 CSoutput.t74 4.06363
R1267 CSoutput.n109 CSoutput.t18 4.06363
R1268 CSoutput.n111 CSoutput.t56 4.06363
R1269 CSoutput.n111 CSoutput.t42 4.06363
R1270 CSoutput.n113 CSoutput.t156 4.06363
R1271 CSoutput.n113 CSoutput.t96 4.06363
R1272 CSoutput.n115 CSoutput.t24 4.06363
R1273 CSoutput.n115 CSoutput.t16 4.06363
R1274 CSoutput.n79 CSoutput.t30 4.06363
R1275 CSoutput.n79 CSoutput.t17 4.06363
R1276 CSoutput.n80 CSoutput.t83 4.06363
R1277 CSoutput.n80 CSoutput.t153 4.06363
R1278 CSoutput.n82 CSoutput.t15 4.06363
R1279 CSoutput.n82 CSoutput.t90 4.06363
R1280 CSoutput.n84 CSoutput.t45 4.06363
R1281 CSoutput.n84 CSoutput.t64 4.06363
R1282 CSoutput.n86 CSoutput.t46 4.06363
R1283 CSoutput.n86 CSoutput.t77 4.06363
R1284 CSoutput.n88 CSoutput.t61 4.06363
R1285 CSoutput.n88 CSoutput.t35 4.06363
R1286 CSoutput.n90 CSoutput.t165 4.06363
R1287 CSoutput.n90 CSoutput.t97 4.06363
R1288 CSoutput.n92 CSoutput.t2 4.06363
R1289 CSoutput.n92 CSoutput.t89 4.06363
R1290 CSoutput.n94 CSoutput.t44 4.06363
R1291 CSoutput.n94 CSoutput.t37 4.06363
R1292 CSoutput.n96 CSoutput.t93 4.06363
R1293 CSoutput.n96 CSoutput.t76 4.06363
R1294 CSoutput.n44 CSoutput.n43 3.79402
R1295 CSoutput.n49 CSoutput.n48 3.79402
R1296 CSoutput.n397 CSoutput.n396 3.78008
R1297 CSoutput.n348 CSoutput.n138 3.19963
R1298 CSoutput.n369 CSoutput.t116 2.82907
R1299 CSoutput.n369 CSoutput.t106 2.82907
R1300 CSoutput.n367 CSoutput.t117 2.82907
R1301 CSoutput.n367 CSoutput.t145 2.82907
R1302 CSoutput.n365 CSoutput.t137 2.82907
R1303 CSoutput.n365 CSoutput.t114 2.82907
R1304 CSoutput.n363 CSoutput.t147 2.82907
R1305 CSoutput.n363 CSoutput.t121 2.82907
R1306 CSoutput.n361 CSoutput.t150 2.82907
R1307 CSoutput.n361 CSoutput.t140 2.82907
R1308 CSoutput.n360 CSoutput.t112 2.82907
R1309 CSoutput.n360 CSoutput.t126 2.82907
R1310 CSoutput.n358 CSoutput.t148 2.82907
R1311 CSoutput.n358 CSoutput.t113 2.82907
R1312 CSoutput.n356 CSoutput.t146 2.82907
R1313 CSoutput.n356 CSoutput.t120 2.82907
R1314 CSoutput.n354 CSoutput.t110 2.82907
R1315 CSoutput.n354 CSoutput.t143 2.82907
R1316 CSoutput.n352 CSoutput.t122 2.82907
R1317 CSoutput.n352 CSoutput.t128 2.82907
R1318 CSoutput.n350 CSoutput.t105 2.82907
R1319 CSoutput.n350 CSoutput.t107 2.82907
R1320 CSoutput.n349 CSoutput.t142 2.82907
R1321 CSoutput.n349 CSoutput.t134 2.82907
R1322 CSoutput.n384 CSoutput.t130 2.82907
R1323 CSoutput.n384 CSoutput.t124 2.82907
R1324 CSoutput.n385 CSoutput.t104 2.82907
R1325 CSoutput.n385 CSoutput.t135 2.82907
R1326 CSoutput.n387 CSoutput.t139 2.82907
R1327 CSoutput.n387 CSoutput.t119 2.82907
R1328 CSoutput.n389 CSoutput.t125 2.82907
R1329 CSoutput.n389 CSoutput.t129 2.82907
R1330 CSoutput.n391 CSoutput.t133 2.82907
R1331 CSoutput.n391 CSoutput.t144 2.82907
R1332 CSoutput.n393 CSoutput.t149 2.82907
R1333 CSoutput.n393 CSoutput.t108 2.82907
R1334 CSoutput.n373 CSoutput.t136 2.82907
R1335 CSoutput.n373 CSoutput.t131 2.82907
R1336 CSoutput.n374 CSoutput.t111 2.82907
R1337 CSoutput.n374 CSoutput.t109 2.82907
R1338 CSoutput.n376 CSoutput.t151 2.82907
R1339 CSoutput.n376 CSoutput.t127 2.82907
R1340 CSoutput.n378 CSoutput.t132 2.82907
R1341 CSoutput.n378 CSoutput.t141 2.82907
R1342 CSoutput.n380 CSoutput.t138 2.82907
R1343 CSoutput.n380 CSoutput.t118 2.82907
R1344 CSoutput.n382 CSoutput.t123 2.82907
R1345 CSoutput.n382 CSoutput.t115 2.82907
R1346 CSoutput.n396 CSoutput.n372 2.75627
R1347 CSoutput.n75 CSoutput.n1 2.45513
R1348 CSoutput.n229 CSoutput.n227 2.251
R1349 CSoutput.n229 CSoutput.n226 2.251
R1350 CSoutput.n229 CSoutput.n225 2.251
R1351 CSoutput.n229 CSoutput.n224 2.251
R1352 CSoutput.n198 CSoutput.n197 2.251
R1353 CSoutput.n198 CSoutput.n196 2.251
R1354 CSoutput.n198 CSoutput.n195 2.251
R1355 CSoutput.n198 CSoutput.n194 2.251
R1356 CSoutput.n271 CSoutput.n270 2.251
R1357 CSoutput.n236 CSoutput.n234 2.251
R1358 CSoutput.n236 CSoutput.n233 2.251
R1359 CSoutput.n236 CSoutput.n232 2.251
R1360 CSoutput.n254 CSoutput.n236 2.251
R1361 CSoutput.n242 CSoutput.n241 2.251
R1362 CSoutput.n242 CSoutput.n240 2.251
R1363 CSoutput.n242 CSoutput.n239 2.251
R1364 CSoutput.n242 CSoutput.n238 2.251
R1365 CSoutput.n268 CSoutput.n208 2.251
R1366 CSoutput.n263 CSoutput.n261 2.251
R1367 CSoutput.n263 CSoutput.n260 2.251
R1368 CSoutput.n263 CSoutput.n259 2.251
R1369 CSoutput.n263 CSoutput.n258 2.251
R1370 CSoutput.n164 CSoutput.n163 2.251
R1371 CSoutput.n164 CSoutput.n162 2.251
R1372 CSoutput.n164 CSoutput.n161 2.251
R1373 CSoutput.n164 CSoutput.n160 2.251
R1374 CSoutput.n281 CSoutput.n280 2.251
R1375 CSoutput.n198 CSoutput.n178 2.2505
R1376 CSoutput.n193 CSoutput.n178 2.2505
R1377 CSoutput.n191 CSoutput.n178 2.2505
R1378 CSoutput.n190 CSoutput.n178 2.2505
R1379 CSoutput.n275 CSoutput.n178 2.2505
R1380 CSoutput.n273 CSoutput.n178 2.2505
R1381 CSoutput.n271 CSoutput.n178 2.2505
R1382 CSoutput.n201 CSoutput.n178 2.2505
R1383 CSoutput.n200 CSoutput.n178 2.2505
R1384 CSoutput.n204 CSoutput.n178 2.2505
R1385 CSoutput.n203 CSoutput.n178 2.2505
R1386 CSoutput.n186 CSoutput.n178 2.2505
R1387 CSoutput.n278 CSoutput.n178 2.2505
R1388 CSoutput.n278 CSoutput.n277 2.2505
R1389 CSoutput.n242 CSoutput.n213 2.2505
R1390 CSoutput.n223 CSoutput.n213 2.2505
R1391 CSoutput.n244 CSoutput.n213 2.2505
R1392 CSoutput.n222 CSoutput.n213 2.2505
R1393 CSoutput.n246 CSoutput.n213 2.2505
R1394 CSoutput.n213 CSoutput.n207 2.2505
R1395 CSoutput.n268 CSoutput.n213 2.2505
R1396 CSoutput.n266 CSoutput.n213 2.2505
R1397 CSoutput.n248 CSoutput.n213 2.2505
R1398 CSoutput.n220 CSoutput.n213 2.2505
R1399 CSoutput.n250 CSoutput.n213 2.2505
R1400 CSoutput.n219 CSoutput.n213 2.2505
R1401 CSoutput.n264 CSoutput.n213 2.2505
R1402 CSoutput.n264 CSoutput.n217 2.2505
R1403 CSoutput.n164 CSoutput.n144 2.2505
R1404 CSoutput.n159 CSoutput.n144 2.2505
R1405 CSoutput.n157 CSoutput.n144 2.2505
R1406 CSoutput.n156 CSoutput.n144 2.2505
R1407 CSoutput.n285 CSoutput.n144 2.2505
R1408 CSoutput.n283 CSoutput.n144 2.2505
R1409 CSoutput.n281 CSoutput.n144 2.2505
R1410 CSoutput.n167 CSoutput.n144 2.2505
R1411 CSoutput.n166 CSoutput.n144 2.2505
R1412 CSoutput.n170 CSoutput.n144 2.2505
R1413 CSoutput.n169 CSoutput.n144 2.2505
R1414 CSoutput.n152 CSoutput.n144 2.2505
R1415 CSoutput.n288 CSoutput.n144 2.2505
R1416 CSoutput.n288 CSoutput.n287 2.2505
R1417 CSoutput.n206 CSoutput.n199 2.25024
R1418 CSoutput.n206 CSoutput.n192 2.25024
R1419 CSoutput.n274 CSoutput.n206 2.25024
R1420 CSoutput.n206 CSoutput.n202 2.25024
R1421 CSoutput.n206 CSoutput.n205 2.25024
R1422 CSoutput.n206 CSoutput.n173 2.25024
R1423 CSoutput.n256 CSoutput.n253 2.25024
R1424 CSoutput.n256 CSoutput.n252 2.25024
R1425 CSoutput.n256 CSoutput.n251 2.25024
R1426 CSoutput.n256 CSoutput.n218 2.25024
R1427 CSoutput.n256 CSoutput.n255 2.25024
R1428 CSoutput.n257 CSoutput.n256 2.25024
R1429 CSoutput.n172 CSoutput.n165 2.25024
R1430 CSoutput.n172 CSoutput.n158 2.25024
R1431 CSoutput.n284 CSoutput.n172 2.25024
R1432 CSoutput.n172 CSoutput.n168 2.25024
R1433 CSoutput.n172 CSoutput.n171 2.25024
R1434 CSoutput.n172 CSoutput.n139 2.25024
R1435 CSoutput.n273 CSoutput.n183 1.50111
R1436 CSoutput.n221 CSoutput.n207 1.50111
R1437 CSoutput.n283 CSoutput.n149 1.50111
R1438 CSoutput.n229 CSoutput.n228 1.501
R1439 CSoutput.n236 CSoutput.n235 1.501
R1440 CSoutput.n263 CSoutput.n262 1.501
R1441 CSoutput.n277 CSoutput.n188 1.12536
R1442 CSoutput.n277 CSoutput.n189 1.12536
R1443 CSoutput.n277 CSoutput.n276 1.12536
R1444 CSoutput.n237 CSoutput.n217 1.12536
R1445 CSoutput.n243 CSoutput.n217 1.12536
R1446 CSoutput.n245 CSoutput.n217 1.12536
R1447 CSoutput.n287 CSoutput.n154 1.12536
R1448 CSoutput.n287 CSoutput.n155 1.12536
R1449 CSoutput.n287 CSoutput.n286 1.12536
R1450 CSoutput.n277 CSoutput.n184 1.12536
R1451 CSoutput.n277 CSoutput.n185 1.12536
R1452 CSoutput.n277 CSoutput.n187 1.12536
R1453 CSoutput.n267 CSoutput.n217 1.12536
R1454 CSoutput.n247 CSoutput.n217 1.12536
R1455 CSoutput.n249 CSoutput.n217 1.12536
R1456 CSoutput.n287 CSoutput.n150 1.12536
R1457 CSoutput.n287 CSoutput.n151 1.12536
R1458 CSoutput.n287 CSoutput.n153 1.12536
R1459 CSoutput.n31 CSoutput.n30 0.669944
R1460 CSoutput.n62 CSoutput.n61 0.669944
R1461 CSoutput.n364 CSoutput.n362 0.573776
R1462 CSoutput.n366 CSoutput.n364 0.573776
R1463 CSoutput.n368 CSoutput.n366 0.573776
R1464 CSoutput.n370 CSoutput.n368 0.573776
R1465 CSoutput.n353 CSoutput.n351 0.573776
R1466 CSoutput.n355 CSoutput.n353 0.573776
R1467 CSoutput.n357 CSoutput.n355 0.573776
R1468 CSoutput.n359 CSoutput.n357 0.573776
R1469 CSoutput.n394 CSoutput.n392 0.573776
R1470 CSoutput.n392 CSoutput.n390 0.573776
R1471 CSoutput.n390 CSoutput.n388 0.573776
R1472 CSoutput.n388 CSoutput.n386 0.573776
R1473 CSoutput.n383 CSoutput.n381 0.573776
R1474 CSoutput.n381 CSoutput.n379 0.573776
R1475 CSoutput.n379 CSoutput.n377 0.573776
R1476 CSoutput.n377 CSoutput.n375 0.573776
R1477 CSoutput.n397 CSoutput.n288 0.534303
R1478 CSoutput.n332 CSoutput.n330 0.358259
R1479 CSoutput.n334 CSoutput.n332 0.358259
R1480 CSoutput.n336 CSoutput.n334 0.358259
R1481 CSoutput.n338 CSoutput.n336 0.358259
R1482 CSoutput.n340 CSoutput.n338 0.358259
R1483 CSoutput.n342 CSoutput.n340 0.358259
R1484 CSoutput.n344 CSoutput.n342 0.358259
R1485 CSoutput.n346 CSoutput.n344 0.358259
R1486 CSoutput.n312 CSoutput.n310 0.358259
R1487 CSoutput.n314 CSoutput.n312 0.358259
R1488 CSoutput.n316 CSoutput.n314 0.358259
R1489 CSoutput.n318 CSoutput.n316 0.358259
R1490 CSoutput.n320 CSoutput.n318 0.358259
R1491 CSoutput.n322 CSoutput.n320 0.358259
R1492 CSoutput.n324 CSoutput.n322 0.358259
R1493 CSoutput.n326 CSoutput.n324 0.358259
R1494 CSoutput.n293 CSoutput.n291 0.358259
R1495 CSoutput.n295 CSoutput.n293 0.358259
R1496 CSoutput.n297 CSoutput.n295 0.358259
R1497 CSoutput.n299 CSoutput.n297 0.358259
R1498 CSoutput.n301 CSoutput.n299 0.358259
R1499 CSoutput.n303 CSoutput.n301 0.358259
R1500 CSoutput.n305 CSoutput.n303 0.358259
R1501 CSoutput.n307 CSoutput.n305 0.358259
R1502 CSoutput.n136 CSoutput.n134 0.358259
R1503 CSoutput.n134 CSoutput.n132 0.358259
R1504 CSoutput.n132 CSoutput.n130 0.358259
R1505 CSoutput.n130 CSoutput.n128 0.358259
R1506 CSoutput.n128 CSoutput.n126 0.358259
R1507 CSoutput.n126 CSoutput.n124 0.358259
R1508 CSoutput.n124 CSoutput.n122 0.358259
R1509 CSoutput.n122 CSoutput.n120 0.358259
R1510 CSoutput.n116 CSoutput.n114 0.358259
R1511 CSoutput.n114 CSoutput.n112 0.358259
R1512 CSoutput.n112 CSoutput.n110 0.358259
R1513 CSoutput.n110 CSoutput.n108 0.358259
R1514 CSoutput.n108 CSoutput.n106 0.358259
R1515 CSoutput.n106 CSoutput.n104 0.358259
R1516 CSoutput.n104 CSoutput.n102 0.358259
R1517 CSoutput.n102 CSoutput.n100 0.358259
R1518 CSoutput.n97 CSoutput.n95 0.358259
R1519 CSoutput.n95 CSoutput.n93 0.358259
R1520 CSoutput.n93 CSoutput.n91 0.358259
R1521 CSoutput.n91 CSoutput.n89 0.358259
R1522 CSoutput.n89 CSoutput.n87 0.358259
R1523 CSoutput.n87 CSoutput.n85 0.358259
R1524 CSoutput.n85 CSoutput.n83 0.358259
R1525 CSoutput.n83 CSoutput.n81 0.358259
R1526 CSoutput.n21 CSoutput.n20 0.169105
R1527 CSoutput.n21 CSoutput.n16 0.169105
R1528 CSoutput.n26 CSoutput.n16 0.169105
R1529 CSoutput.n27 CSoutput.n26 0.169105
R1530 CSoutput.n27 CSoutput.n14 0.169105
R1531 CSoutput.n32 CSoutput.n14 0.169105
R1532 CSoutput.n33 CSoutput.n32 0.169105
R1533 CSoutput.n34 CSoutput.n33 0.169105
R1534 CSoutput.n34 CSoutput.n12 0.169105
R1535 CSoutput.n39 CSoutput.n12 0.169105
R1536 CSoutput.n40 CSoutput.n39 0.169105
R1537 CSoutput.n40 CSoutput.n10 0.169105
R1538 CSoutput.n45 CSoutput.n10 0.169105
R1539 CSoutput.n46 CSoutput.n45 0.169105
R1540 CSoutput.n47 CSoutput.n46 0.169105
R1541 CSoutput.n47 CSoutput.n8 0.169105
R1542 CSoutput.n52 CSoutput.n8 0.169105
R1543 CSoutput.n53 CSoutput.n52 0.169105
R1544 CSoutput.n53 CSoutput.n6 0.169105
R1545 CSoutput.n58 CSoutput.n6 0.169105
R1546 CSoutput.n59 CSoutput.n58 0.169105
R1547 CSoutput.n60 CSoutput.n59 0.169105
R1548 CSoutput.n60 CSoutput.n4 0.169105
R1549 CSoutput.n66 CSoutput.n4 0.169105
R1550 CSoutput.n67 CSoutput.n66 0.169105
R1551 CSoutput.n68 CSoutput.n67 0.169105
R1552 CSoutput.n68 CSoutput.n2 0.169105
R1553 CSoutput.n73 CSoutput.n2 0.169105
R1554 CSoutput.n74 CSoutput.n73 0.169105
R1555 CSoutput.n74 CSoutput.n0 0.169105
R1556 CSoutput.n78 CSoutput.n0 0.169105
R1557 CSoutput.n231 CSoutput.n230 0.0910737
R1558 CSoutput.n282 CSoutput.n279 0.0723685
R1559 CSoutput.n236 CSoutput.n231 0.0522944
R1560 CSoutput.n279 CSoutput.n278 0.0499135
R1561 CSoutput.n230 CSoutput.n229 0.0499135
R1562 CSoutput.n264 CSoutput.n263 0.0464294
R1563 CSoutput.n272 CSoutput.n269 0.0391444
R1564 CSoutput.n231 CSoutput.t189 0.023435
R1565 CSoutput.n279 CSoutput.t170 0.02262
R1566 CSoutput.n230 CSoutput.t177 0.02262
R1567 CSoutput CSoutput.n397 0.0052
R1568 CSoutput.n201 CSoutput.n184 0.00365111
R1569 CSoutput.n204 CSoutput.n185 0.00365111
R1570 CSoutput.n187 CSoutput.n186 0.00365111
R1571 CSoutput.n229 CSoutput.n188 0.00365111
R1572 CSoutput.n193 CSoutput.n189 0.00365111
R1573 CSoutput.n276 CSoutput.n190 0.00365111
R1574 CSoutput.n267 CSoutput.n266 0.00365111
R1575 CSoutput.n247 CSoutput.n220 0.00365111
R1576 CSoutput.n249 CSoutput.n219 0.00365111
R1577 CSoutput.n237 CSoutput.n236 0.00365111
R1578 CSoutput.n243 CSoutput.n223 0.00365111
R1579 CSoutput.n245 CSoutput.n222 0.00365111
R1580 CSoutput.n167 CSoutput.n150 0.00365111
R1581 CSoutput.n170 CSoutput.n151 0.00365111
R1582 CSoutput.n153 CSoutput.n152 0.00365111
R1583 CSoutput.n263 CSoutput.n154 0.00365111
R1584 CSoutput.n159 CSoutput.n155 0.00365111
R1585 CSoutput.n286 CSoutput.n156 0.00365111
R1586 CSoutput.n198 CSoutput.n188 0.00340054
R1587 CSoutput.n191 CSoutput.n189 0.00340054
R1588 CSoutput.n276 CSoutput.n275 0.00340054
R1589 CSoutput.n271 CSoutput.n184 0.00340054
R1590 CSoutput.n200 CSoutput.n185 0.00340054
R1591 CSoutput.n203 CSoutput.n187 0.00340054
R1592 CSoutput.n242 CSoutput.n237 0.00340054
R1593 CSoutput.n244 CSoutput.n243 0.00340054
R1594 CSoutput.n246 CSoutput.n245 0.00340054
R1595 CSoutput.n268 CSoutput.n267 0.00340054
R1596 CSoutput.n248 CSoutput.n247 0.00340054
R1597 CSoutput.n250 CSoutput.n249 0.00340054
R1598 CSoutput.n164 CSoutput.n154 0.00340054
R1599 CSoutput.n157 CSoutput.n155 0.00340054
R1600 CSoutput.n286 CSoutput.n285 0.00340054
R1601 CSoutput.n281 CSoutput.n150 0.00340054
R1602 CSoutput.n166 CSoutput.n151 0.00340054
R1603 CSoutput.n169 CSoutput.n153 0.00340054
R1604 CSoutput.n199 CSoutput.n193 0.00252698
R1605 CSoutput.n192 CSoutput.n190 0.00252698
R1606 CSoutput.n274 CSoutput.n273 0.00252698
R1607 CSoutput.n202 CSoutput.n200 0.00252698
R1608 CSoutput.n205 CSoutput.n203 0.00252698
R1609 CSoutput.n278 CSoutput.n173 0.00252698
R1610 CSoutput.n199 CSoutput.n198 0.00252698
R1611 CSoutput.n192 CSoutput.n191 0.00252698
R1612 CSoutput.n275 CSoutput.n274 0.00252698
R1613 CSoutput.n202 CSoutput.n201 0.00252698
R1614 CSoutput.n205 CSoutput.n204 0.00252698
R1615 CSoutput.n186 CSoutput.n173 0.00252698
R1616 CSoutput.n253 CSoutput.n223 0.00252698
R1617 CSoutput.n252 CSoutput.n222 0.00252698
R1618 CSoutput.n251 CSoutput.n207 0.00252698
R1619 CSoutput.n248 CSoutput.n218 0.00252698
R1620 CSoutput.n255 CSoutput.n250 0.00252698
R1621 CSoutput.n264 CSoutput.n257 0.00252698
R1622 CSoutput.n253 CSoutput.n242 0.00252698
R1623 CSoutput.n252 CSoutput.n244 0.00252698
R1624 CSoutput.n251 CSoutput.n246 0.00252698
R1625 CSoutput.n266 CSoutput.n218 0.00252698
R1626 CSoutput.n255 CSoutput.n220 0.00252698
R1627 CSoutput.n257 CSoutput.n219 0.00252698
R1628 CSoutput.n165 CSoutput.n159 0.00252698
R1629 CSoutput.n158 CSoutput.n156 0.00252698
R1630 CSoutput.n284 CSoutput.n283 0.00252698
R1631 CSoutput.n168 CSoutput.n166 0.00252698
R1632 CSoutput.n171 CSoutput.n169 0.00252698
R1633 CSoutput.n288 CSoutput.n139 0.00252698
R1634 CSoutput.n165 CSoutput.n164 0.00252698
R1635 CSoutput.n158 CSoutput.n157 0.00252698
R1636 CSoutput.n285 CSoutput.n284 0.00252698
R1637 CSoutput.n168 CSoutput.n167 0.00252698
R1638 CSoutput.n171 CSoutput.n170 0.00252698
R1639 CSoutput.n152 CSoutput.n139 0.00252698
R1640 CSoutput.n273 CSoutput.n272 0.0020275
R1641 CSoutput.n272 CSoutput.n271 0.0020275
R1642 CSoutput.n269 CSoutput.n207 0.0020275
R1643 CSoutput.n269 CSoutput.n268 0.0020275
R1644 CSoutput.n283 CSoutput.n282 0.0020275
R1645 CSoutput.n282 CSoutput.n281 0.0020275
R1646 CSoutput.n183 CSoutput.n182 0.00166668
R1647 CSoutput.n265 CSoutput.n221 0.00166668
R1648 CSoutput.n149 CSoutput.n148 0.00166668
R1649 CSoutput.n287 CSoutput.n149 0.00133328
R1650 CSoutput.n221 CSoutput.n217 0.00133328
R1651 CSoutput.n277 CSoutput.n183 0.00133328
R1652 CSoutput.n280 CSoutput.n172 0.001
R1653 CSoutput.n258 CSoutput.n172 0.001
R1654 CSoutput.n160 CSoutput.n140 0.001
R1655 CSoutput.n259 CSoutput.n140 0.001
R1656 CSoutput.n161 CSoutput.n141 0.001
R1657 CSoutput.n260 CSoutput.n141 0.001
R1658 CSoutput.n162 CSoutput.n142 0.001
R1659 CSoutput.n261 CSoutput.n142 0.001
R1660 CSoutput.n163 CSoutput.n143 0.001
R1661 CSoutput.n262 CSoutput.n143 0.001
R1662 CSoutput.n256 CSoutput.n208 0.001
R1663 CSoutput.n256 CSoutput.n254 0.001
R1664 CSoutput.n238 CSoutput.n209 0.001
R1665 CSoutput.n232 CSoutput.n209 0.001
R1666 CSoutput.n239 CSoutput.n210 0.001
R1667 CSoutput.n233 CSoutput.n210 0.001
R1668 CSoutput.n240 CSoutput.n211 0.001
R1669 CSoutput.n234 CSoutput.n211 0.001
R1670 CSoutput.n241 CSoutput.n212 0.001
R1671 CSoutput.n235 CSoutput.n212 0.001
R1672 CSoutput.n270 CSoutput.n206 0.001
R1673 CSoutput.n224 CSoutput.n206 0.001
R1674 CSoutput.n194 CSoutput.n174 0.001
R1675 CSoutput.n225 CSoutput.n174 0.001
R1676 CSoutput.n195 CSoutput.n175 0.001
R1677 CSoutput.n226 CSoutput.n175 0.001
R1678 CSoutput.n196 CSoutput.n176 0.001
R1679 CSoutput.n227 CSoutput.n176 0.001
R1680 CSoutput.n197 CSoutput.n177 0.001
R1681 CSoutput.n228 CSoutput.n177 0.001
R1682 CSoutput.n228 CSoutput.n178 0.001
R1683 CSoutput.n227 CSoutput.n179 0.001
R1684 CSoutput.n226 CSoutput.n180 0.001
R1685 CSoutput.n225 CSoutput.t171 0.001
R1686 CSoutput.n224 CSoutput.n181 0.001
R1687 CSoutput.n197 CSoutput.n179 0.001
R1688 CSoutput.n196 CSoutput.n180 0.001
R1689 CSoutput.n195 CSoutput.t171 0.001
R1690 CSoutput.n194 CSoutput.n181 0.001
R1691 CSoutput.n270 CSoutput.n182 0.001
R1692 CSoutput.n235 CSoutput.n213 0.001
R1693 CSoutput.n234 CSoutput.n214 0.001
R1694 CSoutput.n233 CSoutput.n215 0.001
R1695 CSoutput.n232 CSoutput.t178 0.001
R1696 CSoutput.n254 CSoutput.n216 0.001
R1697 CSoutput.n241 CSoutput.n214 0.001
R1698 CSoutput.n240 CSoutput.n215 0.001
R1699 CSoutput.n239 CSoutput.t178 0.001
R1700 CSoutput.n238 CSoutput.n216 0.001
R1701 CSoutput.n265 CSoutput.n208 0.001
R1702 CSoutput.n262 CSoutput.n144 0.001
R1703 CSoutput.n261 CSoutput.n145 0.001
R1704 CSoutput.n260 CSoutput.n146 0.001
R1705 CSoutput.n259 CSoutput.t185 0.001
R1706 CSoutput.n258 CSoutput.n147 0.001
R1707 CSoutput.n163 CSoutput.n145 0.001
R1708 CSoutput.n162 CSoutput.n146 0.001
R1709 CSoutput.n161 CSoutput.t185 0.001
R1710 CSoutput.n160 CSoutput.n147 0.001
R1711 CSoutput.n280 CSoutput.n148 0.001
R1712 gnd.n6795 gnd.n6794 1810.87
R1713 gnd.n4741 gnd.n4740 927.927
R1714 gnd.n7178 gnd.n84 838.452
R1715 gnd.n7327 gnd.n80 838.452
R1716 gnd.n1728 gnd.n1461 838.452
R1717 gnd.n1649 gnd.n1463 838.452
R1718 gnd.n4507 gnd.n1330 838.452
R1719 gnd.n3079 gnd.n1328 838.452
R1720 gnd.n1120 gnd.n1068 838.452
R1721 gnd.n4634 gnd.n1122 838.452
R1722 gnd.n7325 gnd.n86 819.232
R1723 gnd.n155 gnd.n82 819.232
R1724 gnd.n1913 gnd.n1460 819.232
R1725 gnd.n4360 gnd.n1464 819.232
R1726 gnd.n4509 gnd.n1325 819.232
R1727 gnd.n3246 gnd.n1327 819.232
R1728 gnd.n4637 gnd.n4636 819.232
R1729 gnd.n4713 gnd.n1072 819.232
R1730 gnd.n3125 gnd.n1335 771.183
R1731 gnd.n4378 gnd.n1438 771.183
R1732 gnd.n3008 gnd.n2517 771.183
R1733 gnd.n4124 gnd.n1440 771.183
R1734 gnd.n6057 gnd.n1013 766.379
R1735 gnd.n5973 gnd.n1015 766.379
R1736 gnd.n5268 gnd.n5171 766.379
R1737 gnd.n5264 gnd.n5169 766.379
R1738 gnd.n6054 gnd.n4743 756.769
R1739 gnd.n6023 gnd.n1016 756.769
R1740 gnd.n5361 gnd.n5078 756.769
R1741 gnd.n5359 gnd.n5081 756.769
R1742 gnd.n6275 gnd.n762 737.549
R1743 gnd.n6796 gnd.n451 737.549
R1744 gnd.n7006 gnd.n321 737.549
R1745 gnd.n4738 gnd.n930 737.549
R1746 gnd.n765 gnd.n762 585
R1747 gnd.n6273 gnd.n762 585
R1748 gnd.n6271 gnd.n6270 585
R1749 gnd.n6272 gnd.n6271 585
R1750 gnd.n6269 gnd.n764 585
R1751 gnd.n764 gnd.n763 585
R1752 gnd.n6268 gnd.n6267 585
R1753 gnd.n6267 gnd.n6266 585
R1754 gnd.n770 gnd.n769 585
R1755 gnd.n6265 gnd.n770 585
R1756 gnd.n6263 gnd.n6262 585
R1757 gnd.n6264 gnd.n6263 585
R1758 gnd.n6261 gnd.n772 585
R1759 gnd.n772 gnd.n771 585
R1760 gnd.n6260 gnd.n6259 585
R1761 gnd.n6259 gnd.n6258 585
R1762 gnd.n778 gnd.n777 585
R1763 gnd.n6257 gnd.n778 585
R1764 gnd.n6255 gnd.n6254 585
R1765 gnd.n6256 gnd.n6255 585
R1766 gnd.n6253 gnd.n780 585
R1767 gnd.n780 gnd.n779 585
R1768 gnd.n6252 gnd.n6251 585
R1769 gnd.n6251 gnd.n6250 585
R1770 gnd.n786 gnd.n785 585
R1771 gnd.n6249 gnd.n786 585
R1772 gnd.n6247 gnd.n6246 585
R1773 gnd.n6248 gnd.n6247 585
R1774 gnd.n6245 gnd.n788 585
R1775 gnd.n788 gnd.n787 585
R1776 gnd.n6244 gnd.n6243 585
R1777 gnd.n6243 gnd.n6242 585
R1778 gnd.n794 gnd.n793 585
R1779 gnd.n6241 gnd.n794 585
R1780 gnd.n6239 gnd.n6238 585
R1781 gnd.n6240 gnd.n6239 585
R1782 gnd.n6237 gnd.n796 585
R1783 gnd.n796 gnd.n795 585
R1784 gnd.n6236 gnd.n6235 585
R1785 gnd.n6235 gnd.n6234 585
R1786 gnd.n802 gnd.n801 585
R1787 gnd.n6233 gnd.n802 585
R1788 gnd.n6231 gnd.n6230 585
R1789 gnd.n6232 gnd.n6231 585
R1790 gnd.n6229 gnd.n804 585
R1791 gnd.n804 gnd.n803 585
R1792 gnd.n6228 gnd.n6227 585
R1793 gnd.n6227 gnd.n6226 585
R1794 gnd.n810 gnd.n809 585
R1795 gnd.n6225 gnd.n810 585
R1796 gnd.n6223 gnd.n6222 585
R1797 gnd.n6224 gnd.n6223 585
R1798 gnd.n6221 gnd.n812 585
R1799 gnd.n812 gnd.n811 585
R1800 gnd.n6220 gnd.n6219 585
R1801 gnd.n6219 gnd.n6218 585
R1802 gnd.n818 gnd.n817 585
R1803 gnd.n6217 gnd.n818 585
R1804 gnd.n6215 gnd.n6214 585
R1805 gnd.n6216 gnd.n6215 585
R1806 gnd.n6213 gnd.n820 585
R1807 gnd.n820 gnd.n819 585
R1808 gnd.n6212 gnd.n6211 585
R1809 gnd.n6211 gnd.n6210 585
R1810 gnd.n826 gnd.n825 585
R1811 gnd.n6209 gnd.n826 585
R1812 gnd.n6207 gnd.n6206 585
R1813 gnd.n6208 gnd.n6207 585
R1814 gnd.n6205 gnd.n828 585
R1815 gnd.n828 gnd.n827 585
R1816 gnd.n6204 gnd.n6203 585
R1817 gnd.n6203 gnd.n6202 585
R1818 gnd.n834 gnd.n833 585
R1819 gnd.n6201 gnd.n834 585
R1820 gnd.n6199 gnd.n6198 585
R1821 gnd.n6200 gnd.n6199 585
R1822 gnd.n6197 gnd.n836 585
R1823 gnd.n836 gnd.n835 585
R1824 gnd.n6196 gnd.n6195 585
R1825 gnd.n6195 gnd.n6194 585
R1826 gnd.n842 gnd.n841 585
R1827 gnd.n6193 gnd.n842 585
R1828 gnd.n6191 gnd.n6190 585
R1829 gnd.n6192 gnd.n6191 585
R1830 gnd.n6189 gnd.n844 585
R1831 gnd.n844 gnd.n843 585
R1832 gnd.n6188 gnd.n6187 585
R1833 gnd.n6187 gnd.n6186 585
R1834 gnd.n850 gnd.n849 585
R1835 gnd.n6185 gnd.n850 585
R1836 gnd.n6183 gnd.n6182 585
R1837 gnd.n6184 gnd.n6183 585
R1838 gnd.n6181 gnd.n852 585
R1839 gnd.n852 gnd.n851 585
R1840 gnd.n6180 gnd.n6179 585
R1841 gnd.n6179 gnd.n6178 585
R1842 gnd.n858 gnd.n857 585
R1843 gnd.n6177 gnd.n858 585
R1844 gnd.n6175 gnd.n6174 585
R1845 gnd.n6176 gnd.n6175 585
R1846 gnd.n6173 gnd.n860 585
R1847 gnd.n860 gnd.n859 585
R1848 gnd.n6172 gnd.n6171 585
R1849 gnd.n6171 gnd.n6170 585
R1850 gnd.n866 gnd.n865 585
R1851 gnd.n6169 gnd.n866 585
R1852 gnd.n6167 gnd.n6166 585
R1853 gnd.n6168 gnd.n6167 585
R1854 gnd.n6165 gnd.n868 585
R1855 gnd.n868 gnd.n867 585
R1856 gnd.n6164 gnd.n6163 585
R1857 gnd.n6163 gnd.n6162 585
R1858 gnd.n874 gnd.n873 585
R1859 gnd.n6161 gnd.n874 585
R1860 gnd.n6159 gnd.n6158 585
R1861 gnd.n6160 gnd.n6159 585
R1862 gnd.n6157 gnd.n876 585
R1863 gnd.n876 gnd.n875 585
R1864 gnd.n6156 gnd.n6155 585
R1865 gnd.n6155 gnd.n6154 585
R1866 gnd.n882 gnd.n881 585
R1867 gnd.n6153 gnd.n882 585
R1868 gnd.n6151 gnd.n6150 585
R1869 gnd.n6152 gnd.n6151 585
R1870 gnd.n6149 gnd.n884 585
R1871 gnd.n884 gnd.n883 585
R1872 gnd.n6148 gnd.n6147 585
R1873 gnd.n6147 gnd.n6146 585
R1874 gnd.n890 gnd.n889 585
R1875 gnd.n6145 gnd.n890 585
R1876 gnd.n6143 gnd.n6142 585
R1877 gnd.n6144 gnd.n6143 585
R1878 gnd.n6141 gnd.n892 585
R1879 gnd.n892 gnd.n891 585
R1880 gnd.n6140 gnd.n6139 585
R1881 gnd.n6139 gnd.n6138 585
R1882 gnd.n898 gnd.n897 585
R1883 gnd.n6137 gnd.n898 585
R1884 gnd.n6135 gnd.n6134 585
R1885 gnd.n6136 gnd.n6135 585
R1886 gnd.n6133 gnd.n900 585
R1887 gnd.n900 gnd.n899 585
R1888 gnd.n6132 gnd.n6131 585
R1889 gnd.n6131 gnd.n6130 585
R1890 gnd.n906 gnd.n905 585
R1891 gnd.n6129 gnd.n906 585
R1892 gnd.n6127 gnd.n6126 585
R1893 gnd.n6128 gnd.n6127 585
R1894 gnd.n6125 gnd.n908 585
R1895 gnd.n908 gnd.n907 585
R1896 gnd.n6124 gnd.n6123 585
R1897 gnd.n6123 gnd.n6122 585
R1898 gnd.n914 gnd.n913 585
R1899 gnd.n6121 gnd.n914 585
R1900 gnd.n6119 gnd.n6118 585
R1901 gnd.n6120 gnd.n6119 585
R1902 gnd.n6117 gnd.n916 585
R1903 gnd.n916 gnd.n915 585
R1904 gnd.n6116 gnd.n6115 585
R1905 gnd.n6115 gnd.n6114 585
R1906 gnd.n922 gnd.n921 585
R1907 gnd.n6113 gnd.n922 585
R1908 gnd.n6111 gnd.n6110 585
R1909 gnd.n6112 gnd.n6111 585
R1910 gnd.n6109 gnd.n924 585
R1911 gnd.n924 gnd.n923 585
R1912 gnd.n6108 gnd.n6107 585
R1913 gnd.n6107 gnd.n6106 585
R1914 gnd.n6276 gnd.n6275 585
R1915 gnd.n6275 gnd.n6274 585
R1916 gnd.n760 gnd.n759 585
R1917 gnd.n759 gnd.n758 585
R1918 gnd.n6281 gnd.n6280 585
R1919 gnd.n6282 gnd.n6281 585
R1920 gnd.n757 gnd.n756 585
R1921 gnd.n6283 gnd.n757 585
R1922 gnd.n6286 gnd.n6285 585
R1923 gnd.n6285 gnd.n6284 585
R1924 gnd.n754 gnd.n753 585
R1925 gnd.n753 gnd.n752 585
R1926 gnd.n6291 gnd.n6290 585
R1927 gnd.n6292 gnd.n6291 585
R1928 gnd.n751 gnd.n750 585
R1929 gnd.n6293 gnd.n751 585
R1930 gnd.n6296 gnd.n6295 585
R1931 gnd.n6295 gnd.n6294 585
R1932 gnd.n748 gnd.n747 585
R1933 gnd.n747 gnd.n746 585
R1934 gnd.n6301 gnd.n6300 585
R1935 gnd.n6302 gnd.n6301 585
R1936 gnd.n745 gnd.n744 585
R1937 gnd.n6303 gnd.n745 585
R1938 gnd.n6306 gnd.n6305 585
R1939 gnd.n6305 gnd.n6304 585
R1940 gnd.n742 gnd.n741 585
R1941 gnd.n741 gnd.n740 585
R1942 gnd.n6311 gnd.n6310 585
R1943 gnd.n6312 gnd.n6311 585
R1944 gnd.n739 gnd.n738 585
R1945 gnd.n6313 gnd.n739 585
R1946 gnd.n6316 gnd.n6315 585
R1947 gnd.n6315 gnd.n6314 585
R1948 gnd.n736 gnd.n735 585
R1949 gnd.n735 gnd.n734 585
R1950 gnd.n6321 gnd.n6320 585
R1951 gnd.n6322 gnd.n6321 585
R1952 gnd.n733 gnd.n732 585
R1953 gnd.n6323 gnd.n733 585
R1954 gnd.n6326 gnd.n6325 585
R1955 gnd.n6325 gnd.n6324 585
R1956 gnd.n730 gnd.n729 585
R1957 gnd.n729 gnd.n728 585
R1958 gnd.n6331 gnd.n6330 585
R1959 gnd.n6332 gnd.n6331 585
R1960 gnd.n727 gnd.n726 585
R1961 gnd.n6333 gnd.n727 585
R1962 gnd.n6336 gnd.n6335 585
R1963 gnd.n6335 gnd.n6334 585
R1964 gnd.n724 gnd.n723 585
R1965 gnd.n723 gnd.n722 585
R1966 gnd.n6341 gnd.n6340 585
R1967 gnd.n6342 gnd.n6341 585
R1968 gnd.n721 gnd.n720 585
R1969 gnd.n6343 gnd.n721 585
R1970 gnd.n6346 gnd.n6345 585
R1971 gnd.n6345 gnd.n6344 585
R1972 gnd.n718 gnd.n717 585
R1973 gnd.n717 gnd.n716 585
R1974 gnd.n6351 gnd.n6350 585
R1975 gnd.n6352 gnd.n6351 585
R1976 gnd.n715 gnd.n714 585
R1977 gnd.n6353 gnd.n715 585
R1978 gnd.n6356 gnd.n6355 585
R1979 gnd.n6355 gnd.n6354 585
R1980 gnd.n712 gnd.n711 585
R1981 gnd.n711 gnd.n710 585
R1982 gnd.n6361 gnd.n6360 585
R1983 gnd.n6362 gnd.n6361 585
R1984 gnd.n709 gnd.n708 585
R1985 gnd.n6363 gnd.n709 585
R1986 gnd.n6366 gnd.n6365 585
R1987 gnd.n6365 gnd.n6364 585
R1988 gnd.n706 gnd.n705 585
R1989 gnd.n705 gnd.n704 585
R1990 gnd.n6371 gnd.n6370 585
R1991 gnd.n6372 gnd.n6371 585
R1992 gnd.n703 gnd.n702 585
R1993 gnd.n6373 gnd.n703 585
R1994 gnd.n6376 gnd.n6375 585
R1995 gnd.n6375 gnd.n6374 585
R1996 gnd.n700 gnd.n699 585
R1997 gnd.n699 gnd.n698 585
R1998 gnd.n6381 gnd.n6380 585
R1999 gnd.n6382 gnd.n6381 585
R2000 gnd.n697 gnd.n696 585
R2001 gnd.n6383 gnd.n697 585
R2002 gnd.n6386 gnd.n6385 585
R2003 gnd.n6385 gnd.n6384 585
R2004 gnd.n694 gnd.n693 585
R2005 gnd.n693 gnd.n692 585
R2006 gnd.n6391 gnd.n6390 585
R2007 gnd.n6392 gnd.n6391 585
R2008 gnd.n691 gnd.n690 585
R2009 gnd.n6393 gnd.n691 585
R2010 gnd.n6396 gnd.n6395 585
R2011 gnd.n6395 gnd.n6394 585
R2012 gnd.n688 gnd.n687 585
R2013 gnd.n687 gnd.n686 585
R2014 gnd.n6401 gnd.n6400 585
R2015 gnd.n6402 gnd.n6401 585
R2016 gnd.n685 gnd.n684 585
R2017 gnd.n6403 gnd.n685 585
R2018 gnd.n6406 gnd.n6405 585
R2019 gnd.n6405 gnd.n6404 585
R2020 gnd.n682 gnd.n681 585
R2021 gnd.n681 gnd.n680 585
R2022 gnd.n6411 gnd.n6410 585
R2023 gnd.n6412 gnd.n6411 585
R2024 gnd.n679 gnd.n678 585
R2025 gnd.n6413 gnd.n679 585
R2026 gnd.n6416 gnd.n6415 585
R2027 gnd.n6415 gnd.n6414 585
R2028 gnd.n676 gnd.n675 585
R2029 gnd.n675 gnd.n674 585
R2030 gnd.n6421 gnd.n6420 585
R2031 gnd.n6422 gnd.n6421 585
R2032 gnd.n673 gnd.n672 585
R2033 gnd.n6423 gnd.n673 585
R2034 gnd.n6426 gnd.n6425 585
R2035 gnd.n6425 gnd.n6424 585
R2036 gnd.n670 gnd.n669 585
R2037 gnd.n669 gnd.n668 585
R2038 gnd.n6431 gnd.n6430 585
R2039 gnd.n6432 gnd.n6431 585
R2040 gnd.n667 gnd.n666 585
R2041 gnd.n6433 gnd.n667 585
R2042 gnd.n6436 gnd.n6435 585
R2043 gnd.n6435 gnd.n6434 585
R2044 gnd.n664 gnd.n663 585
R2045 gnd.n663 gnd.n662 585
R2046 gnd.n6441 gnd.n6440 585
R2047 gnd.n6442 gnd.n6441 585
R2048 gnd.n661 gnd.n660 585
R2049 gnd.n6443 gnd.n661 585
R2050 gnd.n6446 gnd.n6445 585
R2051 gnd.n6445 gnd.n6444 585
R2052 gnd.n658 gnd.n657 585
R2053 gnd.n657 gnd.n656 585
R2054 gnd.n6451 gnd.n6450 585
R2055 gnd.n6452 gnd.n6451 585
R2056 gnd.n655 gnd.n654 585
R2057 gnd.n6453 gnd.n655 585
R2058 gnd.n6456 gnd.n6455 585
R2059 gnd.n6455 gnd.n6454 585
R2060 gnd.n652 gnd.n651 585
R2061 gnd.n651 gnd.n650 585
R2062 gnd.n6461 gnd.n6460 585
R2063 gnd.n6462 gnd.n6461 585
R2064 gnd.n649 gnd.n648 585
R2065 gnd.n6463 gnd.n649 585
R2066 gnd.n6466 gnd.n6465 585
R2067 gnd.n6465 gnd.n6464 585
R2068 gnd.n646 gnd.n645 585
R2069 gnd.n645 gnd.n644 585
R2070 gnd.n6471 gnd.n6470 585
R2071 gnd.n6472 gnd.n6471 585
R2072 gnd.n643 gnd.n642 585
R2073 gnd.n6473 gnd.n643 585
R2074 gnd.n6476 gnd.n6475 585
R2075 gnd.n6475 gnd.n6474 585
R2076 gnd.n640 gnd.n639 585
R2077 gnd.n639 gnd.n638 585
R2078 gnd.n6481 gnd.n6480 585
R2079 gnd.n6482 gnd.n6481 585
R2080 gnd.n637 gnd.n636 585
R2081 gnd.n6483 gnd.n637 585
R2082 gnd.n6486 gnd.n6485 585
R2083 gnd.n6485 gnd.n6484 585
R2084 gnd.n634 gnd.n633 585
R2085 gnd.n633 gnd.n632 585
R2086 gnd.n6491 gnd.n6490 585
R2087 gnd.n6492 gnd.n6491 585
R2088 gnd.n631 gnd.n630 585
R2089 gnd.n6493 gnd.n631 585
R2090 gnd.n6496 gnd.n6495 585
R2091 gnd.n6495 gnd.n6494 585
R2092 gnd.n628 gnd.n627 585
R2093 gnd.n627 gnd.n626 585
R2094 gnd.n6501 gnd.n6500 585
R2095 gnd.n6502 gnd.n6501 585
R2096 gnd.n625 gnd.n624 585
R2097 gnd.n6503 gnd.n625 585
R2098 gnd.n6506 gnd.n6505 585
R2099 gnd.n6505 gnd.n6504 585
R2100 gnd.n622 gnd.n621 585
R2101 gnd.n621 gnd.n620 585
R2102 gnd.n6511 gnd.n6510 585
R2103 gnd.n6512 gnd.n6511 585
R2104 gnd.n619 gnd.n618 585
R2105 gnd.n6513 gnd.n619 585
R2106 gnd.n6516 gnd.n6515 585
R2107 gnd.n6515 gnd.n6514 585
R2108 gnd.n616 gnd.n615 585
R2109 gnd.n615 gnd.n614 585
R2110 gnd.n6521 gnd.n6520 585
R2111 gnd.n6522 gnd.n6521 585
R2112 gnd.n613 gnd.n612 585
R2113 gnd.n6523 gnd.n613 585
R2114 gnd.n6526 gnd.n6525 585
R2115 gnd.n6525 gnd.n6524 585
R2116 gnd.n610 gnd.n609 585
R2117 gnd.n609 gnd.n608 585
R2118 gnd.n6531 gnd.n6530 585
R2119 gnd.n6532 gnd.n6531 585
R2120 gnd.n607 gnd.n606 585
R2121 gnd.n6533 gnd.n607 585
R2122 gnd.n6536 gnd.n6535 585
R2123 gnd.n6535 gnd.n6534 585
R2124 gnd.n604 gnd.n603 585
R2125 gnd.n603 gnd.n602 585
R2126 gnd.n6541 gnd.n6540 585
R2127 gnd.n6542 gnd.n6541 585
R2128 gnd.n601 gnd.n600 585
R2129 gnd.n6543 gnd.n601 585
R2130 gnd.n6546 gnd.n6545 585
R2131 gnd.n6545 gnd.n6544 585
R2132 gnd.n598 gnd.n597 585
R2133 gnd.n597 gnd.n596 585
R2134 gnd.n6551 gnd.n6550 585
R2135 gnd.n6552 gnd.n6551 585
R2136 gnd.n595 gnd.n594 585
R2137 gnd.n6553 gnd.n595 585
R2138 gnd.n6556 gnd.n6555 585
R2139 gnd.n6555 gnd.n6554 585
R2140 gnd.n592 gnd.n591 585
R2141 gnd.n591 gnd.n590 585
R2142 gnd.n6561 gnd.n6560 585
R2143 gnd.n6562 gnd.n6561 585
R2144 gnd.n589 gnd.n588 585
R2145 gnd.n6563 gnd.n589 585
R2146 gnd.n6566 gnd.n6565 585
R2147 gnd.n6565 gnd.n6564 585
R2148 gnd.n586 gnd.n585 585
R2149 gnd.n585 gnd.n584 585
R2150 gnd.n6571 gnd.n6570 585
R2151 gnd.n6572 gnd.n6571 585
R2152 gnd.n583 gnd.n582 585
R2153 gnd.n6573 gnd.n583 585
R2154 gnd.n6576 gnd.n6575 585
R2155 gnd.n6575 gnd.n6574 585
R2156 gnd.n580 gnd.n579 585
R2157 gnd.n579 gnd.n578 585
R2158 gnd.n6581 gnd.n6580 585
R2159 gnd.n6582 gnd.n6581 585
R2160 gnd.n577 gnd.n576 585
R2161 gnd.n6583 gnd.n577 585
R2162 gnd.n6586 gnd.n6585 585
R2163 gnd.n6585 gnd.n6584 585
R2164 gnd.n574 gnd.n573 585
R2165 gnd.n573 gnd.n572 585
R2166 gnd.n6591 gnd.n6590 585
R2167 gnd.n6592 gnd.n6591 585
R2168 gnd.n571 gnd.n570 585
R2169 gnd.n6593 gnd.n571 585
R2170 gnd.n6596 gnd.n6595 585
R2171 gnd.n6595 gnd.n6594 585
R2172 gnd.n568 gnd.n567 585
R2173 gnd.n567 gnd.n566 585
R2174 gnd.n6601 gnd.n6600 585
R2175 gnd.n6602 gnd.n6601 585
R2176 gnd.n565 gnd.n564 585
R2177 gnd.n6603 gnd.n565 585
R2178 gnd.n6606 gnd.n6605 585
R2179 gnd.n6605 gnd.n6604 585
R2180 gnd.n562 gnd.n561 585
R2181 gnd.n561 gnd.n560 585
R2182 gnd.n6611 gnd.n6610 585
R2183 gnd.n6612 gnd.n6611 585
R2184 gnd.n559 gnd.n558 585
R2185 gnd.n6613 gnd.n559 585
R2186 gnd.n6616 gnd.n6615 585
R2187 gnd.n6615 gnd.n6614 585
R2188 gnd.n556 gnd.n555 585
R2189 gnd.n555 gnd.n554 585
R2190 gnd.n6621 gnd.n6620 585
R2191 gnd.n6622 gnd.n6621 585
R2192 gnd.n553 gnd.n552 585
R2193 gnd.n6623 gnd.n553 585
R2194 gnd.n6626 gnd.n6625 585
R2195 gnd.n6625 gnd.n6624 585
R2196 gnd.n550 gnd.n549 585
R2197 gnd.n549 gnd.n548 585
R2198 gnd.n6631 gnd.n6630 585
R2199 gnd.n6632 gnd.n6631 585
R2200 gnd.n547 gnd.n546 585
R2201 gnd.n6633 gnd.n547 585
R2202 gnd.n6636 gnd.n6635 585
R2203 gnd.n6635 gnd.n6634 585
R2204 gnd.n544 gnd.n543 585
R2205 gnd.n543 gnd.n542 585
R2206 gnd.n6641 gnd.n6640 585
R2207 gnd.n6642 gnd.n6641 585
R2208 gnd.n541 gnd.n540 585
R2209 gnd.n6643 gnd.n541 585
R2210 gnd.n6646 gnd.n6645 585
R2211 gnd.n6645 gnd.n6644 585
R2212 gnd.n538 gnd.n537 585
R2213 gnd.n537 gnd.n536 585
R2214 gnd.n6651 gnd.n6650 585
R2215 gnd.n6652 gnd.n6651 585
R2216 gnd.n535 gnd.n534 585
R2217 gnd.n6653 gnd.n535 585
R2218 gnd.n6656 gnd.n6655 585
R2219 gnd.n6655 gnd.n6654 585
R2220 gnd.n532 gnd.n531 585
R2221 gnd.n531 gnd.n530 585
R2222 gnd.n6661 gnd.n6660 585
R2223 gnd.n6662 gnd.n6661 585
R2224 gnd.n529 gnd.n528 585
R2225 gnd.n6663 gnd.n529 585
R2226 gnd.n6666 gnd.n6665 585
R2227 gnd.n6665 gnd.n6664 585
R2228 gnd.n526 gnd.n525 585
R2229 gnd.n525 gnd.n524 585
R2230 gnd.n6671 gnd.n6670 585
R2231 gnd.n6672 gnd.n6671 585
R2232 gnd.n523 gnd.n522 585
R2233 gnd.n6673 gnd.n523 585
R2234 gnd.n6676 gnd.n6675 585
R2235 gnd.n6675 gnd.n6674 585
R2236 gnd.n520 gnd.n519 585
R2237 gnd.n519 gnd.n518 585
R2238 gnd.n6681 gnd.n6680 585
R2239 gnd.n6682 gnd.n6681 585
R2240 gnd.n517 gnd.n516 585
R2241 gnd.n6683 gnd.n517 585
R2242 gnd.n6686 gnd.n6685 585
R2243 gnd.n6685 gnd.n6684 585
R2244 gnd.n514 gnd.n513 585
R2245 gnd.n513 gnd.n512 585
R2246 gnd.n6691 gnd.n6690 585
R2247 gnd.n6692 gnd.n6691 585
R2248 gnd.n511 gnd.n510 585
R2249 gnd.n6693 gnd.n511 585
R2250 gnd.n6696 gnd.n6695 585
R2251 gnd.n6695 gnd.n6694 585
R2252 gnd.n508 gnd.n507 585
R2253 gnd.n507 gnd.n506 585
R2254 gnd.n6701 gnd.n6700 585
R2255 gnd.n6702 gnd.n6701 585
R2256 gnd.n505 gnd.n504 585
R2257 gnd.n6703 gnd.n505 585
R2258 gnd.n6706 gnd.n6705 585
R2259 gnd.n6705 gnd.n6704 585
R2260 gnd.n502 gnd.n501 585
R2261 gnd.n501 gnd.n500 585
R2262 gnd.n6711 gnd.n6710 585
R2263 gnd.n6712 gnd.n6711 585
R2264 gnd.n499 gnd.n498 585
R2265 gnd.n6713 gnd.n499 585
R2266 gnd.n6716 gnd.n6715 585
R2267 gnd.n6715 gnd.n6714 585
R2268 gnd.n496 gnd.n495 585
R2269 gnd.n495 gnd.n494 585
R2270 gnd.n6721 gnd.n6720 585
R2271 gnd.n6722 gnd.n6721 585
R2272 gnd.n493 gnd.n492 585
R2273 gnd.n6723 gnd.n493 585
R2274 gnd.n6726 gnd.n6725 585
R2275 gnd.n6725 gnd.n6724 585
R2276 gnd.n490 gnd.n489 585
R2277 gnd.n489 gnd.n488 585
R2278 gnd.n6731 gnd.n6730 585
R2279 gnd.n6732 gnd.n6731 585
R2280 gnd.n487 gnd.n486 585
R2281 gnd.n6733 gnd.n487 585
R2282 gnd.n6736 gnd.n6735 585
R2283 gnd.n6735 gnd.n6734 585
R2284 gnd.n484 gnd.n483 585
R2285 gnd.n483 gnd.n482 585
R2286 gnd.n6741 gnd.n6740 585
R2287 gnd.n6742 gnd.n6741 585
R2288 gnd.n481 gnd.n480 585
R2289 gnd.n6743 gnd.n481 585
R2290 gnd.n6746 gnd.n6745 585
R2291 gnd.n6745 gnd.n6744 585
R2292 gnd.n478 gnd.n477 585
R2293 gnd.n477 gnd.n476 585
R2294 gnd.n6751 gnd.n6750 585
R2295 gnd.n6752 gnd.n6751 585
R2296 gnd.n475 gnd.n474 585
R2297 gnd.n6753 gnd.n475 585
R2298 gnd.n6756 gnd.n6755 585
R2299 gnd.n6755 gnd.n6754 585
R2300 gnd.n472 gnd.n471 585
R2301 gnd.n471 gnd.n470 585
R2302 gnd.n6761 gnd.n6760 585
R2303 gnd.n6762 gnd.n6761 585
R2304 gnd.n469 gnd.n468 585
R2305 gnd.n6763 gnd.n469 585
R2306 gnd.n6766 gnd.n6765 585
R2307 gnd.n6765 gnd.n6764 585
R2308 gnd.n466 gnd.n465 585
R2309 gnd.n465 gnd.n464 585
R2310 gnd.n6771 gnd.n6770 585
R2311 gnd.n6772 gnd.n6771 585
R2312 gnd.n463 gnd.n462 585
R2313 gnd.n6773 gnd.n463 585
R2314 gnd.n6776 gnd.n6775 585
R2315 gnd.n6775 gnd.n6774 585
R2316 gnd.n460 gnd.n459 585
R2317 gnd.n459 gnd.n458 585
R2318 gnd.n6781 gnd.n6780 585
R2319 gnd.n6782 gnd.n6781 585
R2320 gnd.n457 gnd.n456 585
R2321 gnd.n6783 gnd.n457 585
R2322 gnd.n6786 gnd.n6785 585
R2323 gnd.n6785 gnd.n6784 585
R2324 gnd.n454 gnd.n453 585
R2325 gnd.n453 gnd.n452 585
R2326 gnd.n6792 gnd.n6791 585
R2327 gnd.n6793 gnd.n6792 585
R2328 gnd.n6790 gnd.n451 585
R2329 gnd.n6794 gnd.n451 585
R2330 gnd.n326 gnd.n325 585
R2331 gnd.n7004 gnd.n326 585
R2332 gnd.n7002 gnd.n7001 585
R2333 gnd.n7003 gnd.n7002 585
R2334 gnd.n329 gnd.n328 585
R2335 gnd.n328 gnd.n327 585
R2336 gnd.n6997 gnd.n6996 585
R2337 gnd.n6996 gnd.n6995 585
R2338 gnd.n332 gnd.n331 585
R2339 gnd.n6994 gnd.n332 585
R2340 gnd.n6992 gnd.n6991 585
R2341 gnd.n6993 gnd.n6992 585
R2342 gnd.n335 gnd.n334 585
R2343 gnd.n334 gnd.n333 585
R2344 gnd.n6987 gnd.n6986 585
R2345 gnd.n6986 gnd.n6985 585
R2346 gnd.n338 gnd.n337 585
R2347 gnd.n6984 gnd.n338 585
R2348 gnd.n6982 gnd.n6981 585
R2349 gnd.n6983 gnd.n6982 585
R2350 gnd.n341 gnd.n340 585
R2351 gnd.n340 gnd.n339 585
R2352 gnd.n6977 gnd.n6976 585
R2353 gnd.n6976 gnd.n6975 585
R2354 gnd.n344 gnd.n343 585
R2355 gnd.n6974 gnd.n344 585
R2356 gnd.n6972 gnd.n6971 585
R2357 gnd.n6973 gnd.n6972 585
R2358 gnd.n347 gnd.n346 585
R2359 gnd.n346 gnd.n345 585
R2360 gnd.n6967 gnd.n6966 585
R2361 gnd.n6966 gnd.n6965 585
R2362 gnd.n350 gnd.n349 585
R2363 gnd.n6964 gnd.n350 585
R2364 gnd.n6962 gnd.n6961 585
R2365 gnd.n6963 gnd.n6962 585
R2366 gnd.n353 gnd.n352 585
R2367 gnd.n352 gnd.n351 585
R2368 gnd.n6957 gnd.n6956 585
R2369 gnd.n6956 gnd.n6955 585
R2370 gnd.n356 gnd.n355 585
R2371 gnd.n6954 gnd.n356 585
R2372 gnd.n6952 gnd.n6951 585
R2373 gnd.n6953 gnd.n6952 585
R2374 gnd.n359 gnd.n358 585
R2375 gnd.n358 gnd.n357 585
R2376 gnd.n6947 gnd.n6946 585
R2377 gnd.n6946 gnd.n6945 585
R2378 gnd.n362 gnd.n361 585
R2379 gnd.n6944 gnd.n362 585
R2380 gnd.n6942 gnd.n6941 585
R2381 gnd.n6943 gnd.n6942 585
R2382 gnd.n365 gnd.n364 585
R2383 gnd.n364 gnd.n363 585
R2384 gnd.n6937 gnd.n6936 585
R2385 gnd.n6936 gnd.n6935 585
R2386 gnd.n368 gnd.n367 585
R2387 gnd.n6934 gnd.n368 585
R2388 gnd.n6932 gnd.n6931 585
R2389 gnd.n6933 gnd.n6932 585
R2390 gnd.n371 gnd.n370 585
R2391 gnd.n370 gnd.n369 585
R2392 gnd.n6927 gnd.n6926 585
R2393 gnd.n6926 gnd.n6925 585
R2394 gnd.n374 gnd.n373 585
R2395 gnd.n6924 gnd.n374 585
R2396 gnd.n6922 gnd.n6921 585
R2397 gnd.n6923 gnd.n6922 585
R2398 gnd.n377 gnd.n376 585
R2399 gnd.n376 gnd.n375 585
R2400 gnd.n6917 gnd.n6916 585
R2401 gnd.n6916 gnd.n6915 585
R2402 gnd.n380 gnd.n379 585
R2403 gnd.n6914 gnd.n380 585
R2404 gnd.n6912 gnd.n6911 585
R2405 gnd.n6913 gnd.n6912 585
R2406 gnd.n383 gnd.n382 585
R2407 gnd.n382 gnd.n381 585
R2408 gnd.n6907 gnd.n6906 585
R2409 gnd.n6906 gnd.n6905 585
R2410 gnd.n386 gnd.n385 585
R2411 gnd.n6904 gnd.n386 585
R2412 gnd.n6902 gnd.n6901 585
R2413 gnd.n6903 gnd.n6902 585
R2414 gnd.n389 gnd.n388 585
R2415 gnd.n388 gnd.n387 585
R2416 gnd.n6897 gnd.n6896 585
R2417 gnd.n6896 gnd.n6895 585
R2418 gnd.n392 gnd.n391 585
R2419 gnd.n6894 gnd.n392 585
R2420 gnd.n6892 gnd.n6891 585
R2421 gnd.n6893 gnd.n6892 585
R2422 gnd.n395 gnd.n394 585
R2423 gnd.n394 gnd.n393 585
R2424 gnd.n6887 gnd.n6886 585
R2425 gnd.n6886 gnd.n6885 585
R2426 gnd.n398 gnd.n397 585
R2427 gnd.n6884 gnd.n398 585
R2428 gnd.n6882 gnd.n6881 585
R2429 gnd.n6883 gnd.n6882 585
R2430 gnd.n401 gnd.n400 585
R2431 gnd.n400 gnd.n399 585
R2432 gnd.n6877 gnd.n6876 585
R2433 gnd.n6876 gnd.n6875 585
R2434 gnd.n404 gnd.n403 585
R2435 gnd.n6874 gnd.n404 585
R2436 gnd.n6872 gnd.n6871 585
R2437 gnd.n6873 gnd.n6872 585
R2438 gnd.n407 gnd.n406 585
R2439 gnd.n406 gnd.n405 585
R2440 gnd.n6867 gnd.n6866 585
R2441 gnd.n6866 gnd.n6865 585
R2442 gnd.n410 gnd.n409 585
R2443 gnd.n6864 gnd.n410 585
R2444 gnd.n6862 gnd.n6861 585
R2445 gnd.n6863 gnd.n6862 585
R2446 gnd.n413 gnd.n412 585
R2447 gnd.n412 gnd.n411 585
R2448 gnd.n6857 gnd.n6856 585
R2449 gnd.n6856 gnd.n6855 585
R2450 gnd.n416 gnd.n415 585
R2451 gnd.n6854 gnd.n416 585
R2452 gnd.n6852 gnd.n6851 585
R2453 gnd.n6853 gnd.n6852 585
R2454 gnd.n419 gnd.n418 585
R2455 gnd.n418 gnd.n417 585
R2456 gnd.n6847 gnd.n6846 585
R2457 gnd.n6846 gnd.n6845 585
R2458 gnd.n422 gnd.n421 585
R2459 gnd.n6844 gnd.n422 585
R2460 gnd.n6842 gnd.n6841 585
R2461 gnd.n6843 gnd.n6842 585
R2462 gnd.n425 gnd.n424 585
R2463 gnd.n424 gnd.n423 585
R2464 gnd.n6837 gnd.n6836 585
R2465 gnd.n6836 gnd.n6835 585
R2466 gnd.n428 gnd.n427 585
R2467 gnd.n6834 gnd.n428 585
R2468 gnd.n6832 gnd.n6831 585
R2469 gnd.n6833 gnd.n6832 585
R2470 gnd.n431 gnd.n430 585
R2471 gnd.n430 gnd.n429 585
R2472 gnd.n6827 gnd.n6826 585
R2473 gnd.n6826 gnd.n6825 585
R2474 gnd.n434 gnd.n433 585
R2475 gnd.n6824 gnd.n434 585
R2476 gnd.n6822 gnd.n6821 585
R2477 gnd.n6823 gnd.n6822 585
R2478 gnd.n437 gnd.n436 585
R2479 gnd.n436 gnd.n435 585
R2480 gnd.n6817 gnd.n6816 585
R2481 gnd.n6816 gnd.n6815 585
R2482 gnd.n440 gnd.n439 585
R2483 gnd.n6814 gnd.n440 585
R2484 gnd.n6812 gnd.n6811 585
R2485 gnd.n6813 gnd.n6812 585
R2486 gnd.n443 gnd.n442 585
R2487 gnd.n442 gnd.n441 585
R2488 gnd.n6807 gnd.n6806 585
R2489 gnd.n6806 gnd.n6805 585
R2490 gnd.n446 gnd.n445 585
R2491 gnd.n6804 gnd.n446 585
R2492 gnd.n6802 gnd.n6801 585
R2493 gnd.n6803 gnd.n6802 585
R2494 gnd.n449 gnd.n448 585
R2495 gnd.n448 gnd.n447 585
R2496 gnd.n6797 gnd.n6796 585
R2497 gnd.n6796 gnd.n6795 585
R2498 gnd.n4507 gnd.n4506 585
R2499 gnd.n4508 gnd.n4507 585
R2500 gnd.n1315 gnd.n1314 585
R2501 gnd.n3239 gnd.n1315 585
R2502 gnd.n4516 gnd.n4515 585
R2503 gnd.n4515 gnd.n4514 585
R2504 gnd.n4517 gnd.n1309 585
R2505 gnd.n2943 gnd.n1309 585
R2506 gnd.n4519 gnd.n4518 585
R2507 gnd.n4520 gnd.n4519 585
R2508 gnd.n1294 gnd.n1293 585
R2509 gnd.n2934 gnd.n1294 585
R2510 gnd.n4528 gnd.n4527 585
R2511 gnd.n4527 gnd.n4526 585
R2512 gnd.n4529 gnd.n1288 585
R2513 gnd.n2930 gnd.n1288 585
R2514 gnd.n4531 gnd.n4530 585
R2515 gnd.n4532 gnd.n4531 585
R2516 gnd.n1272 gnd.n1271 585
R2517 gnd.n2923 gnd.n1272 585
R2518 gnd.n4540 gnd.n4539 585
R2519 gnd.n4539 gnd.n4538 585
R2520 gnd.n4541 gnd.n1266 585
R2521 gnd.n2960 gnd.n1266 585
R2522 gnd.n4543 gnd.n4542 585
R2523 gnd.n4544 gnd.n4543 585
R2524 gnd.n1252 gnd.n1251 585
R2525 gnd.n2915 gnd.n1252 585
R2526 gnd.n4552 gnd.n4551 585
R2527 gnd.n4551 gnd.n4550 585
R2528 gnd.n4553 gnd.n1246 585
R2529 gnd.n2907 gnd.n1246 585
R2530 gnd.n4555 gnd.n4554 585
R2531 gnd.n4556 gnd.n4555 585
R2532 gnd.n1233 gnd.n1232 585
R2533 gnd.n2868 gnd.n1233 585
R2534 gnd.n4565 gnd.n4564 585
R2535 gnd.n4564 gnd.n4563 585
R2536 gnd.n4566 gnd.n1228 585
R2537 gnd.n2876 gnd.n1228 585
R2538 gnd.n4568 gnd.n4567 585
R2539 gnd.n4569 gnd.n4568 585
R2540 gnd.n1217 gnd.n1216 585
R2541 gnd.n2854 gnd.n1217 585
R2542 gnd.n4578 gnd.n4577 585
R2543 gnd.n4577 gnd.n4576 585
R2544 gnd.n4579 gnd.n1209 585
R2545 gnd.n2887 gnd.n1209 585
R2546 gnd.n4581 gnd.n4580 585
R2547 gnd.n4582 gnd.n4581 585
R2548 gnd.n1210 gnd.n1208 585
R2549 gnd.n2893 gnd.n1208 585
R2550 gnd.n1193 gnd.n1192 585
R2551 gnd.n2611 gnd.n1193 585
R2552 gnd.n4592 gnd.n4591 585
R2553 gnd.n4591 gnd.n4590 585
R2554 gnd.n4593 gnd.n1187 585
R2555 gnd.n2837 gnd.n1187 585
R2556 gnd.n4595 gnd.n4594 585
R2557 gnd.n4596 gnd.n4595 585
R2558 gnd.n1171 gnd.n1170 585
R2559 gnd.n2825 gnd.n1171 585
R2560 gnd.n4604 gnd.n4603 585
R2561 gnd.n4603 gnd.n4602 585
R2562 gnd.n4605 gnd.n1165 585
R2563 gnd.n2816 gnd.n1165 585
R2564 gnd.n4607 gnd.n4606 585
R2565 gnd.n4608 gnd.n4607 585
R2566 gnd.n1151 gnd.n1150 585
R2567 gnd.n2808 gnd.n1151 585
R2568 gnd.n4616 gnd.n4615 585
R2569 gnd.n4615 gnd.n4614 585
R2570 gnd.n4617 gnd.n1146 585
R2571 gnd.n2800 gnd.n1146 585
R2572 gnd.n4619 gnd.n4618 585
R2573 gnd.n4620 gnd.n4619 585
R2574 gnd.n1129 gnd.n1127 585
R2575 gnd.n2747 gnd.n1129 585
R2576 gnd.n4628 gnd.n4627 585
R2577 gnd.n4627 gnd.n4626 585
R2578 gnd.n1128 gnd.n1125 585
R2579 gnd.n2753 gnd.n1128 585
R2580 gnd.n4632 gnd.n1123 585
R2581 gnd.n2667 gnd.n1123 585
R2582 gnd.n4634 gnd.n4633 585
R2583 gnd.n4635 gnd.n4634 585
R2584 gnd.n2686 gnd.n1122 585
R2585 gnd.n2688 gnd.n2687 585
R2586 gnd.n2690 gnd.n2689 585
R2587 gnd.n2694 gnd.n2683 585
R2588 gnd.n2696 gnd.n2695 585
R2589 gnd.n2698 gnd.n2697 585
R2590 gnd.n2700 gnd.n2699 585
R2591 gnd.n2704 gnd.n2681 585
R2592 gnd.n2706 gnd.n2705 585
R2593 gnd.n2708 gnd.n2707 585
R2594 gnd.n2710 gnd.n2709 585
R2595 gnd.n2714 gnd.n2679 585
R2596 gnd.n2716 gnd.n2715 585
R2597 gnd.n2718 gnd.n2717 585
R2598 gnd.n2720 gnd.n2719 585
R2599 gnd.n2676 gnd.n2675 585
R2600 gnd.n2724 gnd.n2677 585
R2601 gnd.n2725 gnd.n2672 585
R2602 gnd.n2726 gnd.n1068 585
R2603 gnd.n4715 gnd.n1068 585
R2604 gnd.n3080 gnd.n3079 585
R2605 gnd.n3077 gnd.n3071 585
R2606 gnd.n3087 gnd.n3068 585
R2607 gnd.n3088 gnd.n3066 585
R2608 gnd.n3065 gnd.n3058 585
R2609 gnd.n3095 gnd.n3057 585
R2610 gnd.n3096 gnd.n3056 585
R2611 gnd.n3054 gnd.n3046 585
R2612 gnd.n3103 gnd.n3045 585
R2613 gnd.n3104 gnd.n3043 585
R2614 gnd.n3042 gnd.n3035 585
R2615 gnd.n3111 gnd.n3034 585
R2616 gnd.n3112 gnd.n3033 585
R2617 gnd.n3031 gnd.n3024 585
R2618 gnd.n3119 gnd.n3023 585
R2619 gnd.n3120 gnd.n3021 585
R2620 gnd.n3020 gnd.n3016 585
R2621 gnd.n3018 gnd.n3017 585
R2622 gnd.n1332 gnd.n1330 585
R2623 gnd.n2459 gnd.n1330 585
R2624 gnd.n2495 gnd.n1328 585
R2625 gnd.n4508 gnd.n1328 585
R2626 gnd.n3238 gnd.n3237 585
R2627 gnd.n3239 gnd.n3238 585
R2628 gnd.n2494 gnd.n1318 585
R2629 gnd.n4514 gnd.n1318 585
R2630 gnd.n2946 gnd.n2944 585
R2631 gnd.n2944 gnd.n2943 585
R2632 gnd.n2947 gnd.n1307 585
R2633 gnd.n4520 gnd.n1307 585
R2634 gnd.n2948 gnd.n2586 585
R2635 gnd.n2934 gnd.n2586 585
R2636 gnd.n2584 gnd.n1296 585
R2637 gnd.n4526 gnd.n1296 585
R2638 gnd.n2952 gnd.n2583 585
R2639 gnd.n2930 gnd.n2583 585
R2640 gnd.n2953 gnd.n1286 585
R2641 gnd.n4532 gnd.n1286 585
R2642 gnd.n2954 gnd.n2582 585
R2643 gnd.n2923 gnd.n2582 585
R2644 gnd.n2579 gnd.n1275 585
R2645 gnd.n4538 gnd.n1275 585
R2646 gnd.n2959 gnd.n2958 585
R2647 gnd.n2960 gnd.n2959 585
R2648 gnd.n2578 gnd.n1265 585
R2649 gnd.n4544 gnd.n1265 585
R2650 gnd.n2914 gnd.n2913 585
R2651 gnd.n2915 gnd.n2914 585
R2652 gnd.n2594 gnd.n1254 585
R2653 gnd.n4550 gnd.n1254 585
R2654 gnd.n2909 gnd.n2908 585
R2655 gnd.n2908 gnd.n2907 585
R2656 gnd.n2596 gnd.n1244 585
R2657 gnd.n4556 gnd.n1244 585
R2658 gnd.n2870 gnd.n2869 585
R2659 gnd.n2869 gnd.n2868 585
R2660 gnd.n2631 gnd.n1236 585
R2661 gnd.n4563 gnd.n1236 585
R2662 gnd.n2875 gnd.n2874 585
R2663 gnd.n2876 gnd.n2875 585
R2664 gnd.n2630 gnd.n1227 585
R2665 gnd.n4569 gnd.n1227 585
R2666 gnd.n2853 gnd.n2852 585
R2667 gnd.n2854 gnd.n2853 585
R2668 gnd.n2618 gnd.n1219 585
R2669 gnd.n4576 gnd.n1219 585
R2670 gnd.n2889 gnd.n2888 585
R2671 gnd.n2888 gnd.n2887 585
R2672 gnd.n2890 gnd.n1206 585
R2673 gnd.n4582 gnd.n1206 585
R2674 gnd.n2892 gnd.n2891 585
R2675 gnd.n2893 gnd.n2892 585
R2676 gnd.n2614 gnd.n2613 585
R2677 gnd.n2613 gnd.n2611 585
R2678 gnd.n2833 gnd.n1195 585
R2679 gnd.n4590 gnd.n1195 585
R2680 gnd.n2835 gnd.n2834 585
R2681 gnd.n2837 gnd.n2835 585
R2682 gnd.n2642 gnd.n1185 585
R2683 gnd.n4596 gnd.n1185 585
R2684 gnd.n2827 gnd.n2826 585
R2685 gnd.n2826 gnd.n2825 585
R2686 gnd.n2644 gnd.n1174 585
R2687 gnd.n4602 gnd.n1174 585
R2688 gnd.n2815 gnd.n2814 585
R2689 gnd.n2816 gnd.n2815 585
R2690 gnd.n2649 gnd.n1164 585
R2691 gnd.n4608 gnd.n1164 585
R2692 gnd.n2810 gnd.n2809 585
R2693 gnd.n2809 gnd.n2808 585
R2694 gnd.n2651 gnd.n1153 585
R2695 gnd.n4614 gnd.n1153 585
R2696 gnd.n2736 gnd.n2655 585
R2697 gnd.n2800 gnd.n2655 585
R2698 gnd.n2737 gnd.n1144 585
R2699 gnd.n4620 gnd.n1144 585
R2700 gnd.n2749 gnd.n2748 585
R2701 gnd.n2748 gnd.n2747 585
R2702 gnd.n2750 gnd.n1132 585
R2703 gnd.n4626 gnd.n1132 585
R2704 gnd.n2752 gnd.n2751 585
R2705 gnd.n2753 gnd.n2752 585
R2706 gnd.n2670 gnd.n2669 585
R2707 gnd.n2669 gnd.n2667 585
R2708 gnd.n2728 gnd.n1120 585
R2709 gnd.n4635 gnd.n1120 585
R2710 gnd.n165 gnd.n84 585
R2711 gnd.n7326 gnd.n84 585
R2712 gnd.n7246 gnd.n7245 585
R2713 gnd.n7247 gnd.n7246 585
R2714 gnd.n164 gnd.n163 585
R2715 gnd.n173 gnd.n163 585
R2716 gnd.n7174 gnd.n7173 585
R2717 gnd.n7173 gnd.n7172 585
R2718 gnd.n168 gnd.n167 585
R2719 gnd.n7059 gnd.n168 585
R2720 gnd.n7161 gnd.n7160 585
R2721 gnd.n7162 gnd.n7161 585
R2722 gnd.n184 gnd.n183 585
R2723 gnd.n7065 gnd.n183 585
R2724 gnd.n7156 gnd.n7155 585
R2725 gnd.n7155 gnd.n7154 585
R2726 gnd.n187 gnd.n186 585
R2727 gnd.n7048 gnd.n187 585
R2728 gnd.n7145 gnd.n7144 585
R2729 gnd.n7146 gnd.n7145 585
R2730 gnd.n199 gnd.n198 585
R2731 gnd.n7074 gnd.n198 585
R2732 gnd.n7140 gnd.n7139 585
R2733 gnd.n7139 gnd.n7138 585
R2734 gnd.n202 gnd.n201 585
R2735 gnd.n7078 gnd.n202 585
R2736 gnd.n7129 gnd.n7128 585
R2737 gnd.n7130 gnd.n7129 585
R2738 gnd.n216 gnd.n215 585
R2739 gnd.n7084 gnd.n215 585
R2740 gnd.n7124 gnd.n7123 585
R2741 gnd.n7123 gnd.n7122 585
R2742 gnd.n219 gnd.n218 585
R2743 gnd.n4282 gnd.n219 585
R2744 gnd.n7100 gnd.n7099 585
R2745 gnd.n7099 gnd.n7098 585
R2746 gnd.n7101 gnd.n248 585
R2747 gnd.n7094 gnd.n248 585
R2748 gnd.n4289 gnd.n246 585
R2749 gnd.n4290 gnd.n4289 585
R2750 gnd.n7105 gnd.n245 585
R2751 gnd.n1518 gnd.n245 585
R2752 gnd.n7106 gnd.n244 585
R2753 gnd.n4309 gnd.n244 585
R2754 gnd.n7107 gnd.n243 585
R2755 gnd.n4314 gnd.n243 585
R2756 gnd.n240 gnd.n238 585
R2757 gnd.n4298 gnd.n238 585
R2758 gnd.n7112 gnd.n7111 585
R2759 gnd.n7113 gnd.n7112 585
R2760 gnd.n239 gnd.n237 585
R2761 gnd.n4268 gnd.n237 585
R2762 gnd.n4331 gnd.n4330 585
R2763 gnd.n4330 gnd.n4329 585
R2764 gnd.n1495 gnd.n1494 585
R2765 gnd.n4326 gnd.n1495 585
R2766 gnd.n4335 gnd.n1493 585
R2767 gnd.n1532 gnd.n1493 585
R2768 gnd.n4336 gnd.n1492 585
R2769 gnd.n4260 gnd.n1492 585
R2770 gnd.n4337 gnd.n1491 585
R2771 gnd.n4213 gnd.n1491 585
R2772 gnd.n4249 gnd.n1489 585
R2773 gnd.n4250 gnd.n4249 585
R2774 gnd.n4341 gnd.n1488 585
R2775 gnd.n4222 gnd.n1488 585
R2776 gnd.n4342 gnd.n1487 585
R2777 gnd.n4164 gnd.n1487 585
R2778 gnd.n4343 gnd.n1486 585
R2779 gnd.n4207 gnd.n1486 585
R2780 gnd.n1567 gnd.n1484 585
R2781 gnd.n1568 gnd.n1567 585
R2782 gnd.n4347 gnd.n1483 585
R2783 gnd.n4197 gnd.n1483 585
R2784 gnd.n4348 gnd.n1482 585
R2785 gnd.n4185 gnd.n1482 585
R2786 gnd.n4349 gnd.n1481 585
R2787 gnd.n1586 gnd.n1481 585
R2788 gnd.n1478 gnd.n1476 585
R2789 gnd.n4176 gnd.n1476 585
R2790 gnd.n4354 gnd.n4353 585
R2791 gnd.n4355 gnd.n4354 585
R2792 gnd.n1477 gnd.n1475 585
R2793 gnd.n4148 gnd.n1475 585
R2794 gnd.n1645 gnd.n1463 585
R2795 gnd.n4361 gnd.n1463 585
R2796 gnd.n1649 gnd.n1648 585
R2797 gnd.n1651 gnd.n1642 585
R2798 gnd.n1654 gnd.n1653 585
R2799 gnd.n1635 gnd.n1634 585
R2800 gnd.n1668 gnd.n1667 585
R2801 gnd.n1670 gnd.n1633 585
R2802 gnd.n1673 gnd.n1672 585
R2803 gnd.n1626 gnd.n1625 585
R2804 gnd.n1687 gnd.n1686 585
R2805 gnd.n1689 gnd.n1624 585
R2806 gnd.n1692 gnd.n1691 585
R2807 gnd.n1617 gnd.n1616 585
R2808 gnd.n1706 gnd.n1705 585
R2809 gnd.n1708 gnd.n1615 585
R2810 gnd.n1711 gnd.n1710 585
R2811 gnd.n1608 gnd.n1607 585
R2812 gnd.n1725 gnd.n1724 585
R2813 gnd.n1727 gnd.n1606 585
R2814 gnd.n1729 gnd.n1728 585
R2815 gnd.n1728 gnd.n1451 585
R2816 gnd.n7215 gnd.n80 585
R2817 gnd.n7216 gnd.n7214 585
R2818 gnd.n7217 gnd.n7210 585
R2819 gnd.n7208 gnd.n7206 585
R2820 gnd.n7221 gnd.n7205 585
R2821 gnd.n7222 gnd.n7203 585
R2822 gnd.n7223 gnd.n7202 585
R2823 gnd.n7200 gnd.n7198 585
R2824 gnd.n7227 gnd.n7197 585
R2825 gnd.n7228 gnd.n7195 585
R2826 gnd.n7229 gnd.n7194 585
R2827 gnd.n7192 gnd.n7190 585
R2828 gnd.n7233 gnd.n7189 585
R2829 gnd.n7234 gnd.n7187 585
R2830 gnd.n7235 gnd.n7186 585
R2831 gnd.n7184 gnd.n7182 585
R2832 gnd.n7239 gnd.n7181 585
R2833 gnd.n7240 gnd.n7179 585
R2834 gnd.n7241 gnd.n7178 585
R2835 gnd.n7178 gnd.n94 585
R2836 gnd.n7328 gnd.n7327 585
R2837 gnd.n7327 gnd.n7326 585
R2838 gnd.n79 gnd.n77 585
R2839 gnd.n7247 gnd.n79 585
R2840 gnd.n7332 gnd.n76 585
R2841 gnd.n173 gnd.n76 585
R2842 gnd.n7333 gnd.n75 585
R2843 gnd.n7172 gnd.n75 585
R2844 gnd.n7334 gnd.n74 585
R2845 gnd.n7059 gnd.n74 585
R2846 gnd.n181 gnd.n72 585
R2847 gnd.n7162 gnd.n181 585
R2848 gnd.n7338 gnd.n71 585
R2849 gnd.n7065 gnd.n71 585
R2850 gnd.n7339 gnd.n70 585
R2851 gnd.n7154 gnd.n70 585
R2852 gnd.n7340 gnd.n69 585
R2853 gnd.n7048 gnd.n69 585
R2854 gnd.n196 gnd.n67 585
R2855 gnd.n7146 gnd.n196 585
R2856 gnd.n7344 gnd.n66 585
R2857 gnd.n7074 gnd.n66 585
R2858 gnd.n7345 gnd.n65 585
R2859 gnd.n7138 gnd.n65 585
R2860 gnd.n7346 gnd.n64 585
R2861 gnd.n7078 gnd.n64 585
R2862 gnd.n213 gnd.n62 585
R2863 gnd.n7130 gnd.n213 585
R2864 gnd.n7350 gnd.n61 585
R2865 gnd.n7084 gnd.n61 585
R2866 gnd.n7351 gnd.n60 585
R2867 gnd.n7122 gnd.n60 585
R2868 gnd.n7352 gnd.n59 585
R2869 gnd.n4282 gnd.n59 585
R2870 gnd.n250 gnd.n57 585
R2871 gnd.n7098 gnd.n250 585
R2872 gnd.n7356 gnd.n56 585
R2873 gnd.n7094 gnd.n56 585
R2874 gnd.n7357 gnd.n55 585
R2875 gnd.n4290 gnd.n55 585
R2876 gnd.n7358 gnd.n54 585
R2877 gnd.n1518 gnd.n54 585
R2878 gnd.n1511 gnd.n52 585
R2879 gnd.n4309 gnd.n1511 585
R2880 gnd.n4316 gnd.n4315 585
R2881 gnd.n4315 gnd.n4314 585
R2882 gnd.n4318 gnd.n1510 585
R2883 gnd.n4298 gnd.n1510 585
R2884 gnd.n4319 gnd.n235 585
R2885 gnd.n7113 gnd.n235 585
R2886 gnd.n4320 gnd.n1509 585
R2887 gnd.n4268 gnd.n1509 585
R2888 gnd.n1506 gnd.n1498 585
R2889 gnd.n4329 gnd.n1498 585
R2890 gnd.n4325 gnd.n4324 585
R2891 gnd.n4326 gnd.n4325 585
R2892 gnd.n1505 gnd.n1504 585
R2893 gnd.n1532 gnd.n1504 585
R2894 gnd.n4215 gnd.n1531 585
R2895 gnd.n4260 gnd.n1531 585
R2896 gnd.n4216 gnd.n4214 585
R2897 gnd.n4214 gnd.n4213 585
R2898 gnd.n1551 gnd.n1541 585
R2899 gnd.n4250 gnd.n1541 585
R2900 gnd.n4221 gnd.n4220 585
R2901 gnd.n4222 gnd.n4221 585
R2902 gnd.n1550 gnd.n1549 585
R2903 gnd.n4164 gnd.n1549 585
R2904 gnd.n4209 gnd.n4208 585
R2905 gnd.n4208 gnd.n4207 585
R2906 gnd.n1554 gnd.n1553 585
R2907 gnd.n1568 gnd.n1554 585
R2908 gnd.n1590 gnd.n1566 585
R2909 gnd.n4197 gnd.n1566 585
R2910 gnd.n4184 gnd.n4183 585
R2911 gnd.n4185 gnd.n4184 585
R2912 gnd.n1589 gnd.n1588 585
R2913 gnd.n1588 gnd.n1586 585
R2914 gnd.n4178 gnd.n4177 585
R2915 gnd.n4177 gnd.n4176 585
R2916 gnd.n1592 gnd.n1473 585
R2917 gnd.n4355 gnd.n1473 585
R2918 gnd.n4147 gnd.n4146 585
R2919 gnd.n4148 gnd.n4147 585
R2920 gnd.n1597 gnd.n1461 585
R2921 gnd.n4361 gnd.n1461 585
R2922 gnd.n6058 gnd.n6057 585
R2923 gnd.n6057 gnd.n6056 585
R2924 gnd.n6059 gnd.n1008 585
R2925 gnd.n5966 gnd.n1008 585
R2926 gnd.n6061 gnd.n6060 585
R2927 gnd.n6062 gnd.n6061 585
R2928 gnd.n1009 gnd.n1007 585
R2929 gnd.n1007 gnd.n1003 585
R2930 gnd.n988 gnd.n987 585
R2931 gnd.n992 gnd.n988 585
R2932 gnd.n6072 gnd.n6071 585
R2933 gnd.n6071 gnd.n6070 585
R2934 gnd.n6073 gnd.n982 585
R2935 gnd.n5955 gnd.n982 585
R2936 gnd.n6075 gnd.n6074 585
R2937 gnd.n6076 gnd.n6075 585
R2938 gnd.n983 gnd.n981 585
R2939 gnd.n981 gnd.n977 585
R2940 gnd.n963 gnd.n962 585
R2941 gnd.n5948 gnd.n963 585
R2942 gnd.n6086 gnd.n6085 585
R2943 gnd.n6085 gnd.n6084 585
R2944 gnd.n6087 gnd.n957 585
R2945 gnd.n5615 gnd.n957 585
R2946 gnd.n6089 gnd.n6088 585
R2947 gnd.n6090 gnd.n6089 585
R2948 gnd.n958 gnd.n956 585
R2949 gnd.n956 gnd.n952 585
R2950 gnd.n940 gnd.n939 585
R2951 gnd.n5623 gnd.n940 585
R2952 gnd.n6100 gnd.n6099 585
R2953 gnd.n6099 gnd.n6098 585
R2954 gnd.n6101 gnd.n934 585
R2955 gnd.n4835 gnd.n934 585
R2956 gnd.n6103 gnd.n6102 585
R2957 gnd.n6104 gnd.n6103 585
R2958 gnd.n935 gnd.n933 585
R2959 gnd.n5632 gnd.n933 585
R2960 gnd.n5597 gnd.n4851 585
R2961 gnd.n4851 gnd.n4841 585
R2962 gnd.n5599 gnd.n5598 585
R2963 gnd.n5600 gnd.n5599 585
R2964 gnd.n4852 gnd.n4850 585
R2965 gnd.n4860 gnd.n4850 585
R2966 gnd.n5573 gnd.n4872 585
R2967 gnd.n4872 gnd.n4859 585
R2968 gnd.n5575 gnd.n5574 585
R2969 gnd.n5576 gnd.n5575 585
R2970 gnd.n4873 gnd.n4871 585
R2971 gnd.n4871 gnd.n4867 585
R2972 gnd.n5561 gnd.n5560 585
R2973 gnd.n5560 gnd.n5559 585
R2974 gnd.n4878 gnd.n4877 585
R2975 gnd.n4887 gnd.n4878 585
R2976 gnd.n5550 gnd.n5549 585
R2977 gnd.n5549 gnd.n5548 585
R2978 gnd.n4885 gnd.n4884 585
R2979 gnd.n5536 gnd.n4885 585
R2980 gnd.n4974 gnd.n4973 585
R2981 gnd.n4974 gnd.n4894 585
R2982 gnd.n5493 gnd.n5492 585
R2983 gnd.n5492 gnd.n5491 585
R2984 gnd.n5494 gnd.n4968 585
R2985 gnd.n4979 gnd.n4968 585
R2986 gnd.n5496 gnd.n5495 585
R2987 gnd.n5497 gnd.n5496 585
R2988 gnd.n4969 gnd.n4967 585
R2989 gnd.n4992 gnd.n4967 585
R2990 gnd.n4952 gnd.n4951 585
R2991 gnd.n4955 gnd.n4952 585
R2992 gnd.n5507 gnd.n5506 585
R2993 gnd.n5506 gnd.n5505 585
R2994 gnd.n5508 gnd.n4946 585
R2995 gnd.n5467 gnd.n4946 585
R2996 gnd.n5510 gnd.n5509 585
R2997 gnd.n5511 gnd.n5510 585
R2998 gnd.n4947 gnd.n4945 585
R2999 gnd.n5006 gnd.n4945 585
R3000 gnd.n5459 gnd.n5458 585
R3001 gnd.n5458 gnd.n5457 585
R3002 gnd.n5003 gnd.n5002 585
R3003 gnd.n5441 gnd.n5003 585
R3004 gnd.n5428 gnd.n5022 585
R3005 gnd.n5022 gnd.n5021 585
R3006 gnd.n5430 gnd.n5429 585
R3007 gnd.n5431 gnd.n5430 585
R3008 gnd.n5023 gnd.n5020 585
R3009 gnd.n5029 gnd.n5020 585
R3010 gnd.n5409 gnd.n5408 585
R3011 gnd.n5410 gnd.n5409 585
R3012 gnd.n5040 gnd.n5039 585
R3013 gnd.n5039 gnd.n5035 585
R3014 gnd.n5399 gnd.n5398 585
R3015 gnd.n5400 gnd.n5399 585
R3016 gnd.n5050 gnd.n5049 585
R3017 gnd.n5055 gnd.n5049 585
R3018 gnd.n5377 gnd.n5068 585
R3019 gnd.n5068 gnd.n5054 585
R3020 gnd.n5379 gnd.n5378 585
R3021 gnd.n5380 gnd.n5379 585
R3022 gnd.n5069 gnd.n5067 585
R3023 gnd.n5067 gnd.n5063 585
R3024 gnd.n5368 gnd.n5367 585
R3025 gnd.n5369 gnd.n5368 585
R3026 gnd.n5076 gnd.n5075 585
R3027 gnd.n5080 gnd.n5075 585
R3028 gnd.n5345 gnd.n5097 585
R3029 gnd.n5097 gnd.n5079 585
R3030 gnd.n5347 gnd.n5346 585
R3031 gnd.n5348 gnd.n5347 585
R3032 gnd.n5098 gnd.n5096 585
R3033 gnd.n5096 gnd.n5087 585
R3034 gnd.n5340 gnd.n5339 585
R3035 gnd.n5339 gnd.n5338 585
R3036 gnd.n5145 gnd.n5144 585
R3037 gnd.n5146 gnd.n5145 585
R3038 gnd.n5299 gnd.n5298 585
R3039 gnd.n5300 gnd.n5299 585
R3040 gnd.n5155 gnd.n5154 585
R3041 gnd.n5154 gnd.n5153 585
R3042 gnd.n5294 gnd.n5293 585
R3043 gnd.n5293 gnd.n5292 585
R3044 gnd.n5158 gnd.n5157 585
R3045 gnd.n5159 gnd.n5158 585
R3046 gnd.n5283 gnd.n5282 585
R3047 gnd.n5284 gnd.n5283 585
R3048 gnd.n5166 gnd.n5165 585
R3049 gnd.n5275 gnd.n5165 585
R3050 gnd.n5278 gnd.n5277 585
R3051 gnd.n5277 gnd.n5276 585
R3052 gnd.n5169 gnd.n5168 585
R3053 gnd.n5170 gnd.n5169 585
R3054 gnd.n5264 gnd.n5263 585
R3055 gnd.n5262 gnd.n5188 585
R3056 gnd.n5261 gnd.n5187 585
R3057 gnd.n5266 gnd.n5187 585
R3058 gnd.n5260 gnd.n5259 585
R3059 gnd.n5258 gnd.n5257 585
R3060 gnd.n5256 gnd.n5255 585
R3061 gnd.n5254 gnd.n5253 585
R3062 gnd.n5252 gnd.n5251 585
R3063 gnd.n5250 gnd.n5249 585
R3064 gnd.n5248 gnd.n5247 585
R3065 gnd.n5246 gnd.n5245 585
R3066 gnd.n5244 gnd.n5243 585
R3067 gnd.n5242 gnd.n5241 585
R3068 gnd.n5240 gnd.n5239 585
R3069 gnd.n5238 gnd.n5237 585
R3070 gnd.n5236 gnd.n5235 585
R3071 gnd.n5234 gnd.n5233 585
R3072 gnd.n5232 gnd.n5231 585
R3073 gnd.n5230 gnd.n5229 585
R3074 gnd.n5228 gnd.n5227 585
R3075 gnd.n5226 gnd.n5225 585
R3076 gnd.n5224 gnd.n5223 585
R3077 gnd.n5222 gnd.n5221 585
R3078 gnd.n5220 gnd.n5219 585
R3079 gnd.n5218 gnd.n5217 585
R3080 gnd.n5175 gnd.n5174 585
R3081 gnd.n5269 gnd.n5268 585
R3082 gnd.n5974 gnd.n5973 585
R3083 gnd.n5975 gnd.n4820 585
R3084 gnd.n5977 gnd.n5976 585
R3085 gnd.n5979 gnd.n4819 585
R3086 gnd.n5981 gnd.n5980 585
R3087 gnd.n5982 gnd.n4810 585
R3088 gnd.n5984 gnd.n5983 585
R3089 gnd.n5986 gnd.n4808 585
R3090 gnd.n5988 gnd.n5987 585
R3091 gnd.n5989 gnd.n4803 585
R3092 gnd.n5991 gnd.n5990 585
R3093 gnd.n5993 gnd.n4801 585
R3094 gnd.n5995 gnd.n5994 585
R3095 gnd.n5996 gnd.n4796 585
R3096 gnd.n5998 gnd.n5997 585
R3097 gnd.n6000 gnd.n4794 585
R3098 gnd.n6002 gnd.n6001 585
R3099 gnd.n6003 gnd.n4789 585
R3100 gnd.n6005 gnd.n6004 585
R3101 gnd.n6007 gnd.n4787 585
R3102 gnd.n6009 gnd.n6008 585
R3103 gnd.n6010 gnd.n4782 585
R3104 gnd.n6012 gnd.n6011 585
R3105 gnd.n6014 gnd.n4780 585
R3106 gnd.n6016 gnd.n6015 585
R3107 gnd.n6017 gnd.n4778 585
R3108 gnd.n6018 gnd.n1013 585
R3109 gnd.n4741 gnd.n1013 585
R3110 gnd.n5969 gnd.n1015 585
R3111 gnd.n6056 gnd.n1015 585
R3112 gnd.n5968 gnd.n5967 585
R3113 gnd.n5967 gnd.n5966 585
R3114 gnd.n5965 gnd.n1005 585
R3115 gnd.n6062 gnd.n1005 585
R3116 gnd.n5959 gnd.n4825 585
R3117 gnd.n5959 gnd.n1003 585
R3118 gnd.n5961 gnd.n5960 585
R3119 gnd.n5960 gnd.n992 585
R3120 gnd.n5958 gnd.n990 585
R3121 gnd.n6070 gnd.n990 585
R3122 gnd.n5957 gnd.n5956 585
R3123 gnd.n5956 gnd.n5955 585
R3124 gnd.n4827 gnd.n979 585
R3125 gnd.n6076 gnd.n979 585
R3126 gnd.n5951 gnd.n5950 585
R3127 gnd.n5950 gnd.n977 585
R3128 gnd.n5949 gnd.n4829 585
R3129 gnd.n5949 gnd.n5948 585
R3130 gnd.n5614 gnd.n965 585
R3131 gnd.n6084 gnd.n965 585
R3132 gnd.n5617 gnd.n5616 585
R3133 gnd.n5616 gnd.n5615 585
R3134 gnd.n5618 gnd.n954 585
R3135 gnd.n6090 gnd.n954 585
R3136 gnd.n5620 gnd.n5619 585
R3137 gnd.n5620 gnd.n952 585
R3138 gnd.n5625 gnd.n5624 585
R3139 gnd.n5624 gnd.n5623 585
R3140 gnd.n5626 gnd.n942 585
R3141 gnd.n6098 gnd.n942 585
R3142 gnd.n5628 gnd.n5627 585
R3143 gnd.n5627 gnd.n4835 585
R3144 gnd.n5629 gnd.n932 585
R3145 gnd.n6104 gnd.n932 585
R3146 gnd.n5631 gnd.n5630 585
R3147 gnd.n5632 gnd.n5631 585
R3148 gnd.n4844 gnd.n4843 585
R3149 gnd.n4843 gnd.n4841 585
R3150 gnd.n5602 gnd.n5601 585
R3151 gnd.n5601 gnd.n5600 585
R3152 gnd.n4847 gnd.n4846 585
R3153 gnd.n4860 gnd.n4847 585
R3154 gnd.n5524 gnd.n5523 585
R3155 gnd.n5523 gnd.n4859 585
R3156 gnd.n5525 gnd.n4869 585
R3157 gnd.n5576 gnd.n4869 585
R3158 gnd.n5527 gnd.n5526 585
R3159 gnd.n5526 gnd.n4867 585
R3160 gnd.n5528 gnd.n4880 585
R3161 gnd.n5559 gnd.n4880 585
R3162 gnd.n5530 gnd.n5529 585
R3163 gnd.n5529 gnd.n4887 585
R3164 gnd.n5531 gnd.n4886 585
R3165 gnd.n5548 gnd.n4886 585
R3166 gnd.n5533 gnd.n5532 585
R3167 gnd.n5536 gnd.n5533 585
R3168 gnd.n4897 gnd.n4896 585
R3169 gnd.n4896 gnd.n4894 585
R3170 gnd.n4976 gnd.n4975 585
R3171 gnd.n5491 gnd.n4975 585
R3172 gnd.n4978 gnd.n4977 585
R3173 gnd.n4979 gnd.n4978 585
R3174 gnd.n4989 gnd.n4965 585
R3175 gnd.n5497 gnd.n4965 585
R3176 gnd.n4991 gnd.n4990 585
R3177 gnd.n4992 gnd.n4991 585
R3178 gnd.n4988 gnd.n4987 585
R3179 gnd.n4988 gnd.n4955 585
R3180 gnd.n4986 gnd.n4953 585
R3181 gnd.n5505 gnd.n4953 585
R3182 gnd.n4942 gnd.n4940 585
R3183 gnd.n5467 gnd.n4942 585
R3184 gnd.n5513 gnd.n5512 585
R3185 gnd.n5512 gnd.n5511 585
R3186 gnd.n4941 gnd.n4939 585
R3187 gnd.n5006 gnd.n4941 585
R3188 gnd.n5438 gnd.n5005 585
R3189 gnd.n5457 gnd.n5005 585
R3190 gnd.n5440 gnd.n5439 585
R3191 gnd.n5441 gnd.n5440 585
R3192 gnd.n5015 gnd.n5014 585
R3193 gnd.n5021 gnd.n5014 585
R3194 gnd.n5433 gnd.n5432 585
R3195 gnd.n5432 gnd.n5431 585
R3196 gnd.n5018 gnd.n5017 585
R3197 gnd.n5029 gnd.n5018 585
R3198 gnd.n5318 gnd.n5037 585
R3199 gnd.n5410 gnd.n5037 585
R3200 gnd.n5320 gnd.n5319 585
R3201 gnd.n5319 gnd.n5035 585
R3202 gnd.n5321 gnd.n5048 585
R3203 gnd.n5400 gnd.n5048 585
R3204 gnd.n5323 gnd.n5322 585
R3205 gnd.n5323 gnd.n5055 585
R3206 gnd.n5325 gnd.n5324 585
R3207 gnd.n5324 gnd.n5054 585
R3208 gnd.n5326 gnd.n5065 585
R3209 gnd.n5380 gnd.n5065 585
R3210 gnd.n5328 gnd.n5327 585
R3211 gnd.n5327 gnd.n5063 585
R3212 gnd.n5329 gnd.n5074 585
R3213 gnd.n5369 gnd.n5074 585
R3214 gnd.n5331 gnd.n5330 585
R3215 gnd.n5331 gnd.n5080 585
R3216 gnd.n5333 gnd.n5332 585
R3217 gnd.n5332 gnd.n5079 585
R3218 gnd.n5334 gnd.n5095 585
R3219 gnd.n5348 gnd.n5095 585
R3220 gnd.n5335 gnd.n5148 585
R3221 gnd.n5148 gnd.n5087 585
R3222 gnd.n5337 gnd.n5336 585
R3223 gnd.n5338 gnd.n5337 585
R3224 gnd.n5149 gnd.n5147 585
R3225 gnd.n5147 gnd.n5146 585
R3226 gnd.n5302 gnd.n5301 585
R3227 gnd.n5301 gnd.n5300 585
R3228 gnd.n5152 gnd.n5151 585
R3229 gnd.n5153 gnd.n5152 585
R3230 gnd.n5291 gnd.n5290 585
R3231 gnd.n5292 gnd.n5291 585
R3232 gnd.n5161 gnd.n5160 585
R3233 gnd.n5160 gnd.n5159 585
R3234 gnd.n5286 gnd.n5285 585
R3235 gnd.n5285 gnd.n5284 585
R3236 gnd.n5164 gnd.n5163 585
R3237 gnd.n5275 gnd.n5164 585
R3238 gnd.n5274 gnd.n5273 585
R3239 gnd.n5276 gnd.n5274 585
R3240 gnd.n5172 gnd.n5171 585
R3241 gnd.n5171 gnd.n5170 585
R3242 gnd.n6054 gnd.n6053 585
R3243 gnd.n6055 gnd.n6054 585
R3244 gnd.n4744 gnd.n4742 585
R3245 gnd.n4742 gnd.n1014 585
R3246 gnd.n1002 gnd.n1001 585
R3247 gnd.n1006 gnd.n1002 585
R3248 gnd.n6065 gnd.n6064 585
R3249 gnd.n6064 gnd.n6063 585
R3250 gnd.n6066 gnd.n994 585
R3251 gnd.n5936 gnd.n994 585
R3252 gnd.n6068 gnd.n6067 585
R3253 gnd.n6069 gnd.n6068 585
R3254 gnd.n995 gnd.n993 585
R3255 gnd.n993 gnd.n989 585
R3256 gnd.n976 gnd.n975 585
R3257 gnd.n980 gnd.n976 585
R3258 gnd.n6079 gnd.n6078 585
R3259 gnd.n6078 gnd.n6077 585
R3260 gnd.n6080 gnd.n968 585
R3261 gnd.n5947 gnd.n968 585
R3262 gnd.n6082 gnd.n6081 585
R3263 gnd.n6083 gnd.n6082 585
R3264 gnd.n969 gnd.n967 585
R3265 gnd.n967 gnd.n964 585
R3266 gnd.n951 gnd.n950 585
R3267 gnd.n955 gnd.n951 585
R3268 gnd.n6093 gnd.n6092 585
R3269 gnd.n6092 gnd.n6091 585
R3270 gnd.n6094 gnd.n945 585
R3271 gnd.n5622 gnd.n945 585
R3272 gnd.n6096 gnd.n6095 585
R3273 gnd.n6097 gnd.n6096 585
R3274 gnd.n946 gnd.n944 585
R3275 gnd.n944 gnd.n941 585
R3276 gnd.n5641 gnd.n5640 585
R3277 gnd.n5642 gnd.n5641 585
R3278 gnd.n4837 gnd.n4836 585
R3279 gnd.n4836 gnd.n931 585
R3280 gnd.n5635 gnd.n5634 585
R3281 gnd.n5634 gnd.n5633 585
R3282 gnd.n4840 gnd.n4839 585
R3283 gnd.n4849 gnd.n4840 585
R3284 gnd.n5584 gnd.n4862 585
R3285 gnd.n4862 gnd.n4848 585
R3286 gnd.n5586 gnd.n5585 585
R3287 gnd.n5587 gnd.n5586 585
R3288 gnd.n4863 gnd.n4861 585
R3289 gnd.n4870 gnd.n4861 585
R3290 gnd.n5579 gnd.n5578 585
R3291 gnd.n5578 gnd.n5577 585
R3292 gnd.n4866 gnd.n4865 585
R3293 gnd.n5558 gnd.n4866 585
R3294 gnd.n5544 gnd.n4889 585
R3295 gnd.n4889 gnd.n4879 585
R3296 gnd.n5546 gnd.n5545 585
R3297 gnd.n5547 gnd.n5546 585
R3298 gnd.n4890 gnd.n4888 585
R3299 gnd.n5535 gnd.n4888 585
R3300 gnd.n5539 gnd.n5538 585
R3301 gnd.n5538 gnd.n5537 585
R3302 gnd.n4893 gnd.n4892 585
R3303 gnd.n5490 gnd.n4893 585
R3304 gnd.n4983 gnd.n4982 585
R3305 gnd.n4984 gnd.n4983 585
R3306 gnd.n4963 gnd.n4962 585
R3307 gnd.n4966 gnd.n4963 585
R3308 gnd.n5500 gnd.n5499 585
R3309 gnd.n5499 gnd.n5498 585
R3310 gnd.n5501 gnd.n4957 585
R3311 gnd.n4993 gnd.n4957 585
R3312 gnd.n5503 gnd.n5502 585
R3313 gnd.n5504 gnd.n5503 585
R3314 gnd.n4958 gnd.n4956 585
R3315 gnd.n5468 gnd.n4956 585
R3316 gnd.n5452 gnd.n5451 585
R3317 gnd.n5451 gnd.n4944 585
R3318 gnd.n5453 gnd.n5008 585
R3319 gnd.n5008 gnd.n4943 585
R3320 gnd.n5455 gnd.n5454 585
R3321 gnd.n5456 gnd.n5455 585
R3322 gnd.n5009 gnd.n5007 585
R3323 gnd.n5007 gnd.n5004 585
R3324 gnd.n5444 gnd.n5443 585
R3325 gnd.n5443 gnd.n5442 585
R3326 gnd.n5012 gnd.n5011 585
R3327 gnd.n5019 gnd.n5012 585
R3328 gnd.n5418 gnd.n5417 585
R3329 gnd.n5419 gnd.n5418 585
R3330 gnd.n5031 gnd.n5030 585
R3331 gnd.n5038 gnd.n5030 585
R3332 gnd.n5413 gnd.n5412 585
R3333 gnd.n5412 gnd.n5411 585
R3334 gnd.n5034 gnd.n5033 585
R3335 gnd.n5401 gnd.n5034 585
R3336 gnd.n5388 gnd.n5058 585
R3337 gnd.n5058 gnd.n5057 585
R3338 gnd.n5390 gnd.n5389 585
R3339 gnd.n5391 gnd.n5390 585
R3340 gnd.n5059 gnd.n5056 585
R3341 gnd.n5066 gnd.n5056 585
R3342 gnd.n5383 gnd.n5382 585
R3343 gnd.n5382 gnd.n5381 585
R3344 gnd.n5062 gnd.n5061 585
R3345 gnd.n5370 gnd.n5062 585
R3346 gnd.n5357 gnd.n5083 585
R3347 gnd.n5083 gnd.n5082 585
R3348 gnd.n5359 gnd.n5358 585
R3349 gnd.n5360 gnd.n5359 585
R3350 gnd.n5353 gnd.n5081 585
R3351 gnd.n5352 gnd.n5351 585
R3352 gnd.n5086 gnd.n5085 585
R3353 gnd.n5349 gnd.n5086 585
R3354 gnd.n5108 gnd.n5107 585
R3355 gnd.n5111 gnd.n5110 585
R3356 gnd.n5109 gnd.n5104 585
R3357 gnd.n5116 gnd.n5115 585
R3358 gnd.n5118 gnd.n5117 585
R3359 gnd.n5121 gnd.n5120 585
R3360 gnd.n5119 gnd.n5102 585
R3361 gnd.n5126 gnd.n5125 585
R3362 gnd.n5128 gnd.n5127 585
R3363 gnd.n5131 gnd.n5130 585
R3364 gnd.n5129 gnd.n5100 585
R3365 gnd.n5136 gnd.n5135 585
R3366 gnd.n5140 gnd.n5137 585
R3367 gnd.n5141 gnd.n5078 585
R3368 gnd.n6023 gnd.n6022 585
R3369 gnd.n6025 gnd.n4773 585
R3370 gnd.n6027 gnd.n6026 585
R3371 gnd.n6028 gnd.n4766 585
R3372 gnd.n6030 gnd.n6029 585
R3373 gnd.n6032 gnd.n4764 585
R3374 gnd.n6034 gnd.n6033 585
R3375 gnd.n6035 gnd.n4759 585
R3376 gnd.n6037 gnd.n6036 585
R3377 gnd.n6039 gnd.n4757 585
R3378 gnd.n6041 gnd.n6040 585
R3379 gnd.n6042 gnd.n4752 585
R3380 gnd.n6044 gnd.n6043 585
R3381 gnd.n6046 gnd.n4750 585
R3382 gnd.n6048 gnd.n6047 585
R3383 gnd.n6049 gnd.n4748 585
R3384 gnd.n6050 gnd.n4743 585
R3385 gnd.n4743 gnd.n4741 585
R3386 gnd.n5930 gnd.n1016 585
R3387 gnd.n6055 gnd.n1016 585
R3388 gnd.n5932 gnd.n5931 585
R3389 gnd.n5932 gnd.n1014 585
R3390 gnd.n5934 gnd.n5933 585
R3391 gnd.n5933 gnd.n1006 585
R3392 gnd.n5935 gnd.n1004 585
R3393 gnd.n6063 gnd.n1004 585
R3394 gnd.n5938 gnd.n5937 585
R3395 gnd.n5937 gnd.n5936 585
R3396 gnd.n5939 gnd.n991 585
R3397 gnd.n6069 gnd.n991 585
R3398 gnd.n5941 gnd.n5940 585
R3399 gnd.n5941 gnd.n989 585
R3400 gnd.n5943 gnd.n5942 585
R3401 gnd.n5942 gnd.n980 585
R3402 gnd.n5944 gnd.n978 585
R3403 gnd.n6077 gnd.n978 585
R3404 gnd.n5946 gnd.n5945 585
R3405 gnd.n5947 gnd.n5946 585
R3406 gnd.n5659 gnd.n966 585
R3407 gnd.n6083 gnd.n966 585
R3408 gnd.n5658 gnd.n5657 585
R3409 gnd.n5657 gnd.n964 585
R3410 gnd.n5656 gnd.n5654 585
R3411 gnd.n5656 gnd.n955 585
R3412 gnd.n5652 gnd.n953 585
R3413 gnd.n6091 gnd.n953 585
R3414 gnd.n5621 gnd.n4830 585
R3415 gnd.n5622 gnd.n5621 585
R3416 gnd.n5646 gnd.n943 585
R3417 gnd.n6097 gnd.n943 585
R3418 gnd.n5645 gnd.n5644 585
R3419 gnd.n5644 gnd.n941 585
R3420 gnd.n5643 gnd.n4832 585
R3421 gnd.n5643 gnd.n5642 585
R3422 gnd.n5593 gnd.n4834 585
R3423 gnd.n4834 gnd.n931 585
R3424 gnd.n5594 gnd.n4842 585
R3425 gnd.n5633 gnd.n4842 585
R3426 gnd.n5591 gnd.n5590 585
R3427 gnd.n5590 gnd.n4849 585
R3428 gnd.n5589 gnd.n4856 585
R3429 gnd.n5589 gnd.n4848 585
R3430 gnd.n5588 gnd.n4858 585
R3431 gnd.n5588 gnd.n5587 585
R3432 gnd.n5567 gnd.n4857 585
R3433 gnd.n4870 gnd.n4857 585
R3434 gnd.n5566 gnd.n4868 585
R3435 gnd.n5577 gnd.n4868 585
R3436 gnd.n5557 gnd.n4875 585
R3437 gnd.n5558 gnd.n5557 585
R3438 gnd.n5556 gnd.n5555 585
R3439 gnd.n5556 gnd.n4879 585
R3440 gnd.n5554 gnd.n4881 585
R3441 gnd.n5547 gnd.n4881 585
R3442 gnd.n5534 gnd.n4882 585
R3443 gnd.n5535 gnd.n5534 585
R3444 gnd.n5487 gnd.n4895 585
R3445 gnd.n5537 gnd.n4895 585
R3446 gnd.n5489 gnd.n5488 585
R3447 gnd.n5490 gnd.n5489 585
R3448 gnd.n5482 gnd.n4985 585
R3449 gnd.n4985 gnd.n4984 585
R3450 gnd.n5480 gnd.n5479 585
R3451 gnd.n5479 gnd.n4966 585
R3452 gnd.n5477 gnd.n4964 585
R3453 gnd.n5498 gnd.n4964 585
R3454 gnd.n4995 gnd.n4994 585
R3455 gnd.n4994 gnd.n4993 585
R3456 gnd.n5471 gnd.n4954 585
R3457 gnd.n5504 gnd.n4954 585
R3458 gnd.n5470 gnd.n5469 585
R3459 gnd.n5469 gnd.n5468 585
R3460 gnd.n5466 gnd.n4997 585
R3461 gnd.n5466 gnd.n4944 585
R3462 gnd.n5465 gnd.n5464 585
R3463 gnd.n5465 gnd.n4943 585
R3464 gnd.n5000 gnd.n4999 585
R3465 gnd.n5456 gnd.n4999 585
R3466 gnd.n5424 gnd.n5423 585
R3467 gnd.n5423 gnd.n5004 585
R3468 gnd.n5425 gnd.n5013 585
R3469 gnd.n5442 gnd.n5013 585
R3470 gnd.n5422 gnd.n5421 585
R3471 gnd.n5421 gnd.n5019 585
R3472 gnd.n5420 gnd.n5027 585
R3473 gnd.n5420 gnd.n5419 585
R3474 gnd.n5405 gnd.n5028 585
R3475 gnd.n5038 gnd.n5028 585
R3476 gnd.n5404 gnd.n5036 585
R3477 gnd.n5411 gnd.n5036 585
R3478 gnd.n5403 gnd.n5402 585
R3479 gnd.n5402 gnd.n5401 585
R3480 gnd.n5047 gnd.n5044 585
R3481 gnd.n5057 gnd.n5047 585
R3482 gnd.n5393 gnd.n5392 585
R3483 gnd.n5392 gnd.n5391 585
R3484 gnd.n5053 gnd.n5052 585
R3485 gnd.n5066 gnd.n5053 585
R3486 gnd.n5373 gnd.n5064 585
R3487 gnd.n5381 gnd.n5064 585
R3488 gnd.n5372 gnd.n5371 585
R3489 gnd.n5371 gnd.n5370 585
R3490 gnd.n5073 gnd.n5071 585
R3491 gnd.n5082 gnd.n5073 585
R3492 gnd.n5362 gnd.n5361 585
R3493 gnd.n5361 gnd.n5360 585
R3494 gnd.n4510 gnd.n4509 585
R3495 gnd.n4509 gnd.n4508 585
R3496 gnd.n4511 gnd.n1320 585
R3497 gnd.n3239 gnd.n1320 585
R3498 gnd.n4513 gnd.n4512 585
R3499 gnd.n4514 gnd.n4513 585
R3500 gnd.n1304 gnd.n1303 585
R3501 gnd.n2943 gnd.n1304 585
R3502 gnd.n4522 gnd.n4521 585
R3503 gnd.n4521 gnd.n4520 585
R3504 gnd.n4523 gnd.n1298 585
R3505 gnd.n2934 gnd.n1298 585
R3506 gnd.n4525 gnd.n4524 585
R3507 gnd.n4526 gnd.n4525 585
R3508 gnd.n1283 gnd.n1282 585
R3509 gnd.n2930 gnd.n1283 585
R3510 gnd.n4534 gnd.n4533 585
R3511 gnd.n4533 gnd.n4532 585
R3512 gnd.n4535 gnd.n1277 585
R3513 gnd.n2923 gnd.n1277 585
R3514 gnd.n4537 gnd.n4536 585
R3515 gnd.n4538 gnd.n4537 585
R3516 gnd.n1262 gnd.n1261 585
R3517 gnd.n2960 gnd.n1262 585
R3518 gnd.n4546 gnd.n4545 585
R3519 gnd.n4545 gnd.n4544 585
R3520 gnd.n4547 gnd.n1256 585
R3521 gnd.n2915 gnd.n1256 585
R3522 gnd.n4549 gnd.n4548 585
R3523 gnd.n4550 gnd.n4549 585
R3524 gnd.n1241 gnd.n1240 585
R3525 gnd.n2907 gnd.n1241 585
R3526 gnd.n4558 gnd.n4557 585
R3527 gnd.n4557 gnd.n4556 585
R3528 gnd.n4559 gnd.n1238 585
R3529 gnd.n2868 gnd.n1238 585
R3530 gnd.n4562 gnd.n4561 585
R3531 gnd.n4563 gnd.n4562 585
R3532 gnd.n1239 gnd.n1224 585
R3533 gnd.n2876 gnd.n1224 585
R3534 gnd.n4571 gnd.n4570 585
R3535 gnd.n4570 gnd.n4569 585
R3536 gnd.n4572 gnd.n1221 585
R3537 gnd.n2854 gnd.n1221 585
R3538 gnd.n4575 gnd.n4574 585
R3539 gnd.n4576 gnd.n4575 585
R3540 gnd.n1222 gnd.n1203 585
R3541 gnd.n2887 gnd.n1203 585
R3542 gnd.n4584 gnd.n4583 585
R3543 gnd.n4583 gnd.n4582 585
R3544 gnd.n4585 gnd.n1201 585
R3545 gnd.n2893 gnd.n1201 585
R3546 gnd.n4587 gnd.n1197 585
R3547 gnd.n2611 gnd.n1197 585
R3548 gnd.n4589 gnd.n4588 585
R3549 gnd.n4590 gnd.n4589 585
R3550 gnd.n1182 gnd.n1181 585
R3551 gnd.n2837 gnd.n1182 585
R3552 gnd.n4598 gnd.n4597 585
R3553 gnd.n4597 gnd.n4596 585
R3554 gnd.n4599 gnd.n1176 585
R3555 gnd.n2825 gnd.n1176 585
R3556 gnd.n4601 gnd.n4600 585
R3557 gnd.n4602 gnd.n4601 585
R3558 gnd.n1161 gnd.n1160 585
R3559 gnd.n2816 gnd.n1161 585
R3560 gnd.n4610 gnd.n4609 585
R3561 gnd.n4609 gnd.n4608 585
R3562 gnd.n4611 gnd.n1155 585
R3563 gnd.n2808 gnd.n1155 585
R3564 gnd.n4613 gnd.n4612 585
R3565 gnd.n4614 gnd.n4613 585
R3566 gnd.n1141 gnd.n1140 585
R3567 gnd.n2800 gnd.n1141 585
R3568 gnd.n4622 gnd.n4621 585
R3569 gnd.n4621 gnd.n4620 585
R3570 gnd.n4623 gnd.n1135 585
R3571 gnd.n2747 gnd.n1135 585
R3572 gnd.n4625 gnd.n4624 585
R3573 gnd.n4626 gnd.n4625 585
R3574 gnd.n1136 gnd.n1134 585
R3575 gnd.n2753 gnd.n1134 585
R3576 gnd.n2666 gnd.n2665 585
R3577 gnd.n2667 gnd.n2666 585
R3578 gnd.n2661 gnd.n1072 585
R3579 gnd.n4635 gnd.n1072 585
R3580 gnd.n4713 gnd.n4712 585
R3581 gnd.n4711 gnd.n1071 585
R3582 gnd.n4710 gnd.n1070 585
R3583 gnd.n4715 gnd.n1070 585
R3584 gnd.n4709 gnd.n4708 585
R3585 gnd.n4707 gnd.n4706 585
R3586 gnd.n4705 gnd.n4704 585
R3587 gnd.n4703 gnd.n4702 585
R3588 gnd.n4701 gnd.n4700 585
R3589 gnd.n4699 gnd.n4698 585
R3590 gnd.n4697 gnd.n4696 585
R3591 gnd.n4695 gnd.n4694 585
R3592 gnd.n4693 gnd.n4692 585
R3593 gnd.n4691 gnd.n4690 585
R3594 gnd.n4689 gnd.n4688 585
R3595 gnd.n4687 gnd.n4686 585
R3596 gnd.n4685 gnd.n4684 585
R3597 gnd.n4683 gnd.n4682 585
R3598 gnd.n4681 gnd.n4680 585
R3599 gnd.n4678 gnd.n4677 585
R3600 gnd.n4676 gnd.n4675 585
R3601 gnd.n4674 gnd.n4673 585
R3602 gnd.n4672 gnd.n4671 585
R3603 gnd.n4670 gnd.n4669 585
R3604 gnd.n4668 gnd.n4667 585
R3605 gnd.n4666 gnd.n4665 585
R3606 gnd.n4664 gnd.n4663 585
R3607 gnd.n4662 gnd.n4661 585
R3608 gnd.n4660 gnd.n4659 585
R3609 gnd.n4658 gnd.n4657 585
R3610 gnd.n4656 gnd.n4655 585
R3611 gnd.n4654 gnd.n4653 585
R3612 gnd.n4652 gnd.n4651 585
R3613 gnd.n4650 gnd.n4649 585
R3614 gnd.n4648 gnd.n4647 585
R3615 gnd.n4646 gnd.n4645 585
R3616 gnd.n4644 gnd.n4643 585
R3617 gnd.n4642 gnd.n1111 585
R3618 gnd.n1115 gnd.n1112 585
R3619 gnd.n4638 gnd.n4637 585
R3620 gnd.n3246 gnd.n3245 585
R3621 gnd.n3248 gnd.n2489 585
R3622 gnd.n3250 gnd.n3249 585
R3623 gnd.n3251 gnd.n2482 585
R3624 gnd.n3253 gnd.n3252 585
R3625 gnd.n3255 gnd.n2480 585
R3626 gnd.n3257 gnd.n3256 585
R3627 gnd.n3258 gnd.n2475 585
R3628 gnd.n3260 gnd.n3259 585
R3629 gnd.n3262 gnd.n2473 585
R3630 gnd.n3264 gnd.n3263 585
R3631 gnd.n3265 gnd.n2468 585
R3632 gnd.n3267 gnd.n3266 585
R3633 gnd.n3269 gnd.n2466 585
R3634 gnd.n3271 gnd.n3270 585
R3635 gnd.n3272 gnd.n2461 585
R3636 gnd.n3274 gnd.n3273 585
R3637 gnd.n3276 gnd.n2460 585
R3638 gnd.n3277 gnd.n2403 585
R3639 gnd.n3280 gnd.n3279 585
R3640 gnd.n2404 gnd.n2396 585
R3641 gnd.n2432 gnd.n2397 585
R3642 gnd.n2434 gnd.n2433 585
R3643 gnd.n2436 gnd.n2435 585
R3644 gnd.n2438 gnd.n2437 585
R3645 gnd.n2440 gnd.n2439 585
R3646 gnd.n2442 gnd.n2441 585
R3647 gnd.n2444 gnd.n2443 585
R3648 gnd.n2446 gnd.n2445 585
R3649 gnd.n2448 gnd.n2447 585
R3650 gnd.n2450 gnd.n2449 585
R3651 gnd.n2452 gnd.n2451 585
R3652 gnd.n2454 gnd.n2453 585
R3653 gnd.n2455 gnd.n2414 585
R3654 gnd.n2457 gnd.n2456 585
R3655 gnd.n2415 gnd.n2413 585
R3656 gnd.n2416 gnd.n1325 585
R3657 gnd.n2459 gnd.n1325 585
R3658 gnd.n3242 gnd.n1327 585
R3659 gnd.n4508 gnd.n1327 585
R3660 gnd.n3241 gnd.n3240 585
R3661 gnd.n3240 gnd.n3239 585
R3662 gnd.n2493 gnd.n1317 585
R3663 gnd.n4514 gnd.n1317 585
R3664 gnd.n2942 gnd.n2941 585
R3665 gnd.n2943 gnd.n2942 585
R3666 gnd.n2587 gnd.n1306 585
R3667 gnd.n4520 gnd.n1306 585
R3668 gnd.n2936 gnd.n2935 585
R3669 gnd.n2935 gnd.n2934 585
R3670 gnd.n2933 gnd.n1295 585
R3671 gnd.n4526 gnd.n1295 585
R3672 gnd.n2932 gnd.n2931 585
R3673 gnd.n2931 gnd.n2930 585
R3674 gnd.n2589 gnd.n1285 585
R3675 gnd.n4532 gnd.n1285 585
R3676 gnd.n2925 gnd.n2924 585
R3677 gnd.n2924 gnd.n2923 585
R3678 gnd.n2922 gnd.n1274 585
R3679 gnd.n4538 gnd.n1274 585
R3680 gnd.n2921 gnd.n2577 585
R3681 gnd.n2960 gnd.n2577 585
R3682 gnd.n2591 gnd.n1264 585
R3683 gnd.n4544 gnd.n1264 585
R3684 gnd.n2917 gnd.n2916 585
R3685 gnd.n2916 gnd.n2915 585
R3686 gnd.n2593 gnd.n1253 585
R3687 gnd.n4550 gnd.n1253 585
R3688 gnd.n2864 gnd.n2597 585
R3689 gnd.n2907 gnd.n2597 585
R3690 gnd.n2865 gnd.n1243 585
R3691 gnd.n4556 gnd.n1243 585
R3692 gnd.n2867 gnd.n2866 585
R3693 gnd.n2868 gnd.n2867 585
R3694 gnd.n2633 gnd.n1235 585
R3695 gnd.n4563 gnd.n1235 585
R3696 gnd.n2858 gnd.n2629 585
R3697 gnd.n2876 gnd.n2629 585
R3698 gnd.n2857 gnd.n1226 585
R3699 gnd.n4569 gnd.n1226 585
R3700 gnd.n2856 gnd.n2855 585
R3701 gnd.n2855 gnd.n2854 585
R3702 gnd.n2635 gnd.n1218 585
R3703 gnd.n4576 gnd.n1218 585
R3704 gnd.n2846 gnd.n2619 585
R3705 gnd.n2887 gnd.n2619 585
R3706 gnd.n2845 gnd.n1205 585
R3707 gnd.n4582 gnd.n1205 585
R3708 gnd.n2844 gnd.n2612 585
R3709 gnd.n2893 gnd.n2612 585
R3710 gnd.n2639 gnd.n2638 585
R3711 gnd.n2638 gnd.n2611 585
R3712 gnd.n2840 gnd.n1194 585
R3713 gnd.n4590 gnd.n1194 585
R3714 gnd.n2839 gnd.n2838 585
R3715 gnd.n2838 gnd.n2837 585
R3716 gnd.n2641 gnd.n1184 585
R3717 gnd.n4596 gnd.n1184 585
R3718 gnd.n2824 gnd.n2823 585
R3719 gnd.n2825 gnd.n2824 585
R3720 gnd.n2645 gnd.n1173 585
R3721 gnd.n4602 gnd.n1173 585
R3722 gnd.n2818 gnd.n2817 585
R3723 gnd.n2817 gnd.n2816 585
R3724 gnd.n2647 gnd.n1163 585
R3725 gnd.n4608 gnd.n1163 585
R3726 gnd.n2807 gnd.n2806 585
R3727 gnd.n2808 gnd.n2807 585
R3728 gnd.n2652 gnd.n1152 585
R3729 gnd.n4614 gnd.n1152 585
R3730 gnd.n2802 gnd.n2801 585
R3731 gnd.n2801 gnd.n2800 585
R3732 gnd.n2654 gnd.n1143 585
R3733 gnd.n4620 gnd.n1143 585
R3734 gnd.n2746 gnd.n2745 585
R3735 gnd.n2747 gnd.n2746 585
R3736 gnd.n2738 gnd.n1131 585
R3737 gnd.n4626 gnd.n1131 585
R3738 gnd.n2741 gnd.n2668 585
R3739 gnd.n2753 gnd.n2668 585
R3740 gnd.n2740 gnd.n1117 585
R3741 gnd.n2667 gnd.n1117 585
R3742 gnd.n4636 gnd.n1118 585
R3743 gnd.n4636 gnd.n4635 585
R3744 gnd.n7325 gnd.n7324 585
R3745 gnd.n7326 gnd.n7325 585
R3746 gnd.n87 gnd.n85 585
R3747 gnd.n7247 gnd.n85 585
R3748 gnd.n7169 gnd.n174 585
R3749 gnd.n174 gnd.n173 585
R3750 gnd.n7171 gnd.n7170 585
R3751 gnd.n7172 gnd.n7171 585
R3752 gnd.n175 gnd.n172 585
R3753 gnd.n7059 gnd.n172 585
R3754 gnd.n7164 gnd.n7163 585
R3755 gnd.n7163 gnd.n7162 585
R3756 gnd.n178 gnd.n177 585
R3757 gnd.n7065 gnd.n178 585
R3758 gnd.n7153 gnd.n7152 585
R3759 gnd.n7154 gnd.n7153 585
R3760 gnd.n191 gnd.n190 585
R3761 gnd.n7048 gnd.n190 585
R3762 gnd.n7148 gnd.n7147 585
R3763 gnd.n7147 gnd.n7146 585
R3764 gnd.n194 gnd.n193 585
R3765 gnd.n7074 gnd.n194 585
R3766 gnd.n7137 gnd.n7136 585
R3767 gnd.n7138 gnd.n7137 585
R3768 gnd.n207 gnd.n206 585
R3769 gnd.n7078 gnd.n206 585
R3770 gnd.n7132 gnd.n7131 585
R3771 gnd.n7131 gnd.n7130 585
R3772 gnd.n210 gnd.n209 585
R3773 gnd.n7084 gnd.n210 585
R3774 gnd.n7121 gnd.n7120 585
R3775 gnd.n7122 gnd.n7121 585
R3776 gnd.n223 gnd.n222 585
R3777 gnd.n4282 gnd.n222 585
R3778 gnd.n7097 gnd.n7096 585
R3779 gnd.n7098 gnd.n7097 585
R3780 gnd.n7095 gnd.n254 585
R3781 gnd.n7095 gnd.n7094 585
R3782 gnd.n253 gnd.n252 585
R3783 gnd.n4290 gnd.n252 585
R3784 gnd.n1515 gnd.n1514 585
R3785 gnd.n1518 gnd.n1514 585
R3786 gnd.n4310 gnd.n1516 585
R3787 gnd.n4310 gnd.n4309 585
R3788 gnd.n4313 gnd.n4312 585
R3789 gnd.n4314 gnd.n4313 585
R3790 gnd.n4311 gnd.n232 585
R3791 gnd.n4298 gnd.n232 585
R3792 gnd.n7115 gnd.n7114 585
R3793 gnd.n7114 gnd.n7113 585
R3794 gnd.n7116 gnd.n231 585
R3795 gnd.n4268 gnd.n231 585
R3796 gnd.n4328 gnd.n230 585
R3797 gnd.n4329 gnd.n4328 585
R3798 gnd.n4327 gnd.n1501 585
R3799 gnd.n4327 gnd.n4326 585
R3800 gnd.n4257 gnd.n1500 585
R3801 gnd.n1532 gnd.n1500 585
R3802 gnd.n4259 gnd.n4258 585
R3803 gnd.n4260 gnd.n4259 585
R3804 gnd.n1535 gnd.n1534 585
R3805 gnd.n4213 gnd.n1534 585
R3806 gnd.n4252 gnd.n4251 585
R3807 gnd.n4251 gnd.n4250 585
R3808 gnd.n1538 gnd.n1537 585
R3809 gnd.n4222 gnd.n1538 585
R3810 gnd.n4204 gnd.n1559 585
R3811 gnd.n4164 gnd.n1559 585
R3812 gnd.n4206 gnd.n4205 585
R3813 gnd.n4207 gnd.n4206 585
R3814 gnd.n1560 gnd.n1558 585
R3815 gnd.n1568 gnd.n1558 585
R3816 gnd.n4199 gnd.n4198 585
R3817 gnd.n4198 gnd.n4197 585
R3818 gnd.n1563 gnd.n1562 585
R3819 gnd.n4185 gnd.n1563 585
R3820 gnd.n1585 gnd.n1584 585
R3821 gnd.n1586 gnd.n1585 585
R3822 gnd.n1470 gnd.n1469 585
R3823 gnd.n4176 gnd.n1470 585
R3824 gnd.n4357 gnd.n4356 585
R3825 gnd.n4356 gnd.n4355 585
R3826 gnd.n4358 gnd.n1465 585
R3827 gnd.n4148 gnd.n1465 585
R3828 gnd.n4360 gnd.n4359 585
R3829 gnd.n4361 gnd.n4360 585
R3830 gnd.n1840 gnd.n1464 585
R3831 gnd.n1843 gnd.n1842 585
R3832 gnd.n1838 gnd.n1837 585
R3833 gnd.n1837 gnd.n1451 585
R3834 gnd.n1848 gnd.n1847 585
R3835 gnd.n1850 gnd.n1836 585
R3836 gnd.n1853 gnd.n1852 585
R3837 gnd.n1834 gnd.n1833 585
R3838 gnd.n1858 gnd.n1857 585
R3839 gnd.n1860 gnd.n1832 585
R3840 gnd.n1863 gnd.n1862 585
R3841 gnd.n1830 gnd.n1829 585
R3842 gnd.n1869 gnd.n1868 585
R3843 gnd.n1871 gnd.n1828 585
R3844 gnd.n1872 gnd.n1825 585
R3845 gnd.n1875 gnd.n1874 585
R3846 gnd.n1827 gnd.n1822 585
R3847 gnd.n1956 gnd.n1955 585
R3848 gnd.n1953 gnd.n1882 585
R3849 gnd.n1951 gnd.n1950 585
R3850 gnd.n1949 gnd.n1883 585
R3851 gnd.n1948 gnd.n1947 585
R3852 gnd.n1945 gnd.n1888 585
R3853 gnd.n1943 gnd.n1942 585
R3854 gnd.n1941 gnd.n1889 585
R3855 gnd.n1940 gnd.n1939 585
R3856 gnd.n1937 gnd.n1894 585
R3857 gnd.n1935 gnd.n1934 585
R3858 gnd.n1933 gnd.n1895 585
R3859 gnd.n1932 gnd.n1931 585
R3860 gnd.n1929 gnd.n1900 585
R3861 gnd.n1927 gnd.n1926 585
R3862 gnd.n1925 gnd.n1901 585
R3863 gnd.n1924 gnd.n1923 585
R3864 gnd.n1921 gnd.n1906 585
R3865 gnd.n1919 gnd.n1918 585
R3866 gnd.n1910 gnd.n1907 585
R3867 gnd.n1914 gnd.n1913 585
R3868 gnd.n156 gnd.n155 585
R3869 gnd.n7254 gnd.n151 585
R3870 gnd.n7256 gnd.n7255 585
R3871 gnd.n7258 gnd.n149 585
R3872 gnd.n7260 gnd.n7259 585
R3873 gnd.n7261 gnd.n144 585
R3874 gnd.n7263 gnd.n7262 585
R3875 gnd.n7265 gnd.n142 585
R3876 gnd.n7267 gnd.n7266 585
R3877 gnd.n7268 gnd.n137 585
R3878 gnd.n7270 gnd.n7269 585
R3879 gnd.n7272 gnd.n135 585
R3880 gnd.n7274 gnd.n7273 585
R3881 gnd.n7275 gnd.n130 585
R3882 gnd.n7277 gnd.n7276 585
R3883 gnd.n7279 gnd.n128 585
R3884 gnd.n7281 gnd.n7280 585
R3885 gnd.n7282 gnd.n123 585
R3886 gnd.n7284 gnd.n7283 585
R3887 gnd.n7286 gnd.n121 585
R3888 gnd.n7288 gnd.n7287 585
R3889 gnd.n7292 gnd.n116 585
R3890 gnd.n7294 gnd.n7293 585
R3891 gnd.n7296 gnd.n114 585
R3892 gnd.n7298 gnd.n7297 585
R3893 gnd.n7299 gnd.n109 585
R3894 gnd.n7301 gnd.n7300 585
R3895 gnd.n7303 gnd.n107 585
R3896 gnd.n7305 gnd.n7304 585
R3897 gnd.n7306 gnd.n102 585
R3898 gnd.n7308 gnd.n7307 585
R3899 gnd.n7310 gnd.n100 585
R3900 gnd.n7312 gnd.n7311 585
R3901 gnd.n7313 gnd.n95 585
R3902 gnd.n7315 gnd.n7314 585
R3903 gnd.n7317 gnd.n92 585
R3904 gnd.n7319 gnd.n7318 585
R3905 gnd.n7320 gnd.n90 585
R3906 gnd.n7321 gnd.n86 585
R3907 gnd.n94 gnd.n86 585
R3908 gnd.n7250 gnd.n82 585
R3909 gnd.n7326 gnd.n82 585
R3910 gnd.n7249 gnd.n7248 585
R3911 gnd.n7248 gnd.n7247 585
R3912 gnd.n161 gnd.n160 585
R3913 gnd.n173 gnd.n161 585
R3914 gnd.n7058 gnd.n170 585
R3915 gnd.n7172 gnd.n170 585
R3916 gnd.n7061 gnd.n7060 585
R3917 gnd.n7060 gnd.n7059 585
R3918 gnd.n7062 gnd.n180 585
R3919 gnd.n7162 gnd.n180 585
R3920 gnd.n7064 gnd.n7063 585
R3921 gnd.n7065 gnd.n7064 585
R3922 gnd.n7046 gnd.n189 585
R3923 gnd.n7154 gnd.n189 585
R3924 gnd.n7050 gnd.n7049 585
R3925 gnd.n7049 gnd.n7048 585
R3926 gnd.n269 gnd.n195 585
R3927 gnd.n7146 gnd.n195 585
R3928 gnd.n7076 gnd.n7075 585
R3929 gnd.n7075 gnd.n7074 585
R3930 gnd.n7077 gnd.n204 585
R3931 gnd.n7138 gnd.n204 585
R3932 gnd.n7080 gnd.n7079 585
R3933 gnd.n7079 gnd.n7078 585
R3934 gnd.n7081 gnd.n212 585
R3935 gnd.n7130 gnd.n212 585
R3936 gnd.n7083 gnd.n7082 585
R3937 gnd.n7084 gnd.n7083 585
R3938 gnd.n263 gnd.n221 585
R3939 gnd.n7122 gnd.n221 585
R3940 gnd.n4284 gnd.n4283 585
R3941 gnd.n4283 gnd.n4282 585
R3942 gnd.n4285 gnd.n249 585
R3943 gnd.n7098 gnd.n249 585
R3944 gnd.n4286 gnd.n256 585
R3945 gnd.n7094 gnd.n256 585
R3946 gnd.n4291 gnd.n4287 585
R3947 gnd.n4291 gnd.n4290 585
R3948 gnd.n4293 gnd.n4292 585
R3949 gnd.n4292 gnd.n1518 585
R3950 gnd.n4294 gnd.n1517 585
R3951 gnd.n4309 gnd.n1517 585
R3952 gnd.n4295 gnd.n1512 585
R3953 gnd.n4314 gnd.n1512 585
R3954 gnd.n4297 gnd.n4296 585
R3955 gnd.n4298 gnd.n4297 585
R3956 gnd.n1523 gnd.n234 585
R3957 gnd.n7113 gnd.n234 585
R3958 gnd.n4270 gnd.n4269 585
R3959 gnd.n4269 gnd.n4268 585
R3960 gnd.n4267 gnd.n1497 585
R3961 gnd.n4329 gnd.n1497 585
R3962 gnd.n4266 gnd.n1503 585
R3963 gnd.n4326 gnd.n1503 585
R3964 gnd.n1529 gnd.n1525 585
R3965 gnd.n1532 gnd.n1529 585
R3966 gnd.n4262 gnd.n4261 585
R3967 gnd.n4261 gnd.n4260 585
R3968 gnd.n1528 gnd.n1527 585
R3969 gnd.n4213 gnd.n1528 585
R3970 gnd.n4162 gnd.n1540 585
R3971 gnd.n4250 gnd.n1540 585
R3972 gnd.n4163 gnd.n1548 585
R3973 gnd.n4222 gnd.n1548 585
R3974 gnd.n4166 gnd.n4165 585
R3975 gnd.n4165 gnd.n4164 585
R3976 gnd.n4167 gnd.n1556 585
R3977 gnd.n4207 gnd.n1556 585
R3978 gnd.n4169 gnd.n4168 585
R3979 gnd.n4168 gnd.n1568 585
R3980 gnd.n4170 gnd.n1565 585
R3981 gnd.n4197 gnd.n1565 585
R3982 gnd.n4171 gnd.n1587 585
R3983 gnd.n4185 gnd.n1587 585
R3984 gnd.n4172 gnd.n1593 585
R3985 gnd.n1593 gnd.n1586 585
R3986 gnd.n4174 gnd.n4173 585
R3987 gnd.n4176 gnd.n4174 585
R3988 gnd.n1594 gnd.n1472 585
R3989 gnd.n4355 gnd.n1472 585
R3990 gnd.n4150 gnd.n4149 585
R3991 gnd.n4149 gnd.n4148 585
R3992 gnd.n1596 gnd.n1460 585
R3993 gnd.n4361 gnd.n1460 585
R3994 gnd.n3976 gnd.n1967 585
R3995 gnd.n1967 gnd.n1786 585
R3996 gnd.n3978 gnd.n3977 585
R3997 gnd.n3979 gnd.n3978 585
R3998 gnd.n3887 gnd.n1966 585
R3999 gnd.n3850 gnd.n1966 585
R4000 gnd.n3886 gnd.n3885 585
R4001 gnd.n3885 gnd.n3884 585
R4002 gnd.n1969 gnd.n1968 585
R4003 gnd.n3847 gnd.n1969 585
R4004 gnd.n3867 gnd.n3866 585
R4005 gnd.n3868 gnd.n3867 585
R4006 gnd.n3865 gnd.n1980 585
R4007 gnd.n1980 gnd.n1977 585
R4008 gnd.n3864 gnd.n3863 585
R4009 gnd.n3863 gnd.n3862 585
R4010 gnd.n1982 gnd.n1981 585
R4011 gnd.n3836 gnd.n1982 585
R4012 gnd.n3819 gnd.n3818 585
R4013 gnd.n3818 gnd.n1993 585
R4014 gnd.n3820 gnd.n2004 585
R4015 gnd.n3804 gnd.n2004 585
R4016 gnd.n3822 gnd.n3821 585
R4017 gnd.n3823 gnd.n3822 585
R4018 gnd.n3817 gnd.n2003 585
R4019 gnd.n2003 gnd.n1999 585
R4020 gnd.n3816 gnd.n3815 585
R4021 gnd.n3815 gnd.n3814 585
R4022 gnd.n2006 gnd.n2005 585
R4023 gnd.n3795 gnd.n2006 585
R4024 gnd.n3779 gnd.n3778 585
R4025 gnd.n3778 gnd.n2015 585
R4026 gnd.n3780 gnd.n2025 585
R4027 gnd.n3765 gnd.n2025 585
R4028 gnd.n3782 gnd.n3781 585
R4029 gnd.n3783 gnd.n3782 585
R4030 gnd.n3777 gnd.n2024 585
R4031 gnd.n2024 gnd.n2021 585
R4032 gnd.n3776 gnd.n3775 585
R4033 gnd.n3775 gnd.t173 585
R4034 gnd.n2027 gnd.n2026 585
R4035 gnd.n3756 gnd.n2027 585
R4036 gnd.n3740 gnd.n3739 585
R4037 gnd.n3739 gnd.n2038 585
R4038 gnd.n3741 gnd.n2048 585
R4039 gnd.n3725 gnd.n2048 585
R4040 gnd.n3743 gnd.n3742 585
R4041 gnd.n3744 gnd.n3743 585
R4042 gnd.n3738 gnd.n2047 585
R4043 gnd.n2047 gnd.n2044 585
R4044 gnd.n3737 gnd.n3736 585
R4045 gnd.n3736 gnd.n3735 585
R4046 gnd.n2050 gnd.n2049 585
R4047 gnd.n3716 gnd.n2050 585
R4048 gnd.n3700 gnd.n3699 585
R4049 gnd.n3699 gnd.n2061 585
R4050 gnd.n3701 gnd.n2070 585
R4051 gnd.n3686 gnd.n2070 585
R4052 gnd.n3703 gnd.n3702 585
R4053 gnd.n3704 gnd.n3703 585
R4054 gnd.n3698 gnd.n2069 585
R4055 gnd.n3692 gnd.n2069 585
R4056 gnd.n3697 gnd.n3696 585
R4057 gnd.n3696 gnd.n3695 585
R4058 gnd.n2072 gnd.n2071 585
R4059 gnd.n3645 gnd.n2072 585
R4060 gnd.n3673 gnd.n3672 585
R4061 gnd.n3674 gnd.n3673 585
R4062 gnd.n3671 gnd.n2085 585
R4063 gnd.n3666 gnd.n2085 585
R4064 gnd.n3670 gnd.n3669 585
R4065 gnd.n3669 gnd.n3668 585
R4066 gnd.n2087 gnd.n2086 585
R4067 gnd.n3653 gnd.n2087 585
R4068 gnd.n3638 gnd.n2106 585
R4069 gnd.n2106 gnd.n2097 585
R4070 gnd.n3640 gnd.n3639 585
R4071 gnd.n3641 gnd.n3640 585
R4072 gnd.n3637 gnd.n2105 585
R4073 gnd.n2111 gnd.n2105 585
R4074 gnd.n3636 gnd.n3635 585
R4075 gnd.n3635 gnd.n3634 585
R4076 gnd.n2108 gnd.n2107 585
R4077 gnd.n3375 gnd.n2108 585
R4078 gnd.n3623 gnd.n3622 585
R4079 gnd.n3624 gnd.n3623 585
R4080 gnd.n3621 gnd.n2121 585
R4081 gnd.n2121 gnd.n2118 585
R4082 gnd.n3620 gnd.n3619 585
R4083 gnd.n3619 gnd.n3618 585
R4084 gnd.n2123 gnd.n2122 585
R4085 gnd.n3383 gnd.n2123 585
R4086 gnd.n3591 gnd.n3590 585
R4087 gnd.n3592 gnd.n3591 585
R4088 gnd.n3589 gnd.n2136 585
R4089 gnd.n2136 gnd.n2133 585
R4090 gnd.n3588 gnd.n3587 585
R4091 gnd.n3587 gnd.n3586 585
R4092 gnd.n2138 gnd.n2137 585
R4093 gnd.n3390 gnd.n2138 585
R4094 gnd.n3572 gnd.n3571 585
R4095 gnd.n3573 gnd.n3572 585
R4096 gnd.n3570 gnd.n2150 585
R4097 gnd.n3565 gnd.n2150 585
R4098 gnd.n3569 gnd.n3568 585
R4099 gnd.n3568 gnd.n3567 585
R4100 gnd.n2152 gnd.n2151 585
R4101 gnd.n3554 gnd.n2152 585
R4102 gnd.n3540 gnd.n2174 585
R4103 gnd.n2174 gnd.n2163 585
R4104 gnd.n3542 gnd.n3541 585
R4105 gnd.n3543 gnd.n3542 585
R4106 gnd.n3539 gnd.n2173 585
R4107 gnd.n2173 gnd.n2170 585
R4108 gnd.n3538 gnd.n3537 585
R4109 gnd.n3537 gnd.n3536 585
R4110 gnd.n2176 gnd.n2175 585
R4111 gnd.n3404 gnd.n2176 585
R4112 gnd.n3525 gnd.n3524 585
R4113 gnd.n3526 gnd.n3525 585
R4114 gnd.n3523 gnd.n2187 585
R4115 gnd.n2187 gnd.n2184 585
R4116 gnd.n3522 gnd.n3521 585
R4117 gnd.n3521 gnd.n3520 585
R4118 gnd.n2189 gnd.n2188 585
R4119 gnd.t156 gnd.n2189 585
R4120 gnd.n3507 gnd.n3506 585
R4121 gnd.n3508 gnd.n3507 585
R4122 gnd.n3505 gnd.n2202 585
R4123 gnd.n2202 gnd.n2199 585
R4124 gnd.n3504 gnd.n3503 585
R4125 gnd.n3503 gnd.n3502 585
R4126 gnd.n2204 gnd.n2203 585
R4127 gnd.n2215 gnd.n2204 585
R4128 gnd.n3476 gnd.n3475 585
R4129 gnd.n3475 gnd.n2214 585
R4130 gnd.n3477 gnd.n2224 585
R4131 gnd.n3422 gnd.n2224 585
R4132 gnd.n3479 gnd.n3478 585
R4133 gnd.n3480 gnd.n3479 585
R4134 gnd.n3474 gnd.n2223 585
R4135 gnd.n3469 gnd.n2223 585
R4136 gnd.n3473 gnd.n3472 585
R4137 gnd.n3472 gnd.n3471 585
R4138 gnd.n2226 gnd.n2225 585
R4139 gnd.n2236 gnd.n2226 585
R4140 gnd.n3445 gnd.n3444 585
R4141 gnd.n3444 gnd.n2234 585
R4142 gnd.n3446 gnd.n2246 585
R4143 gnd.n3432 gnd.n2246 585
R4144 gnd.n3448 gnd.n3447 585
R4145 gnd.n3449 gnd.n3448 585
R4146 gnd.n3443 gnd.n2245 585
R4147 gnd.n3438 gnd.n2245 585
R4148 gnd.n3442 gnd.n3441 585
R4149 gnd.n3441 gnd.n3440 585
R4150 gnd.n2248 gnd.n2247 585
R4151 gnd.n3367 gnd.n2248 585
R4152 gnd.n3354 gnd.n2266 585
R4153 gnd.n2266 gnd.n2265 585
R4154 gnd.n3356 gnd.n3355 585
R4155 gnd.n3357 gnd.n3356 585
R4156 gnd.n3353 gnd.n2264 585
R4157 gnd.n2264 gnd.n2260 585
R4158 gnd.n3351 gnd.n3350 585
R4159 gnd.n2288 gnd.n2287 585
R4160 gnd.n3347 gnd.n3346 585
R4161 gnd.n3348 gnd.n3347 585
R4162 gnd.n3345 gnd.n2323 585
R4163 gnd.n3344 gnd.n3343 585
R4164 gnd.n3342 gnd.n3341 585
R4165 gnd.n3340 gnd.n3339 585
R4166 gnd.n3338 gnd.n3337 585
R4167 gnd.n3336 gnd.n3335 585
R4168 gnd.n3334 gnd.n3333 585
R4169 gnd.n3332 gnd.n3331 585
R4170 gnd.n3330 gnd.n3329 585
R4171 gnd.n3328 gnd.n3327 585
R4172 gnd.n3326 gnd.n3325 585
R4173 gnd.n3324 gnd.n3323 585
R4174 gnd.n3322 gnd.n3321 585
R4175 gnd.n3320 gnd.n3319 585
R4176 gnd.n3318 gnd.n3317 585
R4177 gnd.n3316 gnd.n3315 585
R4178 gnd.n3314 gnd.n3313 585
R4179 gnd.n3312 gnd.n3311 585
R4180 gnd.n3310 gnd.n3309 585
R4181 gnd.n3308 gnd.n3307 585
R4182 gnd.n3306 gnd.n3305 585
R4183 gnd.n3304 gnd.n3303 585
R4184 gnd.n3302 gnd.n3301 585
R4185 gnd.n3300 gnd.n3299 585
R4186 gnd.n3298 gnd.n3297 585
R4187 gnd.n3296 gnd.n3295 585
R4188 gnd.n3294 gnd.n3293 585
R4189 gnd.n3292 gnd.n3291 585
R4190 gnd.n3290 gnd.n3289 585
R4191 gnd.n3288 gnd.n3287 585
R4192 gnd.n3286 gnd.n2395 585
R4193 gnd.n2394 gnd.n2393 585
R4194 gnd.n2392 gnd.n2391 585
R4195 gnd.n2389 gnd.n2388 585
R4196 gnd.n2387 gnd.n2386 585
R4197 gnd.n2385 gnd.n2384 585
R4198 gnd.n2383 gnd.n2382 585
R4199 gnd.n2381 gnd.n2380 585
R4200 gnd.n2379 gnd.n2378 585
R4201 gnd.n2377 gnd.n2376 585
R4202 gnd.n2375 gnd.n2374 585
R4203 gnd.n2373 gnd.n2372 585
R4204 gnd.n2371 gnd.n2370 585
R4205 gnd.n2369 gnd.n2368 585
R4206 gnd.n2367 gnd.n2366 585
R4207 gnd.n2365 gnd.n2364 585
R4208 gnd.n2363 gnd.n2362 585
R4209 gnd.n2361 gnd.n2360 585
R4210 gnd.n2359 gnd.n2358 585
R4211 gnd.n2357 gnd.n2356 585
R4212 gnd.n2355 gnd.n2354 585
R4213 gnd.n2353 gnd.n2352 585
R4214 gnd.n2351 gnd.n2350 585
R4215 gnd.n2349 gnd.n2348 585
R4216 gnd.n2347 gnd.n2346 585
R4217 gnd.n2345 gnd.n2344 585
R4218 gnd.n2343 gnd.n2342 585
R4219 gnd.n2341 gnd.n2340 585
R4220 gnd.n2339 gnd.n2338 585
R4221 gnd.n2337 gnd.n2336 585
R4222 gnd.n2335 gnd.n2334 585
R4223 gnd.n2333 gnd.n2332 585
R4224 gnd.n3983 gnd.n3982 585
R4225 gnd.n3985 gnd.n3984 585
R4226 gnd.n3987 gnd.n3986 585
R4227 gnd.n3989 gnd.n3988 585
R4228 gnd.n3991 gnd.n3990 585
R4229 gnd.n3993 gnd.n3992 585
R4230 gnd.n3995 gnd.n3994 585
R4231 gnd.n3997 gnd.n3996 585
R4232 gnd.n3999 gnd.n3998 585
R4233 gnd.n4001 gnd.n4000 585
R4234 gnd.n4003 gnd.n4002 585
R4235 gnd.n4005 gnd.n4004 585
R4236 gnd.n4007 gnd.n4006 585
R4237 gnd.n4009 gnd.n4008 585
R4238 gnd.n4011 gnd.n4010 585
R4239 gnd.n4013 gnd.n4012 585
R4240 gnd.n4015 gnd.n4014 585
R4241 gnd.n4017 gnd.n4016 585
R4242 gnd.n4019 gnd.n4018 585
R4243 gnd.n4021 gnd.n4020 585
R4244 gnd.n4023 gnd.n4022 585
R4245 gnd.n4025 gnd.n4024 585
R4246 gnd.n4027 gnd.n4026 585
R4247 gnd.n4029 gnd.n4028 585
R4248 gnd.n4031 gnd.n4030 585
R4249 gnd.n4033 gnd.n4032 585
R4250 gnd.n4035 gnd.n4034 585
R4251 gnd.n4037 gnd.n4036 585
R4252 gnd.n4039 gnd.n4038 585
R4253 gnd.n4042 gnd.n4041 585
R4254 gnd.n4044 gnd.n4043 585
R4255 gnd.n4046 gnd.n4045 585
R4256 gnd.n4048 gnd.n4047 585
R4257 gnd.n3909 gnd.n1958 585
R4258 gnd.n3911 gnd.n3910 585
R4259 gnd.n3913 gnd.n3912 585
R4260 gnd.n3915 gnd.n3914 585
R4261 gnd.n3918 gnd.n3917 585
R4262 gnd.n3920 gnd.n3919 585
R4263 gnd.n3922 gnd.n3921 585
R4264 gnd.n3924 gnd.n3923 585
R4265 gnd.n3926 gnd.n3925 585
R4266 gnd.n3928 gnd.n3927 585
R4267 gnd.n3930 gnd.n3929 585
R4268 gnd.n3932 gnd.n3931 585
R4269 gnd.n3934 gnd.n3933 585
R4270 gnd.n3936 gnd.n3935 585
R4271 gnd.n3938 gnd.n3937 585
R4272 gnd.n3940 gnd.n3939 585
R4273 gnd.n3942 gnd.n3941 585
R4274 gnd.n3944 gnd.n3943 585
R4275 gnd.n3946 gnd.n3945 585
R4276 gnd.n3948 gnd.n3947 585
R4277 gnd.n3950 gnd.n3949 585
R4278 gnd.n3952 gnd.n3951 585
R4279 gnd.n3954 gnd.n3953 585
R4280 gnd.n3956 gnd.n3955 585
R4281 gnd.n3958 gnd.n3957 585
R4282 gnd.n3960 gnd.n3959 585
R4283 gnd.n3962 gnd.n3961 585
R4284 gnd.n3964 gnd.n3963 585
R4285 gnd.n3966 gnd.n3965 585
R4286 gnd.n3968 gnd.n3967 585
R4287 gnd.n3970 gnd.n3969 585
R4288 gnd.n3972 gnd.n3971 585
R4289 gnd.n3974 gnd.n3973 585
R4290 gnd.n3981 gnd.n1961 585
R4291 gnd.n3981 gnd.n1786 585
R4292 gnd.n3980 gnd.n1963 585
R4293 gnd.n3980 gnd.n3979 585
R4294 gnd.n3843 gnd.n1962 585
R4295 gnd.n3850 gnd.n1962 585
R4296 gnd.n3844 gnd.n1970 585
R4297 gnd.n3884 gnd.n1970 585
R4298 gnd.n3846 gnd.n3845 585
R4299 gnd.n3847 gnd.n3846 585
R4300 gnd.n3842 gnd.n1979 585
R4301 gnd.n3868 gnd.n1979 585
R4302 gnd.n3841 gnd.n3840 585
R4303 gnd.n3840 gnd.n1977 585
R4304 gnd.n3839 gnd.n1984 585
R4305 gnd.n3862 gnd.n1984 585
R4306 gnd.n3838 gnd.n3837 585
R4307 gnd.n3837 gnd.n3836 585
R4308 gnd.n1992 gnd.n1991 585
R4309 gnd.n1993 gnd.n1992 585
R4310 gnd.n3803 gnd.n3802 585
R4311 gnd.n3804 gnd.n3803 585
R4312 gnd.n3801 gnd.n2001 585
R4313 gnd.n3823 gnd.n2001 585
R4314 gnd.n3800 gnd.n3799 585
R4315 gnd.n3799 gnd.n1999 585
R4316 gnd.n3798 gnd.n2008 585
R4317 gnd.n3814 gnd.n2008 585
R4318 gnd.n3797 gnd.n3796 585
R4319 gnd.n3796 gnd.n3795 585
R4320 gnd.n2014 gnd.n2013 585
R4321 gnd.n2015 gnd.n2014 585
R4322 gnd.n3764 gnd.n3763 585
R4323 gnd.n3765 gnd.n3764 585
R4324 gnd.n3762 gnd.n2022 585
R4325 gnd.n3783 gnd.n2022 585
R4326 gnd.n3761 gnd.n3760 585
R4327 gnd.n3760 gnd.n2021 585
R4328 gnd.n3759 gnd.n2029 585
R4329 gnd.t173 gnd.n2029 585
R4330 gnd.n3758 gnd.n3757 585
R4331 gnd.n3757 gnd.n3756 585
R4332 gnd.n2037 gnd.n2036 585
R4333 gnd.n2038 gnd.n2037 585
R4334 gnd.n3724 gnd.n3723 585
R4335 gnd.n3725 gnd.n3724 585
R4336 gnd.n3722 gnd.n2045 585
R4337 gnd.n3744 gnd.n2045 585
R4338 gnd.n3721 gnd.n3720 585
R4339 gnd.n3720 gnd.n2044 585
R4340 gnd.n3719 gnd.n2052 585
R4341 gnd.n3735 gnd.n2052 585
R4342 gnd.n3718 gnd.n3717 585
R4343 gnd.n3717 gnd.n3716 585
R4344 gnd.n2060 gnd.n2059 585
R4345 gnd.n2061 gnd.n2060 585
R4346 gnd.n3688 gnd.n3687 585
R4347 gnd.n3687 gnd.n3686 585
R4348 gnd.n3689 gnd.n2067 585
R4349 gnd.n3704 gnd.n2067 585
R4350 gnd.n3691 gnd.n3690 585
R4351 gnd.n3692 gnd.n3691 585
R4352 gnd.n2077 gnd.n2075 585
R4353 gnd.n3695 gnd.n2075 585
R4354 gnd.n3647 gnd.n3646 585
R4355 gnd.n3646 gnd.n3645 585
R4356 gnd.n3648 gnd.n2083 585
R4357 gnd.n3674 gnd.n2083 585
R4358 gnd.n3649 gnd.n2090 585
R4359 gnd.n3666 gnd.n2090 585
R4360 gnd.n3650 gnd.n2089 585
R4361 gnd.n3668 gnd.n2089 585
R4362 gnd.n3652 gnd.n3651 585
R4363 gnd.n3653 gnd.n3652 585
R4364 gnd.n3644 gnd.n2099 585
R4365 gnd.n2099 gnd.n2097 585
R4366 gnd.n3643 gnd.n3642 585
R4367 gnd.n3642 gnd.n3641 585
R4368 gnd.n2101 gnd.n2100 585
R4369 gnd.n2111 gnd.n2101 585
R4370 gnd.n3373 gnd.n2110 585
R4371 gnd.n3634 gnd.n2110 585
R4372 gnd.n3377 gnd.n3376 585
R4373 gnd.n3376 gnd.n3375 585
R4374 gnd.n3378 gnd.n2119 585
R4375 gnd.n3624 gnd.n2119 585
R4376 gnd.n3380 gnd.n3379 585
R4377 gnd.n3379 gnd.n2118 585
R4378 gnd.n3381 gnd.n2125 585
R4379 gnd.n3618 gnd.n2125 585
R4380 gnd.n3385 gnd.n3384 585
R4381 gnd.n3384 gnd.n3383 585
R4382 gnd.n3386 gnd.n2134 585
R4383 gnd.n3592 gnd.n2134 585
R4384 gnd.n3388 gnd.n3387 585
R4385 gnd.n3387 gnd.n2133 585
R4386 gnd.n3389 gnd.n2140 585
R4387 gnd.n3586 gnd.n2140 585
R4388 gnd.n3392 gnd.n3391 585
R4389 gnd.n3391 gnd.n3390 585
R4390 gnd.n3393 gnd.n2147 585
R4391 gnd.n3573 gnd.n2147 585
R4392 gnd.n3394 gnd.n2155 585
R4393 gnd.n3565 gnd.n2155 585
R4394 gnd.n3395 gnd.n2154 585
R4395 gnd.n3567 gnd.n2154 585
R4396 gnd.n3396 gnd.n2164 585
R4397 gnd.n3554 gnd.n2164 585
R4398 gnd.n3398 gnd.n3397 585
R4399 gnd.n3397 gnd.n2163 585
R4400 gnd.n3399 gnd.n2171 585
R4401 gnd.n3543 gnd.n2171 585
R4402 gnd.n3401 gnd.n3400 585
R4403 gnd.n3400 gnd.n2170 585
R4404 gnd.n3402 gnd.n2178 585
R4405 gnd.n3536 gnd.n2178 585
R4406 gnd.n3406 gnd.n3405 585
R4407 gnd.n3405 gnd.n3404 585
R4408 gnd.n3407 gnd.n2185 585
R4409 gnd.n3526 gnd.n2185 585
R4410 gnd.n3409 gnd.n3408 585
R4411 gnd.n3408 gnd.n2184 585
R4412 gnd.n3410 gnd.n2192 585
R4413 gnd.n3520 gnd.n2192 585
R4414 gnd.n3413 gnd.n3412 585
R4415 gnd.n3412 gnd.t156 585
R4416 gnd.n3414 gnd.n2200 585
R4417 gnd.n3508 gnd.n2200 585
R4418 gnd.n3416 gnd.n3415 585
R4419 gnd.n3415 gnd.n2199 585
R4420 gnd.n3417 gnd.n2206 585
R4421 gnd.n3502 gnd.n2206 585
R4422 gnd.n3419 gnd.n3418 585
R4423 gnd.n3419 gnd.n2215 585
R4424 gnd.n3420 gnd.n3372 585
R4425 gnd.n3420 gnd.n2214 585
R4426 gnd.n3424 gnd.n3423 585
R4427 gnd.n3423 gnd.n3422 585
R4428 gnd.n3425 gnd.n2221 585
R4429 gnd.n3480 gnd.n2221 585
R4430 gnd.n3426 gnd.n2228 585
R4431 gnd.n3469 gnd.n2228 585
R4432 gnd.n3427 gnd.n2227 585
R4433 gnd.n3471 gnd.n2227 585
R4434 gnd.n3429 gnd.n3428 585
R4435 gnd.n3429 gnd.n2236 585
R4436 gnd.n3430 gnd.n3371 585
R4437 gnd.n3430 gnd.n2234 585
R4438 gnd.n3434 gnd.n3433 585
R4439 gnd.n3433 gnd.n3432 585
R4440 gnd.n3435 gnd.n2243 585
R4441 gnd.n3449 gnd.n2243 585
R4442 gnd.n3437 gnd.n3436 585
R4443 gnd.n3438 gnd.n3437 585
R4444 gnd.n3370 gnd.n2250 585
R4445 gnd.n3440 gnd.n2250 585
R4446 gnd.n3369 gnd.n3368 585
R4447 gnd.n3368 gnd.n3367 585
R4448 gnd.n2252 gnd.n2251 585
R4449 gnd.n2265 gnd.n2252 585
R4450 gnd.n2329 gnd.n2262 585
R4451 gnd.n3357 gnd.n2262 585
R4452 gnd.n2331 gnd.n2330 585
R4453 gnd.n2331 gnd.n2260 585
R4454 gnd.n930 gnd.n929 585
R4455 gnd.n4740 gnd.n930 585
R4456 gnd.n7007 gnd.n7006 585
R4457 gnd.n7006 gnd.n7005 585
R4458 gnd.n7010 gnd.n321 585
R4459 gnd.n321 gnd.n320 585
R4460 gnd.n7012 gnd.n7011 585
R4461 gnd.n7013 gnd.n7012 585
R4462 gnd.n319 gnd.n318 585
R4463 gnd.n7014 gnd.n319 585
R4464 gnd.n7017 gnd.n7016 585
R4465 gnd.n7016 gnd.n7015 585
R4466 gnd.n7018 gnd.n313 585
R4467 gnd.n313 gnd.n312 585
R4468 gnd.n7020 gnd.n7019 585
R4469 gnd.n7021 gnd.n7020 585
R4470 gnd.n311 gnd.n310 585
R4471 gnd.n7022 gnd.n311 585
R4472 gnd.n7025 gnd.n7024 585
R4473 gnd.n7024 gnd.n7023 585
R4474 gnd.n7026 gnd.n302 585
R4475 gnd.n302 gnd.n301 585
R4476 gnd.n7028 gnd.n7027 585
R4477 gnd.n7029 gnd.n7028 585
R4478 gnd.n303 gnd.n299 585
R4479 gnd.n7030 gnd.n299 585
R4480 gnd.n7032 gnd.n300 585
R4481 gnd.n7032 gnd.n7031 585
R4482 gnd.n7034 gnd.n298 585
R4483 gnd.n7034 gnd.n7033 585
R4484 gnd.n7036 gnd.n7035 585
R4485 gnd.n7035 gnd.n83 585
R4486 gnd.n7037 gnd.n293 585
R4487 gnd.n293 gnd.n81 585
R4488 gnd.n7039 gnd.n7038 585
R4489 gnd.n7039 gnd.n162 585
R4490 gnd.n7040 gnd.n292 585
R4491 gnd.n7040 gnd.n171 585
R4492 gnd.n7042 gnd.n7041 585
R4493 gnd.n7041 gnd.n169 585
R4494 gnd.n7043 gnd.n287 585
R4495 gnd.n287 gnd.n182 585
R4496 gnd.n7045 gnd.n7044 585
R4497 gnd.n7045 gnd.n179 585
R4498 gnd.n7067 gnd.n286 585
R4499 gnd.n7067 gnd.n7066 585
R4500 gnd.n7069 gnd.n7068 585
R4501 gnd.n7068 gnd.n188 585
R4502 gnd.n7070 gnd.n271 585
R4503 gnd.n271 gnd.n197 585
R4504 gnd.n7072 gnd.n7071 585
R4505 gnd.n7073 gnd.n7072 585
R4506 gnd.n272 gnd.n270 585
R4507 gnd.n270 gnd.n205 585
R4508 gnd.n280 gnd.n279 585
R4509 gnd.n279 gnd.n203 585
R4510 gnd.n278 gnd.n277 585
R4511 gnd.n278 gnd.n214 585
R4512 gnd.n276 gnd.n262 585
R4513 gnd.n262 gnd.n211 585
R4514 gnd.n7086 gnd.n261 585
R4515 gnd.n7086 gnd.n7085 585
R4516 gnd.n7088 gnd.n7087 585
R4517 gnd.n7087 gnd.n220 585
R4518 gnd.n7089 gnd.n258 585
R4519 gnd.n258 gnd.n251 585
R4520 gnd.n7092 gnd.n7091 585
R4521 gnd.n7093 gnd.n7092 585
R4522 gnd.n259 gnd.n257 585
R4523 gnd.n257 gnd.n255 585
R4524 gnd.n4305 gnd.n1520 585
R4525 gnd.n4288 gnd.n1520 585
R4526 gnd.n4307 gnd.n4306 585
R4527 gnd.n4308 gnd.n4307 585
R4528 gnd.n4302 gnd.n1519 585
R4529 gnd.n1519 gnd.n1513 585
R4530 gnd.n4301 gnd.n4300 585
R4531 gnd.n4300 gnd.n4299 585
R4532 gnd.n4235 gnd.n1522 585
R4533 gnd.n1522 gnd.n236 585
R4534 gnd.n4237 gnd.n4236 585
R4535 gnd.n4236 gnd.n233 585
R4536 gnd.n4239 gnd.n4232 585
R4537 gnd.n4232 gnd.n1499 585
R4538 gnd.n4241 gnd.n4240 585
R4539 gnd.n4241 gnd.n1496 585
R4540 gnd.n4242 gnd.n4231 585
R4541 gnd.n4242 gnd.n1502 585
R4542 gnd.n4244 gnd.n4243 585
R4543 gnd.n4243 gnd.n1533 585
R4544 gnd.n4245 gnd.n1543 585
R4545 gnd.n1543 gnd.n1530 585
R4546 gnd.n4247 gnd.n4246 585
R4547 gnd.n4248 gnd.n4247 585
R4548 gnd.n1544 gnd.n1542 585
R4549 gnd.n1542 gnd.n1539 585
R4550 gnd.n4225 gnd.n4224 585
R4551 gnd.n4224 gnd.n4223 585
R4552 gnd.n1547 gnd.n1546 585
R4553 gnd.n1557 gnd.n1547 585
R4554 gnd.n4193 gnd.n1570 585
R4555 gnd.n1570 gnd.n1555 585
R4556 gnd.n4195 gnd.n4194 585
R4557 gnd.n4196 gnd.n4195 585
R4558 gnd.n1571 gnd.n1569 585
R4559 gnd.n1569 gnd.n1564 585
R4560 gnd.n4188 gnd.n4187 585
R4561 gnd.n4187 gnd.n4186 585
R4562 gnd.n1581 gnd.n1573 585
R4563 gnd.n4175 gnd.n1581 585
R4564 gnd.n1580 gnd.n1579 585
R4565 gnd.n1580 gnd.n1474 585
R4566 gnd.n1575 gnd.n1574 585
R4567 gnd.n1574 gnd.n1471 585
R4568 gnd.n1458 gnd.n1457 585
R4569 gnd.n1462 gnd.n1458 585
R4570 gnd.n4364 gnd.n4363 585
R4571 gnd.n4363 gnd.n4362 585
R4572 gnd.n4365 gnd.n1452 585
R4573 gnd.n1459 gnd.n1452 585
R4574 gnd.n4367 gnd.n4366 585
R4575 gnd.n4368 gnd.n4367 585
R4576 gnd.n1449 gnd.n1448 585
R4577 gnd.n4369 gnd.n1449 585
R4578 gnd.n4372 gnd.n4371 585
R4579 gnd.n4371 gnd.n4370 585
R4580 gnd.n4373 gnd.n1443 585
R4581 gnd.n1443 gnd.n1441 585
R4582 gnd.n4375 gnd.n4374 585
R4583 gnd.n4376 gnd.n4375 585
R4584 gnd.n1444 gnd.n1442 585
R4585 gnd.n1442 gnd.n1439 585
R4586 gnd.n4113 gnd.n4112 585
R4587 gnd.n4114 gnd.n4113 585
R4588 gnd.n1753 gnd.n1752 585
R4589 gnd.n4102 gnd.n1752 585
R4590 gnd.n4107 gnd.n4106 585
R4591 gnd.n4106 gnd.n4105 585
R4592 gnd.n1756 gnd.n1755 585
R4593 gnd.n4091 gnd.n1756 585
R4594 gnd.n4089 gnd.n4088 585
R4595 gnd.n4090 gnd.n4089 585
R4596 gnd.n1765 gnd.n1764 585
R4597 gnd.n4079 gnd.n1764 585
R4598 gnd.n4084 gnd.n4083 585
R4599 gnd.n4083 gnd.n4082 585
R4600 gnd.n1768 gnd.n1767 585
R4601 gnd.n4070 gnd.n1768 585
R4602 gnd.n4068 gnd.n4067 585
R4603 gnd.n4069 gnd.n4068 585
R4604 gnd.n1777 gnd.n1776 585
R4605 gnd.n4058 gnd.n1776 585
R4606 gnd.n4063 gnd.n4062 585
R4607 gnd.n4062 gnd.n4061 585
R4608 gnd.n1780 gnd.n1779 585
R4609 gnd.n4049 gnd.n1780 585
R4610 gnd.n3880 gnd.n3879 585
R4611 gnd.n3879 gnd.n3878 585
R4612 gnd.n3881 gnd.n1972 585
R4613 gnd.n1972 gnd.n1964 585
R4614 gnd.n3883 gnd.n3882 585
R4615 gnd.n3884 gnd.n3883 585
R4616 gnd.n1973 gnd.n1971 585
R4617 gnd.n1990 gnd.n1971 585
R4618 gnd.n3872 gnd.n3871 585
R4619 gnd.n3871 gnd.n3870 585
R4620 gnd.n1976 gnd.n1975 585
R4621 gnd.n1983 gnd.n1976 585
R4622 gnd.n3832 gnd.n3831 585
R4623 gnd.n3833 gnd.n3832 585
R4624 gnd.n1995 gnd.n1994 585
R4625 gnd.n2002 gnd.n1994 585
R4626 gnd.n3827 gnd.n3826 585
R4627 gnd.n3826 gnd.n3825 585
R4628 gnd.n1998 gnd.n1997 585
R4629 gnd.n2007 gnd.n1998 585
R4630 gnd.n3791 gnd.n3790 585
R4631 gnd.n3792 gnd.n3791 585
R4632 gnd.n2017 gnd.n2016 585
R4633 gnd.n2035 gnd.n2016 585
R4634 gnd.n3786 gnd.n3785 585
R4635 gnd.n3785 gnd.n3784 585
R4636 gnd.n2020 gnd.n2019 585
R4637 gnd.n2028 gnd.n2020 585
R4638 gnd.n3752 gnd.n3751 585
R4639 gnd.n3753 gnd.n3752 585
R4640 gnd.n2040 gnd.n2039 585
R4641 gnd.n2058 gnd.n2039 585
R4642 gnd.n3747 gnd.n3746 585
R4643 gnd.n3746 gnd.n3745 585
R4644 gnd.n2043 gnd.n2042 585
R4645 gnd.n2051 gnd.n2043 585
R4646 gnd.n3712 gnd.n3711 585
R4647 gnd.n3713 gnd.n3712 585
R4648 gnd.n2063 gnd.n2062 585
R4649 gnd.n3686 gnd.n2062 585
R4650 gnd.n3707 gnd.n3706 585
R4651 gnd.n3706 gnd.n3705 585
R4652 gnd.n2066 gnd.n2065 585
R4653 gnd.n3694 gnd.n2066 585
R4654 gnd.n3662 gnd.n2092 585
R4655 gnd.n2092 gnd.n2084 585
R4656 gnd.n3664 gnd.n3663 585
R4657 gnd.n3665 gnd.n3664 585
R4658 gnd.n2093 gnd.n2091 585
R4659 gnd.n2091 gnd.n2088 585
R4660 gnd.n3657 gnd.n3656 585
R4661 gnd.n3656 gnd.n3655 585
R4662 gnd.n2096 gnd.n2095 585
R4663 gnd.n2102 gnd.n2096 585
R4664 gnd.n3632 gnd.n3631 585
R4665 gnd.n3633 gnd.n3632 585
R4666 gnd.n2114 gnd.n2113 585
R4667 gnd.n3374 gnd.n2113 585
R4668 gnd.n3627 gnd.n3626 585
R4669 gnd.n3626 gnd.n3625 585
R4670 gnd.n2117 gnd.n2116 585
R4671 gnd.n2124 gnd.n2117 585
R4672 gnd.n3581 gnd.n2142 585
R4673 gnd.n2142 gnd.n2135 585
R4674 gnd.n3583 gnd.n3582 585
R4675 gnd.n3584 gnd.n3583 585
R4676 gnd.n2143 gnd.n2141 585
R4677 gnd.n2141 gnd.n2139 585
R4678 gnd.n3576 gnd.n3575 585
R4679 gnd.n3575 gnd.n3574 585
R4680 gnd.n2146 gnd.n2145 585
R4681 gnd.n3566 gnd.n2146 585
R4682 gnd.n3553 gnd.n3552 585
R4683 gnd.n3554 gnd.n3553 585
R4684 gnd.n2166 gnd.n2165 585
R4685 gnd.n2172 gnd.n2165 585
R4686 gnd.n3548 gnd.n3547 585
R4687 gnd.n3547 gnd.n3546 585
R4688 gnd.n2169 gnd.n2168 585
R4689 gnd.n2177 gnd.n2169 585
R4690 gnd.n3516 gnd.n2194 585
R4691 gnd.n2194 gnd.n2186 585
R4692 gnd.n3518 gnd.n3517 585
R4693 gnd.n3519 gnd.n3518 585
R4694 gnd.n2195 gnd.n2193 585
R4695 gnd.n3411 gnd.n2193 585
R4696 gnd.n3511 gnd.n3510 585
R4697 gnd.n3510 gnd.n3509 585
R4698 gnd.n2198 gnd.n2197 585
R4699 gnd.n3501 gnd.n2198 585
R4700 gnd.n3488 gnd.n3487 585
R4701 gnd.n3489 gnd.n3488 585
R4702 gnd.n2217 gnd.n2216 585
R4703 gnd.n3421 gnd.n2216 585
R4704 gnd.n3483 gnd.n3482 585
R4705 gnd.n3482 gnd.n3481 585
R4706 gnd.n2220 gnd.n2219 585
R4707 gnd.n3470 gnd.n2220 585
R4708 gnd.n3457 gnd.n3456 585
R4709 gnd.n3458 gnd.n3457 585
R4710 gnd.n2238 gnd.n2237 585
R4711 gnd.n3431 gnd.n2237 585
R4712 gnd.n3452 gnd.n3451 585
R4713 gnd.n3451 gnd.n3450 585
R4714 gnd.n2241 gnd.n2240 585
R4715 gnd.n3439 gnd.n2241 585
R4716 gnd.n3366 gnd.n3365 585
R4717 gnd.n3367 gnd.n3366 585
R4718 gnd.n2256 gnd.n2255 585
R4719 gnd.n2263 gnd.n2255 585
R4720 gnd.n3361 gnd.n3360 585
R4721 gnd.n3360 gnd.n3359 585
R4722 gnd.n2259 gnd.n2258 585
R4723 gnd.n2322 gnd.n2259 585
R4724 gnd.n3177 gnd.n3176 585
R4725 gnd.n3178 gnd.n3177 585
R4726 gnd.n2533 gnd.n2532 585
R4727 gnd.n3168 gnd.n2532 585
R4728 gnd.n3172 gnd.n3171 585
R4729 gnd.n3171 gnd.n3170 585
R4730 gnd.n2536 gnd.n2535 585
R4731 gnd.n3166 gnd.n2536 585
R4732 gnd.n3163 gnd.n3162 585
R4733 gnd.n3164 gnd.n3163 585
R4734 gnd.n2541 gnd.n2540 585
R4735 gnd.n3154 gnd.n2540 585
R4736 gnd.n3158 gnd.n3157 585
R4737 gnd.n3157 gnd.n3156 585
R4738 gnd.n2544 gnd.n2543 585
R4739 gnd.n3152 gnd.n2544 585
R4740 gnd.n3149 gnd.n3148 585
R4741 gnd.n3150 gnd.n3149 585
R4742 gnd.n2549 gnd.n2548 585
R4743 gnd.n3140 gnd.n2548 585
R4744 gnd.n3144 gnd.n3143 585
R4745 gnd.n3143 gnd.n3142 585
R4746 gnd.n2552 gnd.n2551 585
R4747 gnd.n3138 gnd.n2552 585
R4748 gnd.n3135 gnd.n3134 585
R4749 gnd.n3136 gnd.n3135 585
R4750 gnd.n2555 gnd.n2554 585
R4751 gnd.n2554 gnd.n2553 585
R4752 gnd.n3130 gnd.n3129 585
R4753 gnd.n3129 gnd.n3128 585
R4754 gnd.n2558 gnd.n2557 585
R4755 gnd.n2994 gnd.n2558 585
R4756 gnd.n2992 gnd.n2991 585
R4757 gnd.n2993 gnd.n2992 585
R4758 gnd.n2561 gnd.n2560 585
R4759 gnd.n2560 gnd.n2559 585
R4760 gnd.n2987 gnd.n2986 585
R4761 gnd.n2986 gnd.n1329 585
R4762 gnd.n2985 gnd.n2563 585
R4763 gnd.n2985 gnd.n1326 585
R4764 gnd.n2984 gnd.n2983 585
R4765 gnd.n2984 gnd.n1319 585
R4766 gnd.n2565 gnd.n2564 585
R4767 gnd.n2564 gnd.n1316 585
R4768 gnd.n2979 gnd.n2978 585
R4769 gnd.n2978 gnd.n1308 585
R4770 gnd.n2977 gnd.n2567 585
R4771 gnd.n2977 gnd.n1305 585
R4772 gnd.n2976 gnd.n2975 585
R4773 gnd.n2976 gnd.n1297 585
R4774 gnd.n2569 gnd.n2568 585
R4775 gnd.n2929 gnd.n2568 585
R4776 gnd.n2971 gnd.n2970 585
R4777 gnd.n2970 gnd.n1287 585
R4778 gnd.n2969 gnd.n2571 585
R4779 gnd.n2969 gnd.n1284 585
R4780 gnd.n2968 gnd.n2967 585
R4781 gnd.n2968 gnd.n1276 585
R4782 gnd.n2573 gnd.n2572 585
R4783 gnd.n2572 gnd.n1273 585
R4784 gnd.n2963 gnd.n2962 585
R4785 gnd.n2962 gnd.n2961 585
R4786 gnd.n2576 gnd.n2575 585
R4787 gnd.n2576 gnd.n1263 585
R4788 gnd.n2903 gnd.n2599 585
R4789 gnd.n2599 gnd.n1255 585
R4790 gnd.n2905 gnd.n2904 585
R4791 gnd.n2906 gnd.n2905 585
R4792 gnd.n2600 gnd.n2598 585
R4793 gnd.n2598 gnd.n1245 585
R4794 gnd.n2624 gnd.n2623 585
R4795 gnd.n2624 gnd.n1242 585
R4796 gnd.n2626 gnd.n2625 585
R4797 gnd.n2625 gnd.n1237 585
R4798 gnd.n2628 gnd.n2627 585
R4799 gnd.n2628 gnd.n1234 585
R4800 gnd.n2879 gnd.n2878 585
R4801 gnd.n2878 gnd.n2877 585
R4802 gnd.n2881 gnd.n2880 585
R4803 gnd.n2881 gnd.n1225 585
R4804 gnd.n2883 gnd.n2882 585
R4805 gnd.n2882 gnd.n1220 585
R4806 gnd.n2885 gnd.n2884 585
R4807 gnd.n2886 gnd.n2885 585
R4808 gnd.n2622 gnd.n2621 585
R4809 gnd.n2622 gnd.n1207 585
R4810 gnd.n2620 gnd.n2610 585
R4811 gnd.n2610 gnd.n1204 585
R4812 gnd.n2895 gnd.n2608 585
R4813 gnd.n2895 gnd.n2894 585
R4814 gnd.n2897 gnd.n2896 585
R4815 gnd.n2896 gnd.n1196 585
R4816 gnd.n2609 gnd.n2607 585
R4817 gnd.n2836 gnd.n2609 585
R4818 gnd.n2787 gnd.n2786 585
R4819 gnd.n2787 gnd.n1186 585
R4820 gnd.n2789 gnd.n2788 585
R4821 gnd.n2788 gnd.n1183 585
R4822 gnd.n2790 gnd.n2780 585
R4823 gnd.n2780 gnd.n1175 585
R4824 gnd.n2792 gnd.n2791 585
R4825 gnd.n2792 gnd.n1172 585
R4826 gnd.n2793 gnd.n2779 585
R4827 gnd.n2793 gnd.n2648 585
R4828 gnd.n2795 gnd.n2794 585
R4829 gnd.n2794 gnd.n1162 585
R4830 gnd.n2796 gnd.n2657 585
R4831 gnd.n2657 gnd.n1154 585
R4832 gnd.n2798 gnd.n2797 585
R4833 gnd.n2799 gnd.n2798 585
R4834 gnd.n2658 gnd.n2656 585
R4835 gnd.n2656 gnd.n1145 585
R4836 gnd.n2773 gnd.n2772 585
R4837 gnd.n2772 gnd.n1142 585
R4838 gnd.n2771 gnd.n2660 585
R4839 gnd.n2771 gnd.n1133 585
R4840 gnd.n2770 gnd.n2769 585
R4841 gnd.n2770 gnd.n1130 585
R4842 gnd.n2756 gnd.n2755 585
R4843 gnd.n2755 gnd.n2754 585
R4844 gnd.n2765 gnd.n2764 585
R4845 gnd.n2764 gnd.n1121 585
R4846 gnd.n2763 gnd.n2758 585
R4847 gnd.n2763 gnd.n1119 585
R4848 gnd.n2762 gnd.n2761 585
R4849 gnd.n2762 gnd.n1069 585
R4850 gnd.n1040 gnd.n1039 585
R4851 gnd.n4716 gnd.n1040 585
R4852 gnd.n4719 gnd.n4718 585
R4853 gnd.n4718 gnd.n4717 585
R4854 gnd.n4720 gnd.n1034 585
R4855 gnd.n1034 gnd.n1033 585
R4856 gnd.n4722 gnd.n4721 585
R4857 gnd.n4723 gnd.n4722 585
R4858 gnd.n1032 gnd.n1031 585
R4859 gnd.n4724 gnd.n1032 585
R4860 gnd.n4727 gnd.n4726 585
R4861 gnd.n4726 gnd.n4725 585
R4862 gnd.n4728 gnd.n1026 585
R4863 gnd.n1026 gnd.n1025 585
R4864 gnd.n4730 gnd.n4729 585
R4865 gnd.n4731 gnd.n4730 585
R4866 gnd.n1024 gnd.n1023 585
R4867 gnd.n4732 gnd.n1024 585
R4868 gnd.n4735 gnd.n4734 585
R4869 gnd.n4734 gnd.n4733 585
R4870 gnd.n4736 gnd.n1018 585
R4871 gnd.n1018 gnd.n1017 585
R4872 gnd.n4738 gnd.n4737 585
R4873 gnd.n4739 gnd.n4738 585
R4874 gnd.n4379 gnd.n4378 585
R4875 gnd.n4378 gnd.n4377 585
R4876 gnd.n4380 gnd.n1436 585
R4877 gnd.n4115 gnd.n1436 585
R4878 gnd.n4381 gnd.n1435 585
R4879 gnd.n4101 gnd.n1435 585
R4880 gnd.n4103 gnd.n1433 585
R4881 gnd.n4104 gnd.n4103 585
R4882 gnd.n4385 gnd.n1432 585
R4883 gnd.n1757 gnd.n1432 585
R4884 gnd.n4386 gnd.n1431 585
R4885 gnd.n4092 gnd.n1431 585
R4886 gnd.n4387 gnd.n1430 585
R4887 gnd.n1763 gnd.n1430 585
R4888 gnd.n4080 gnd.n1428 585
R4889 gnd.n4081 gnd.n4080 585
R4890 gnd.n4391 gnd.n1427 585
R4891 gnd.n1769 gnd.n1427 585
R4892 gnd.n4392 gnd.n1426 585
R4893 gnd.n4071 gnd.n1426 585
R4894 gnd.n4393 gnd.n1425 585
R4895 gnd.n1775 gnd.n1425 585
R4896 gnd.n4059 gnd.n1423 585
R4897 gnd.n4060 gnd.n4059 585
R4898 gnd.n4397 gnd.n1422 585
R4899 gnd.n1804 gnd.n1422 585
R4900 gnd.n4398 gnd.n1421 585
R4901 gnd.n4050 gnd.n1421 585
R4902 gnd.n4399 gnd.n1420 585
R4903 gnd.n1965 gnd.n1420 585
R4904 gnd.n3851 gnd.n1418 585
R4905 gnd.n3852 gnd.n3851 585
R4906 gnd.n4403 gnd.n1417 585
R4907 gnd.n3848 gnd.n1417 585
R4908 gnd.n4404 gnd.n1416 585
R4909 gnd.n3869 gnd.n1416 585
R4910 gnd.n4405 gnd.n1415 585
R4911 gnd.n3861 gnd.n1415 585
R4912 gnd.n3834 gnd.n1413 585
R4913 gnd.n3835 gnd.n3834 585
R4914 gnd.n4409 gnd.n1412 585
R4915 gnd.n3805 gnd.n1412 585
R4916 gnd.n4410 gnd.n1411 585
R4917 gnd.n3824 gnd.n1411 585
R4918 gnd.n4411 gnd.n1410 585
R4919 gnd.n3813 gnd.n1410 585
R4920 gnd.n3793 gnd.n1408 585
R4921 gnd.n3794 gnd.n3793 585
R4922 gnd.n4415 gnd.n1407 585
R4923 gnd.n3766 gnd.n1407 585
R4924 gnd.n4416 gnd.n1406 585
R4925 gnd.n2023 gnd.n1406 585
R4926 gnd.n4417 gnd.n1405 585
R4927 gnd.n3774 gnd.n1405 585
R4928 gnd.n3754 gnd.n1403 585
R4929 gnd.n3755 gnd.n3754 585
R4930 gnd.n4421 gnd.n1402 585
R4931 gnd.n3726 gnd.n1402 585
R4932 gnd.n4422 gnd.n1401 585
R4933 gnd.n2046 gnd.n1401 585
R4934 gnd.n4423 gnd.n1400 585
R4935 gnd.n3734 gnd.n1400 585
R4936 gnd.n3714 gnd.n1398 585
R4937 gnd.n3715 gnd.n3714 585
R4938 gnd.n4427 gnd.n1397 585
R4939 gnd.n3685 gnd.n1397 585
R4940 gnd.n4428 gnd.n1396 585
R4941 gnd.n2068 gnd.n1396 585
R4942 gnd.n4429 gnd.n1395 585
R4943 gnd.n3693 gnd.n1395 585
R4944 gnd.n2073 gnd.n1393 585
R4945 gnd.n2074 gnd.n2073 585
R4946 gnd.n4433 gnd.n1392 585
R4947 gnd.n3675 gnd.n1392 585
R4948 gnd.n4434 gnd.n1391 585
R4949 gnd.n3667 gnd.n1391 585
R4950 gnd.n4435 gnd.n1390 585
R4951 gnd.n3654 gnd.n1390 585
R4952 gnd.n2103 gnd.n1388 585
R4953 gnd.n2104 gnd.n2103 585
R4954 gnd.n4439 gnd.n1387 585
R4955 gnd.n2112 gnd.n1387 585
R4956 gnd.n4440 gnd.n1386 585
R4957 gnd.n2109 gnd.n1386 585
R4958 gnd.n4441 gnd.n1385 585
R4959 gnd.n2120 gnd.n1385 585
R4960 gnd.n3616 gnd.n1383 585
R4961 gnd.n3617 gnd.n3616 585
R4962 gnd.n4445 gnd.n1382 585
R4963 gnd.n3382 gnd.n1382 585
R4964 gnd.n4446 gnd.n1381 585
R4965 gnd.n3593 gnd.n1381 585
R4966 gnd.n4447 gnd.n1380 585
R4967 gnd.n3585 gnd.n1380 585
R4968 gnd.n2148 gnd.n1378 585
R4969 gnd.n2149 gnd.n2148 585
R4970 gnd.n4451 gnd.n1377 585
R4971 gnd.n3564 gnd.n1377 585
R4972 gnd.n4452 gnd.n1376 585
R4973 gnd.n2153 gnd.n1376 585
R4974 gnd.n4453 gnd.n1375 585
R4975 gnd.n3555 gnd.n1375 585
R4976 gnd.n3544 gnd.n1373 585
R4977 gnd.n3545 gnd.n3544 585
R4978 gnd.n4457 gnd.n1372 585
R4979 gnd.n3535 gnd.n1372 585
R4980 gnd.n4458 gnd.n1371 585
R4981 gnd.n3403 gnd.n1371 585
R4982 gnd.n4459 gnd.n1370 585
R4983 gnd.n3527 gnd.n1370 585
R4984 gnd.n2190 gnd.n1368 585
R4985 gnd.n2191 gnd.n2190 585
R4986 gnd.n4463 gnd.n1367 585
R4987 gnd.n2201 gnd.n1367 585
R4988 gnd.n4464 gnd.n1366 585
R4989 gnd.n3500 gnd.n1366 585
R4990 gnd.n4465 gnd.n1365 585
R4991 gnd.n2205 gnd.n1365 585
R4992 gnd.n3490 gnd.n1363 585
R4993 gnd.n3491 gnd.n3490 585
R4994 gnd.n4469 gnd.n1362 585
R4995 gnd.n2222 gnd.n1362 585
R4996 gnd.n4470 gnd.n1361 585
R4997 gnd.n3468 gnd.n1361 585
R4998 gnd.n4471 gnd.n1360 585
R4999 gnd.n2235 gnd.n1360 585
R5000 gnd.n3459 gnd.n1358 585
R5001 gnd.n3460 gnd.n3459 585
R5002 gnd.n4475 gnd.n1357 585
R5003 gnd.n2244 gnd.n1357 585
R5004 gnd.n4476 gnd.n1356 585
R5005 gnd.n2242 gnd.n1356 585
R5006 gnd.n4477 gnd.n1355 585
R5007 gnd.n2249 gnd.n1355 585
R5008 gnd.n2253 gnd.n1353 585
R5009 gnd.n2254 gnd.n2253 585
R5010 gnd.n4481 gnd.n1352 585
R5011 gnd.n3358 gnd.n1352 585
R5012 gnd.n4482 gnd.n1351 585
R5013 gnd.n3183 gnd.n1351 585
R5014 gnd.n4483 gnd.n1350 585
R5015 gnd.n2289 gnd.n1350 585
R5016 gnd.n3179 gnd.n1348 585
R5017 gnd.n3180 gnd.n3179 585
R5018 gnd.n4487 gnd.n1347 585
R5019 gnd.n3169 gnd.n1347 585
R5020 gnd.n4488 gnd.n1346 585
R5021 gnd.n3167 gnd.n1346 585
R5022 gnd.n4489 gnd.n1345 585
R5023 gnd.n3165 gnd.n1345 585
R5024 gnd.n2538 gnd.n1343 585
R5025 gnd.n2539 gnd.n2538 585
R5026 gnd.n4493 gnd.n1342 585
R5027 gnd.n3155 gnd.n1342 585
R5028 gnd.n4494 gnd.n1341 585
R5029 gnd.n3153 gnd.n1341 585
R5030 gnd.n4495 gnd.n1340 585
R5031 gnd.n3151 gnd.n1340 585
R5032 gnd.n2546 gnd.n1338 585
R5033 gnd.n2547 gnd.n2546 585
R5034 gnd.n4499 gnd.n1337 585
R5035 gnd.n3141 gnd.n1337 585
R5036 gnd.n4500 gnd.n1336 585
R5037 gnd.n3139 gnd.n1336 585
R5038 gnd.n4501 gnd.n1335 585
R5039 gnd.n3137 gnd.n1335 585
R5040 gnd.n3125 gnd.n3124 585
R5041 gnd.n3123 gnd.n3011 585
R5042 gnd.n3013 gnd.n3010 585
R5043 gnd.n3127 gnd.n3010 585
R5044 gnd.n3116 gnd.n3026 585
R5045 gnd.n3115 gnd.n3027 585
R5046 gnd.n3029 gnd.n3028 585
R5047 gnd.n3108 gnd.n3037 585
R5048 gnd.n3107 gnd.n3038 585
R5049 gnd.n3048 gnd.n3039 585
R5050 gnd.n3100 gnd.n3049 585
R5051 gnd.n3099 gnd.n3050 585
R5052 gnd.n3052 gnd.n3051 585
R5053 gnd.n3092 gnd.n3060 585
R5054 gnd.n3091 gnd.n3061 585
R5055 gnd.n3073 gnd.n3062 585
R5056 gnd.n3084 gnd.n3074 585
R5057 gnd.n3083 gnd.n3076 585
R5058 gnd.n3075 gnd.n2499 585
R5059 gnd.n3232 gnd.n2500 585
R5060 gnd.n3231 gnd.n2501 585
R5061 gnd.n3230 gnd.n2502 585
R5062 gnd.n3004 gnd.n2503 585
R5063 gnd.n3226 gnd.n2505 585
R5064 gnd.n3225 gnd.n2506 585
R5065 gnd.n3224 gnd.n2507 585
R5066 gnd.n3221 gnd.n2512 585
R5067 gnd.n3220 gnd.n2513 585
R5068 gnd.n3219 gnd.n2514 585
R5069 gnd.n3008 gnd.n2515 585
R5070 gnd.n4118 gnd.n1440 585
R5071 gnd.n4377 gnd.n1440 585
R5072 gnd.n4117 gnd.n4116 585
R5073 gnd.n4116 gnd.n4115 585
R5074 gnd.n1751 gnd.n1750 585
R5075 gnd.n4101 gnd.n1751 585
R5076 gnd.n4100 gnd.n4099 585
R5077 gnd.n4104 gnd.n4100 585
R5078 gnd.n1759 gnd.n1758 585
R5079 gnd.n1758 gnd.n1757 585
R5080 gnd.n4094 gnd.n4093 585
R5081 gnd.n4093 gnd.n4092 585
R5082 gnd.n1762 gnd.n1761 585
R5083 gnd.n1763 gnd.n1762 585
R5084 gnd.n4078 gnd.n4077 585
R5085 gnd.n4081 gnd.n4078 585
R5086 gnd.n1771 gnd.n1770 585
R5087 gnd.n1770 gnd.n1769 585
R5088 gnd.n4073 gnd.n4072 585
R5089 gnd.n4072 gnd.n4071 585
R5090 gnd.n1774 gnd.n1773 585
R5091 gnd.n1775 gnd.n1774 585
R5092 gnd.n4057 gnd.n4056 585
R5093 gnd.n4060 gnd.n4057 585
R5094 gnd.n1782 gnd.n1781 585
R5095 gnd.n1804 gnd.n1781 585
R5096 gnd.n4052 gnd.n4051 585
R5097 gnd.n4051 gnd.n4050 585
R5098 gnd.n1785 gnd.n1784 585
R5099 gnd.n1965 gnd.n1785 585
R5100 gnd.n3854 gnd.n3853 585
R5101 gnd.n3853 gnd.n3852 585
R5102 gnd.n3855 gnd.n3849 585
R5103 gnd.n3849 gnd.n3848 585
R5104 gnd.n1987 gnd.n1978 585
R5105 gnd.n3869 gnd.n1978 585
R5106 gnd.n3860 gnd.n3859 585
R5107 gnd.n3861 gnd.n3860 585
R5108 gnd.n1986 gnd.n1985 585
R5109 gnd.n3835 gnd.n1985 585
R5110 gnd.n3807 gnd.n3806 585
R5111 gnd.n3806 gnd.n3805 585
R5112 gnd.n2011 gnd.n2000 585
R5113 gnd.n3824 gnd.n2000 585
R5114 gnd.n3812 gnd.n3811 585
R5115 gnd.n3813 gnd.n3812 585
R5116 gnd.n2010 gnd.n2009 585
R5117 gnd.n3794 gnd.n2009 585
R5118 gnd.n3768 gnd.n3767 585
R5119 gnd.n3767 gnd.n3766 585
R5120 gnd.n2033 gnd.n2031 585
R5121 gnd.n2031 gnd.n2023 585
R5122 gnd.n3773 gnd.n3772 585
R5123 gnd.n3774 gnd.n3773 585
R5124 gnd.n2032 gnd.n2030 585
R5125 gnd.n3755 gnd.n2030 585
R5126 gnd.n3728 gnd.n3727 585
R5127 gnd.n3727 gnd.n3726 585
R5128 gnd.n2056 gnd.n2054 585
R5129 gnd.n2054 gnd.n2046 585
R5130 gnd.n3733 gnd.n3732 585
R5131 gnd.n3734 gnd.n3733 585
R5132 gnd.n2055 gnd.n2053 585
R5133 gnd.n3715 gnd.n2053 585
R5134 gnd.n3684 gnd.n3683 585
R5135 gnd.n3685 gnd.n3684 585
R5136 gnd.n2079 gnd.n2078 585
R5137 gnd.n2078 gnd.n2068 585
R5138 gnd.n3679 gnd.n2076 585
R5139 gnd.n3693 gnd.n2076 585
R5140 gnd.n3678 gnd.n3677 585
R5141 gnd.n3677 gnd.n2074 585
R5142 gnd.n3676 gnd.n2081 585
R5143 gnd.n3676 gnd.n3675 585
R5144 gnd.n3604 gnd.n2082 585
R5145 gnd.n3667 gnd.n2082 585
R5146 gnd.n3602 gnd.n2098 585
R5147 gnd.n3654 gnd.n2098 585
R5148 gnd.n3608 gnd.n3601 585
R5149 gnd.n3601 gnd.n2104 585
R5150 gnd.n3609 gnd.n3600 585
R5151 gnd.n3600 gnd.n2112 585
R5152 gnd.n3610 gnd.n3599 585
R5153 gnd.n3599 gnd.n2109 585
R5154 gnd.n2129 gnd.n2127 585
R5155 gnd.n2127 gnd.n2120 585
R5156 gnd.n3615 gnd.n3614 585
R5157 gnd.n3617 gnd.n3615 585
R5158 gnd.n2128 gnd.n2126 585
R5159 gnd.n3382 gnd.n2126 585
R5160 gnd.n3595 gnd.n3594 585
R5161 gnd.n3594 gnd.n3593 585
R5162 gnd.n2132 gnd.n2131 585
R5163 gnd.n3585 gnd.n2132 585
R5164 gnd.n2159 gnd.n2157 585
R5165 gnd.n2157 gnd.n2149 585
R5166 gnd.n3563 gnd.n3562 585
R5167 gnd.n3564 gnd.n3563 585
R5168 gnd.n2158 gnd.n2156 585
R5169 gnd.n2156 gnd.n2153 585
R5170 gnd.n3557 gnd.n3556 585
R5171 gnd.n3556 gnd.n3555 585
R5172 gnd.n2162 gnd.n2161 585
R5173 gnd.n3545 gnd.n2162 585
R5174 gnd.n3534 gnd.n3533 585
R5175 gnd.n3535 gnd.n3534 585
R5176 gnd.n2180 gnd.n2179 585
R5177 gnd.n3403 gnd.n2179 585
R5178 gnd.n3529 gnd.n3528 585
R5179 gnd.n3528 gnd.n3527 585
R5180 gnd.n2183 gnd.n2182 585
R5181 gnd.n2191 gnd.n2183 585
R5182 gnd.n2210 gnd.n2208 585
R5183 gnd.n2208 gnd.n2201 585
R5184 gnd.n3499 gnd.n3498 585
R5185 gnd.n3500 gnd.n3499 585
R5186 gnd.n2209 gnd.n2207 585
R5187 gnd.n2207 gnd.n2205 585
R5188 gnd.n3493 gnd.n3492 585
R5189 gnd.n3492 gnd.n3491 585
R5190 gnd.n2213 gnd.n2212 585
R5191 gnd.n2222 gnd.n2213 585
R5192 gnd.n3467 gnd.n3466 585
R5193 gnd.n3468 gnd.n3467 585
R5194 gnd.n2230 gnd.n2229 585
R5195 gnd.n2235 gnd.n2229 585
R5196 gnd.n3462 gnd.n3461 585
R5197 gnd.n3461 gnd.n3460 585
R5198 gnd.n2233 gnd.n2232 585
R5199 gnd.n2244 gnd.n2233 585
R5200 gnd.n3190 gnd.n3189 585
R5201 gnd.n3189 gnd.n2242 585
R5202 gnd.n3191 gnd.n3188 585
R5203 gnd.n3188 gnd.n2249 585
R5204 gnd.n3187 gnd.n3185 585
R5205 gnd.n3187 gnd.n2254 585
R5206 gnd.n3195 gnd.n2261 585
R5207 gnd.n3358 gnd.n2261 585
R5208 gnd.n3196 gnd.n3184 585
R5209 gnd.n3184 gnd.n3183 585
R5210 gnd.n3197 gnd.n3182 585
R5211 gnd.n3182 gnd.n2289 585
R5212 gnd.n3181 gnd.n2530 585
R5213 gnd.n3181 gnd.n3180 585
R5214 gnd.n3201 gnd.n2529 585
R5215 gnd.n3169 gnd.n2529 585
R5216 gnd.n3202 gnd.n2528 585
R5217 gnd.n3167 gnd.n2528 585
R5218 gnd.n3203 gnd.n2527 585
R5219 gnd.n3165 gnd.n2527 585
R5220 gnd.n2537 gnd.n2525 585
R5221 gnd.n2539 gnd.n2537 585
R5222 gnd.n3207 gnd.n2524 585
R5223 gnd.n3155 gnd.n2524 585
R5224 gnd.n3208 gnd.n2523 585
R5225 gnd.n3153 gnd.n2523 585
R5226 gnd.n3209 gnd.n2522 585
R5227 gnd.n3151 gnd.n2522 585
R5228 gnd.n2545 gnd.n2520 585
R5229 gnd.n2547 gnd.n2545 585
R5230 gnd.n3213 gnd.n2519 585
R5231 gnd.n3141 gnd.n2519 585
R5232 gnd.n3214 gnd.n2518 585
R5233 gnd.n3139 gnd.n2518 585
R5234 gnd.n3215 gnd.n2517 585
R5235 gnd.n3137 gnd.n2517 585
R5236 gnd.n4125 gnd.n4124 585
R5237 gnd.n4124 gnd.n1450 585
R5238 gnd.n4126 gnd.n4123 585
R5239 gnd.n4121 gnd.n1748 585
R5240 gnd.n4130 gnd.n1747 585
R5241 gnd.n4134 gnd.n1745 585
R5242 gnd.n4135 gnd.n1744 585
R5243 gnd.n1742 gnd.n1740 585
R5244 gnd.n4139 gnd.n1739 585
R5245 gnd.n4140 gnd.n1737 585
R5246 gnd.n4141 gnd.n1736 585
R5247 gnd.n1734 gnd.n1600 585
R5248 gnd.n1733 gnd.n1732 585
R5249 gnd.n1719 gnd.n1602 585
R5250 gnd.n1721 gnd.n1720 585
R5251 gnd.n1717 gnd.n1611 585
R5252 gnd.n1716 gnd.n1715 585
R5253 gnd.n1700 gnd.n1613 585
R5254 gnd.n1702 gnd.n1701 585
R5255 gnd.n1698 gnd.n1620 585
R5256 gnd.n1697 gnd.n1696 585
R5257 gnd.n1681 gnd.n1622 585
R5258 gnd.n1683 gnd.n1682 585
R5259 gnd.n1679 gnd.n1629 585
R5260 gnd.n1678 gnd.n1677 585
R5261 gnd.n1662 gnd.n1631 585
R5262 gnd.n1664 gnd.n1663 585
R5263 gnd.n1660 gnd.n1638 585
R5264 gnd.n1659 gnd.n1658 585
R5265 gnd.n1640 gnd.n1438 585
R5266 gnd.n6274 gnd.n6273 540.215
R5267 gnd.n3973 gnd.n1967 511.721
R5268 gnd.n3982 gnd.n3981 511.721
R5269 gnd.n2332 gnd.n2331 511.721
R5270 gnd.n3350 gnd.n2264 511.721
R5271 gnd.n2327 gnd.t106 389.64
R5272 gnd.n1959 gnd.t56 389.64
R5273 gnd.n2324 gnd.t27 389.64
R5274 gnd.n3907 gnd.t109 389.64
R5275 gnd.n2508 gnd.t96 371.625
R5276 gnd.n7211 gnd.t86 371.625
R5277 gnd.n1604 gnd.t70 371.625
R5278 gnd.n3069 gnd.t93 371.625
R5279 gnd.n1879 gnd.t67 371.625
R5280 gnd.n1908 gnd.t45 371.625
R5281 gnd.n157 gnd.t31 371.625
R5282 gnd.n7289 gnd.t60 371.625
R5283 gnd.n1091 gnd.t132 371.625
R5284 gnd.n1113 gnd.t119 371.625
R5285 gnd.n2673 gnd.t115 371.625
R5286 gnd.n2487 gnd.t63 371.625
R5287 gnd.n2398 gnd.t83 371.625
R5288 gnd.n4131 gnd.t73 371.625
R5289 gnd.n7005 gnd.n7004 368.44
R5290 gnd.n5138 gnd.t49 323.425
R5291 gnd.n4771 gnd.t89 323.425
R5292 gnd.n6795 gnd.n447 301.784
R5293 gnd.n6803 gnd.n447 301.784
R5294 gnd.n6804 gnd.n6803 301.784
R5295 gnd.n6805 gnd.n6804 301.784
R5296 gnd.n6805 gnd.n441 301.784
R5297 gnd.n6813 gnd.n441 301.784
R5298 gnd.n6814 gnd.n6813 301.784
R5299 gnd.n6815 gnd.n6814 301.784
R5300 gnd.n6815 gnd.n435 301.784
R5301 gnd.n6823 gnd.n435 301.784
R5302 gnd.n6824 gnd.n6823 301.784
R5303 gnd.n6825 gnd.n6824 301.784
R5304 gnd.n6825 gnd.n429 301.784
R5305 gnd.n6833 gnd.n429 301.784
R5306 gnd.n6834 gnd.n6833 301.784
R5307 gnd.n6835 gnd.n6834 301.784
R5308 gnd.n6835 gnd.n423 301.784
R5309 gnd.n6843 gnd.n423 301.784
R5310 gnd.n6844 gnd.n6843 301.784
R5311 gnd.n6845 gnd.n6844 301.784
R5312 gnd.n6845 gnd.n417 301.784
R5313 gnd.n6853 gnd.n417 301.784
R5314 gnd.n6854 gnd.n6853 301.784
R5315 gnd.n6855 gnd.n6854 301.784
R5316 gnd.n6855 gnd.n411 301.784
R5317 gnd.n6863 gnd.n411 301.784
R5318 gnd.n6864 gnd.n6863 301.784
R5319 gnd.n6865 gnd.n6864 301.784
R5320 gnd.n6865 gnd.n405 301.784
R5321 gnd.n6873 gnd.n405 301.784
R5322 gnd.n6874 gnd.n6873 301.784
R5323 gnd.n6875 gnd.n6874 301.784
R5324 gnd.n6875 gnd.n399 301.784
R5325 gnd.n6883 gnd.n399 301.784
R5326 gnd.n6884 gnd.n6883 301.784
R5327 gnd.n6885 gnd.n6884 301.784
R5328 gnd.n6885 gnd.n393 301.784
R5329 gnd.n6893 gnd.n393 301.784
R5330 gnd.n6894 gnd.n6893 301.784
R5331 gnd.n6895 gnd.n6894 301.784
R5332 gnd.n6895 gnd.n387 301.784
R5333 gnd.n6903 gnd.n387 301.784
R5334 gnd.n6904 gnd.n6903 301.784
R5335 gnd.n6905 gnd.n6904 301.784
R5336 gnd.n6905 gnd.n381 301.784
R5337 gnd.n6913 gnd.n381 301.784
R5338 gnd.n6914 gnd.n6913 301.784
R5339 gnd.n6915 gnd.n6914 301.784
R5340 gnd.n6915 gnd.n375 301.784
R5341 gnd.n6923 gnd.n375 301.784
R5342 gnd.n6924 gnd.n6923 301.784
R5343 gnd.n6925 gnd.n6924 301.784
R5344 gnd.n6925 gnd.n369 301.784
R5345 gnd.n6933 gnd.n369 301.784
R5346 gnd.n6934 gnd.n6933 301.784
R5347 gnd.n6935 gnd.n6934 301.784
R5348 gnd.n6935 gnd.n363 301.784
R5349 gnd.n6943 gnd.n363 301.784
R5350 gnd.n6944 gnd.n6943 301.784
R5351 gnd.n6945 gnd.n6944 301.784
R5352 gnd.n6945 gnd.n357 301.784
R5353 gnd.n6953 gnd.n357 301.784
R5354 gnd.n6954 gnd.n6953 301.784
R5355 gnd.n6955 gnd.n6954 301.784
R5356 gnd.n6955 gnd.n351 301.784
R5357 gnd.n6963 gnd.n351 301.784
R5358 gnd.n6964 gnd.n6963 301.784
R5359 gnd.n6965 gnd.n6964 301.784
R5360 gnd.n6965 gnd.n345 301.784
R5361 gnd.n6973 gnd.n345 301.784
R5362 gnd.n6974 gnd.n6973 301.784
R5363 gnd.n6975 gnd.n6974 301.784
R5364 gnd.n6975 gnd.n339 301.784
R5365 gnd.n6983 gnd.n339 301.784
R5366 gnd.n6984 gnd.n6983 301.784
R5367 gnd.n6985 gnd.n6984 301.784
R5368 gnd.n6985 gnd.n333 301.784
R5369 gnd.n6993 gnd.n333 301.784
R5370 gnd.n6994 gnd.n6993 301.784
R5371 gnd.n6995 gnd.n6994 301.784
R5372 gnd.n6995 gnd.n327 301.784
R5373 gnd.n7003 gnd.n327 301.784
R5374 gnd.n7004 gnd.n7003 301.784
R5375 gnd.n5916 gnd.n5890 289.615
R5376 gnd.n5884 gnd.n5858 289.615
R5377 gnd.n5852 gnd.n5826 289.615
R5378 gnd.n5821 gnd.n5795 289.615
R5379 gnd.n5789 gnd.n5763 289.615
R5380 gnd.n5757 gnd.n5731 289.615
R5381 gnd.n5725 gnd.n5699 289.615
R5382 gnd.n5694 gnd.n5668 289.615
R5383 gnd.n5212 gnd.t122 279.217
R5384 gnd.n4815 gnd.t35 279.217
R5385 gnd.n2273 gnd.t44 260.649
R5386 gnd.n3899 gnd.t79 260.649
R5387 gnd.n3349 gnd.n3348 256.663
R5388 gnd.n3348 gnd.n2290 256.663
R5389 gnd.n3348 gnd.n2291 256.663
R5390 gnd.n3348 gnd.n2292 256.663
R5391 gnd.n3348 gnd.n2293 256.663
R5392 gnd.n3348 gnd.n2294 256.663
R5393 gnd.n3348 gnd.n2295 256.663
R5394 gnd.n3348 gnd.n2296 256.663
R5395 gnd.n3348 gnd.n2297 256.663
R5396 gnd.n3348 gnd.n2298 256.663
R5397 gnd.n3348 gnd.n2299 256.663
R5398 gnd.n3348 gnd.n2300 256.663
R5399 gnd.n3348 gnd.n2301 256.663
R5400 gnd.n3348 gnd.n2302 256.663
R5401 gnd.n3348 gnd.n2303 256.663
R5402 gnd.n3348 gnd.n2304 256.663
R5403 gnd.n3288 gnd.n3285 256.663
R5404 gnd.n3348 gnd.n2305 256.663
R5405 gnd.n3348 gnd.n2306 256.663
R5406 gnd.n3348 gnd.n2307 256.663
R5407 gnd.n3348 gnd.n2308 256.663
R5408 gnd.n3348 gnd.n2309 256.663
R5409 gnd.n3348 gnd.n2310 256.663
R5410 gnd.n3348 gnd.n2311 256.663
R5411 gnd.n3348 gnd.n2312 256.663
R5412 gnd.n3348 gnd.n2313 256.663
R5413 gnd.n3348 gnd.n2314 256.663
R5414 gnd.n3348 gnd.n2315 256.663
R5415 gnd.n3348 gnd.n2316 256.663
R5416 gnd.n3348 gnd.n2317 256.663
R5417 gnd.n3348 gnd.n2318 256.663
R5418 gnd.n3348 gnd.n2319 256.663
R5419 gnd.n3348 gnd.n2320 256.663
R5420 gnd.n3348 gnd.n2321 256.663
R5421 gnd.n4048 gnd.n1805 256.663
R5422 gnd.n4048 gnd.n1806 256.663
R5423 gnd.n4048 gnd.n1807 256.663
R5424 gnd.n4048 gnd.n1808 256.663
R5425 gnd.n4048 gnd.n1809 256.663
R5426 gnd.n4048 gnd.n1810 256.663
R5427 gnd.n4048 gnd.n1811 256.663
R5428 gnd.n4048 gnd.n1812 256.663
R5429 gnd.n4048 gnd.n1813 256.663
R5430 gnd.n4048 gnd.n1814 256.663
R5431 gnd.n4048 gnd.n1815 256.663
R5432 gnd.n4048 gnd.n1816 256.663
R5433 gnd.n4048 gnd.n1817 256.663
R5434 gnd.n4048 gnd.n1818 256.663
R5435 gnd.n4048 gnd.n1819 256.663
R5436 gnd.n4048 gnd.n1820 256.663
R5437 gnd.n1958 gnd.n1821 256.663
R5438 gnd.n4048 gnd.n1803 256.663
R5439 gnd.n4048 gnd.n1802 256.663
R5440 gnd.n4048 gnd.n1801 256.663
R5441 gnd.n4048 gnd.n1800 256.663
R5442 gnd.n4048 gnd.n1799 256.663
R5443 gnd.n4048 gnd.n1798 256.663
R5444 gnd.n4048 gnd.n1797 256.663
R5445 gnd.n4048 gnd.n1796 256.663
R5446 gnd.n4048 gnd.n1795 256.663
R5447 gnd.n4048 gnd.n1794 256.663
R5448 gnd.n4048 gnd.n1793 256.663
R5449 gnd.n4048 gnd.n1792 256.663
R5450 gnd.n4048 gnd.n1791 256.663
R5451 gnd.n4048 gnd.n1790 256.663
R5452 gnd.n4048 gnd.n1789 256.663
R5453 gnd.n4048 gnd.n1788 256.663
R5454 gnd.n4048 gnd.n1787 256.663
R5455 gnd.n4715 gnd.n1059 242.672
R5456 gnd.n4715 gnd.n1060 242.672
R5457 gnd.n4715 gnd.n1061 242.672
R5458 gnd.n4715 gnd.n1062 242.672
R5459 gnd.n4715 gnd.n1063 242.672
R5460 gnd.n4715 gnd.n1064 242.672
R5461 gnd.n4715 gnd.n1065 242.672
R5462 gnd.n4715 gnd.n1066 242.672
R5463 gnd.n4715 gnd.n1067 242.672
R5464 gnd.n3078 gnd.n2459 242.672
R5465 gnd.n3067 gnd.n2459 242.672
R5466 gnd.n3064 gnd.n2459 242.672
R5467 gnd.n3055 gnd.n2459 242.672
R5468 gnd.n3044 gnd.n2459 242.672
R5469 gnd.n3041 gnd.n2459 242.672
R5470 gnd.n3032 gnd.n2459 242.672
R5471 gnd.n3022 gnd.n2459 242.672
R5472 gnd.n3019 gnd.n2459 242.672
R5473 gnd.n1650 gnd.n1451 242.672
R5474 gnd.n1652 gnd.n1451 242.672
R5475 gnd.n1669 gnd.n1451 242.672
R5476 gnd.n1671 gnd.n1451 242.672
R5477 gnd.n1688 gnd.n1451 242.672
R5478 gnd.n1690 gnd.n1451 242.672
R5479 gnd.n1707 gnd.n1451 242.672
R5480 gnd.n1709 gnd.n1451 242.672
R5481 gnd.n1726 gnd.n1451 242.672
R5482 gnd.n7213 gnd.n94 242.672
R5483 gnd.n7209 gnd.n94 242.672
R5484 gnd.n7204 gnd.n94 242.672
R5485 gnd.n7201 gnd.n94 242.672
R5486 gnd.n7196 gnd.n94 242.672
R5487 gnd.n7193 gnd.n94 242.672
R5488 gnd.n7188 gnd.n94 242.672
R5489 gnd.n7185 gnd.n94 242.672
R5490 gnd.n7180 gnd.n94 242.672
R5491 gnd.n5266 gnd.n5265 242.672
R5492 gnd.n5266 gnd.n5176 242.672
R5493 gnd.n5266 gnd.n5177 242.672
R5494 gnd.n5266 gnd.n5178 242.672
R5495 gnd.n5266 gnd.n5179 242.672
R5496 gnd.n5266 gnd.n5180 242.672
R5497 gnd.n5266 gnd.n5181 242.672
R5498 gnd.n5266 gnd.n5182 242.672
R5499 gnd.n5266 gnd.n5183 242.672
R5500 gnd.n5266 gnd.n5184 242.672
R5501 gnd.n5266 gnd.n5185 242.672
R5502 gnd.n5266 gnd.n5186 242.672
R5503 gnd.n5267 gnd.n5266 242.672
R5504 gnd.n5972 gnd.n4741 242.672
R5505 gnd.n5978 gnd.n4741 242.672
R5506 gnd.n4818 gnd.n4741 242.672
R5507 gnd.n5985 gnd.n4741 242.672
R5508 gnd.n4809 gnd.n4741 242.672
R5509 gnd.n5992 gnd.n4741 242.672
R5510 gnd.n4802 gnd.n4741 242.672
R5511 gnd.n5999 gnd.n4741 242.672
R5512 gnd.n4795 gnd.n4741 242.672
R5513 gnd.n6006 gnd.n4741 242.672
R5514 gnd.n4788 gnd.n4741 242.672
R5515 gnd.n6013 gnd.n4741 242.672
R5516 gnd.n4781 gnd.n4741 242.672
R5517 gnd.n5350 gnd.n5349 242.672
R5518 gnd.n5349 gnd.n5088 242.672
R5519 gnd.n5349 gnd.n5089 242.672
R5520 gnd.n5349 gnd.n5090 242.672
R5521 gnd.n5349 gnd.n5091 242.672
R5522 gnd.n5349 gnd.n5092 242.672
R5523 gnd.n5349 gnd.n5093 242.672
R5524 gnd.n5349 gnd.n5094 242.672
R5525 gnd.n6024 gnd.n4741 242.672
R5526 gnd.n4774 gnd.n4741 242.672
R5527 gnd.n6031 gnd.n4741 242.672
R5528 gnd.n4765 gnd.n4741 242.672
R5529 gnd.n6038 gnd.n4741 242.672
R5530 gnd.n4758 gnd.n4741 242.672
R5531 gnd.n6045 gnd.n4741 242.672
R5532 gnd.n4751 gnd.n4741 242.672
R5533 gnd.n4715 gnd.n4714 242.672
R5534 gnd.n4715 gnd.n1041 242.672
R5535 gnd.n4715 gnd.n1042 242.672
R5536 gnd.n4715 gnd.n1043 242.672
R5537 gnd.n4715 gnd.n1044 242.672
R5538 gnd.n4715 gnd.n1045 242.672
R5539 gnd.n4715 gnd.n1046 242.672
R5540 gnd.n4715 gnd.n1047 242.672
R5541 gnd.n4715 gnd.n1048 242.672
R5542 gnd.n4715 gnd.n1049 242.672
R5543 gnd.n4715 gnd.n1050 242.672
R5544 gnd.n4715 gnd.n1051 242.672
R5545 gnd.n4715 gnd.n1052 242.672
R5546 gnd.n4715 gnd.n1053 242.672
R5547 gnd.n4715 gnd.n1054 242.672
R5548 gnd.n4715 gnd.n1055 242.672
R5549 gnd.n4715 gnd.n1056 242.672
R5550 gnd.n4715 gnd.n1057 242.672
R5551 gnd.n4715 gnd.n1058 242.672
R5552 gnd.n3247 gnd.n2459 242.672
R5553 gnd.n2490 gnd.n2459 242.672
R5554 gnd.n3254 gnd.n2459 242.672
R5555 gnd.n2481 gnd.n2459 242.672
R5556 gnd.n3261 gnd.n2459 242.672
R5557 gnd.n2474 gnd.n2459 242.672
R5558 gnd.n3268 gnd.n2459 242.672
R5559 gnd.n2467 gnd.n2459 242.672
R5560 gnd.n3275 gnd.n2459 242.672
R5561 gnd.n3278 gnd.n2459 242.672
R5562 gnd.n2459 gnd.n2405 242.672
R5563 gnd.n3284 gnd.n2400 242.672
R5564 gnd.n2459 gnd.n2406 242.672
R5565 gnd.n2459 gnd.n2407 242.672
R5566 gnd.n2459 gnd.n2408 242.672
R5567 gnd.n2459 gnd.n2409 242.672
R5568 gnd.n2459 gnd.n2410 242.672
R5569 gnd.n2459 gnd.n2411 242.672
R5570 gnd.n2459 gnd.n2412 242.672
R5571 gnd.n2459 gnd.n2458 242.672
R5572 gnd.n1841 gnd.n1451 242.672
R5573 gnd.n1849 gnd.n1451 242.672
R5574 gnd.n1851 gnd.n1451 242.672
R5575 gnd.n1859 gnd.n1451 242.672
R5576 gnd.n1861 gnd.n1451 242.672
R5577 gnd.n1870 gnd.n1451 242.672
R5578 gnd.n1873 gnd.n1451 242.672
R5579 gnd.n1826 gnd.n1451 242.672
R5580 gnd.n1957 gnd.n1823 242.672
R5581 gnd.n1954 gnd.n1451 242.672
R5582 gnd.n1952 gnd.n1451 242.672
R5583 gnd.n1946 gnd.n1451 242.672
R5584 gnd.n1944 gnd.n1451 242.672
R5585 gnd.n1938 gnd.n1451 242.672
R5586 gnd.n1936 gnd.n1451 242.672
R5587 gnd.n1930 gnd.n1451 242.672
R5588 gnd.n1928 gnd.n1451 242.672
R5589 gnd.n1922 gnd.n1451 242.672
R5590 gnd.n1920 gnd.n1451 242.672
R5591 gnd.n1912 gnd.n1451 242.672
R5592 gnd.n154 gnd.n94 242.672
R5593 gnd.n7257 gnd.n94 242.672
R5594 gnd.n150 gnd.n94 242.672
R5595 gnd.n7264 gnd.n94 242.672
R5596 gnd.n143 gnd.n94 242.672
R5597 gnd.n7271 gnd.n94 242.672
R5598 gnd.n136 gnd.n94 242.672
R5599 gnd.n7278 gnd.n94 242.672
R5600 gnd.n129 gnd.n94 242.672
R5601 gnd.n7285 gnd.n94 242.672
R5602 gnd.n122 gnd.n94 242.672
R5603 gnd.n7295 gnd.n94 242.672
R5604 gnd.n115 gnd.n94 242.672
R5605 gnd.n7302 gnd.n94 242.672
R5606 gnd.n108 gnd.n94 242.672
R5607 gnd.n7309 gnd.n94 242.672
R5608 gnd.n101 gnd.n94 242.672
R5609 gnd.n7316 gnd.n94 242.672
R5610 gnd.n94 gnd.n93 242.672
R5611 gnd.n3127 gnd.n3126 242.672
R5612 gnd.n3127 gnd.n2995 242.672
R5613 gnd.n3127 gnd.n2996 242.672
R5614 gnd.n3127 gnd.n2997 242.672
R5615 gnd.n3127 gnd.n2998 242.672
R5616 gnd.n3127 gnd.n2999 242.672
R5617 gnd.n3127 gnd.n3000 242.672
R5618 gnd.n3127 gnd.n3001 242.672
R5619 gnd.n3127 gnd.n3002 242.672
R5620 gnd.n3127 gnd.n3003 242.672
R5621 gnd.n3127 gnd.n3005 242.672
R5622 gnd.n3127 gnd.n3006 242.672
R5623 gnd.n3127 gnd.n3007 242.672
R5624 gnd.n3127 gnd.n3009 242.672
R5625 gnd.n4122 gnd.n1450 242.672
R5626 gnd.n1746 gnd.n1450 242.672
R5627 gnd.n1743 gnd.n1450 242.672
R5628 gnd.n1738 gnd.n1450 242.672
R5629 gnd.n1735 gnd.n1450 242.672
R5630 gnd.n1601 gnd.n1450 242.672
R5631 gnd.n1718 gnd.n1450 242.672
R5632 gnd.n1612 gnd.n1450 242.672
R5633 gnd.n1699 gnd.n1450 242.672
R5634 gnd.n1621 gnd.n1450 242.672
R5635 gnd.n1680 gnd.n1450 242.672
R5636 gnd.n1630 gnd.n1450 242.672
R5637 gnd.n1661 gnd.n1450 242.672
R5638 gnd.n1639 gnd.n1450 242.672
R5639 gnd.n90 gnd.n86 240.244
R5640 gnd.n7318 gnd.n7317 240.244
R5641 gnd.n7315 gnd.n95 240.244
R5642 gnd.n7311 gnd.n7310 240.244
R5643 gnd.n7308 gnd.n102 240.244
R5644 gnd.n7304 gnd.n7303 240.244
R5645 gnd.n7301 gnd.n109 240.244
R5646 gnd.n7297 gnd.n7296 240.244
R5647 gnd.n7294 gnd.n116 240.244
R5648 gnd.n7287 gnd.n7286 240.244
R5649 gnd.n7284 gnd.n123 240.244
R5650 gnd.n7280 gnd.n7279 240.244
R5651 gnd.n7277 gnd.n130 240.244
R5652 gnd.n7273 gnd.n7272 240.244
R5653 gnd.n7270 gnd.n137 240.244
R5654 gnd.n7266 gnd.n7265 240.244
R5655 gnd.n7263 gnd.n144 240.244
R5656 gnd.n7259 gnd.n7258 240.244
R5657 gnd.n7256 gnd.n151 240.244
R5658 gnd.n4149 gnd.n1460 240.244
R5659 gnd.n4149 gnd.n1472 240.244
R5660 gnd.n4174 gnd.n1472 240.244
R5661 gnd.n4174 gnd.n1593 240.244
R5662 gnd.n1593 gnd.n1587 240.244
R5663 gnd.n1587 gnd.n1565 240.244
R5664 gnd.n4168 gnd.n1565 240.244
R5665 gnd.n4168 gnd.n1556 240.244
R5666 gnd.n4165 gnd.n1556 240.244
R5667 gnd.n4165 gnd.n1548 240.244
R5668 gnd.n1548 gnd.n1540 240.244
R5669 gnd.n1540 gnd.n1528 240.244
R5670 gnd.n4261 gnd.n1528 240.244
R5671 gnd.n4261 gnd.n1529 240.244
R5672 gnd.n1529 gnd.n1503 240.244
R5673 gnd.n1503 gnd.n1497 240.244
R5674 gnd.n4269 gnd.n1497 240.244
R5675 gnd.n4269 gnd.n234 240.244
R5676 gnd.n4297 gnd.n234 240.244
R5677 gnd.n4297 gnd.n1512 240.244
R5678 gnd.n1517 gnd.n1512 240.244
R5679 gnd.n4292 gnd.n1517 240.244
R5680 gnd.n4292 gnd.n4291 240.244
R5681 gnd.n4291 gnd.n256 240.244
R5682 gnd.n256 gnd.n249 240.244
R5683 gnd.n4283 gnd.n249 240.244
R5684 gnd.n4283 gnd.n221 240.244
R5685 gnd.n7083 gnd.n221 240.244
R5686 gnd.n7083 gnd.n212 240.244
R5687 gnd.n7079 gnd.n212 240.244
R5688 gnd.n7079 gnd.n204 240.244
R5689 gnd.n7075 gnd.n204 240.244
R5690 gnd.n7075 gnd.n195 240.244
R5691 gnd.n7049 gnd.n195 240.244
R5692 gnd.n7049 gnd.n189 240.244
R5693 gnd.n7064 gnd.n189 240.244
R5694 gnd.n7064 gnd.n180 240.244
R5695 gnd.n7060 gnd.n180 240.244
R5696 gnd.n7060 gnd.n170 240.244
R5697 gnd.n170 gnd.n161 240.244
R5698 gnd.n7248 gnd.n161 240.244
R5699 gnd.n7248 gnd.n82 240.244
R5700 gnd.n1842 gnd.n1837 240.244
R5701 gnd.n1848 gnd.n1837 240.244
R5702 gnd.n1852 gnd.n1850 240.244
R5703 gnd.n1858 gnd.n1833 240.244
R5704 gnd.n1862 gnd.n1860 240.244
R5705 gnd.n1869 gnd.n1829 240.244
R5706 gnd.n1872 gnd.n1871 240.244
R5707 gnd.n1874 gnd.n1827 240.244
R5708 gnd.n1955 gnd.n1953 240.244
R5709 gnd.n1951 gnd.n1883 240.244
R5710 gnd.n1947 gnd.n1945 240.244
R5711 gnd.n1943 gnd.n1889 240.244
R5712 gnd.n1939 gnd.n1937 240.244
R5713 gnd.n1935 gnd.n1895 240.244
R5714 gnd.n1931 gnd.n1929 240.244
R5715 gnd.n1927 gnd.n1901 240.244
R5716 gnd.n1923 gnd.n1921 240.244
R5717 gnd.n1919 gnd.n1907 240.244
R5718 gnd.n4360 gnd.n1465 240.244
R5719 gnd.n4356 gnd.n1465 240.244
R5720 gnd.n4356 gnd.n1470 240.244
R5721 gnd.n1585 gnd.n1470 240.244
R5722 gnd.n1585 gnd.n1563 240.244
R5723 gnd.n4198 gnd.n1563 240.244
R5724 gnd.n4198 gnd.n1558 240.244
R5725 gnd.n4206 gnd.n1558 240.244
R5726 gnd.n4206 gnd.n1559 240.244
R5727 gnd.n1559 gnd.n1538 240.244
R5728 gnd.n4251 gnd.n1538 240.244
R5729 gnd.n4251 gnd.n1534 240.244
R5730 gnd.n4259 gnd.n1534 240.244
R5731 gnd.n4259 gnd.n1500 240.244
R5732 gnd.n4327 gnd.n1500 240.244
R5733 gnd.n4328 gnd.n4327 240.244
R5734 gnd.n4328 gnd.n231 240.244
R5735 gnd.n7114 gnd.n231 240.244
R5736 gnd.n7114 gnd.n232 240.244
R5737 gnd.n4313 gnd.n232 240.244
R5738 gnd.n4313 gnd.n4310 240.244
R5739 gnd.n4310 gnd.n1514 240.244
R5740 gnd.n1514 gnd.n252 240.244
R5741 gnd.n7095 gnd.n252 240.244
R5742 gnd.n7097 gnd.n7095 240.244
R5743 gnd.n7097 gnd.n222 240.244
R5744 gnd.n7121 gnd.n222 240.244
R5745 gnd.n7121 gnd.n210 240.244
R5746 gnd.n7131 gnd.n210 240.244
R5747 gnd.n7131 gnd.n206 240.244
R5748 gnd.n7137 gnd.n206 240.244
R5749 gnd.n7137 gnd.n194 240.244
R5750 gnd.n7147 gnd.n194 240.244
R5751 gnd.n7147 gnd.n190 240.244
R5752 gnd.n7153 gnd.n190 240.244
R5753 gnd.n7153 gnd.n178 240.244
R5754 gnd.n7163 gnd.n178 240.244
R5755 gnd.n7163 gnd.n172 240.244
R5756 gnd.n7171 gnd.n172 240.244
R5757 gnd.n7171 gnd.n174 240.244
R5758 gnd.n174 gnd.n85 240.244
R5759 gnd.n7325 gnd.n85 240.244
R5760 gnd.n2413 gnd.n1325 240.244
R5761 gnd.n2457 gnd.n2414 240.244
R5762 gnd.n2453 gnd.n2452 240.244
R5763 gnd.n2449 gnd.n2448 240.244
R5764 gnd.n2445 gnd.n2444 240.244
R5765 gnd.n2441 gnd.n2440 240.244
R5766 gnd.n2437 gnd.n2436 240.244
R5767 gnd.n2433 gnd.n2432 240.244
R5768 gnd.n3279 gnd.n2404 240.244
R5769 gnd.n3277 gnd.n3276 240.244
R5770 gnd.n3274 gnd.n2461 240.244
R5771 gnd.n3270 gnd.n3269 240.244
R5772 gnd.n3267 gnd.n2468 240.244
R5773 gnd.n3263 gnd.n3262 240.244
R5774 gnd.n3260 gnd.n2475 240.244
R5775 gnd.n3256 gnd.n3255 240.244
R5776 gnd.n3253 gnd.n2482 240.244
R5777 gnd.n3249 gnd.n3248 240.244
R5778 gnd.n4636 gnd.n1117 240.244
R5779 gnd.n2668 gnd.n1117 240.244
R5780 gnd.n2668 gnd.n1131 240.244
R5781 gnd.n2746 gnd.n1131 240.244
R5782 gnd.n2746 gnd.n1143 240.244
R5783 gnd.n2801 gnd.n1143 240.244
R5784 gnd.n2801 gnd.n1152 240.244
R5785 gnd.n2807 gnd.n1152 240.244
R5786 gnd.n2807 gnd.n1163 240.244
R5787 gnd.n2817 gnd.n1163 240.244
R5788 gnd.n2817 gnd.n1173 240.244
R5789 gnd.n2824 gnd.n1173 240.244
R5790 gnd.n2824 gnd.n1184 240.244
R5791 gnd.n2838 gnd.n1184 240.244
R5792 gnd.n2838 gnd.n1194 240.244
R5793 gnd.n2638 gnd.n1194 240.244
R5794 gnd.n2638 gnd.n2612 240.244
R5795 gnd.n2612 gnd.n1205 240.244
R5796 gnd.n2619 gnd.n1205 240.244
R5797 gnd.n2619 gnd.n1218 240.244
R5798 gnd.n2855 gnd.n1218 240.244
R5799 gnd.n2855 gnd.n1226 240.244
R5800 gnd.n2629 gnd.n1226 240.244
R5801 gnd.n2629 gnd.n1235 240.244
R5802 gnd.n2867 gnd.n1235 240.244
R5803 gnd.n2867 gnd.n1243 240.244
R5804 gnd.n2597 gnd.n1243 240.244
R5805 gnd.n2597 gnd.n1253 240.244
R5806 gnd.n2916 gnd.n1253 240.244
R5807 gnd.n2916 gnd.n1264 240.244
R5808 gnd.n2577 gnd.n1264 240.244
R5809 gnd.n2577 gnd.n1274 240.244
R5810 gnd.n2924 gnd.n1274 240.244
R5811 gnd.n2924 gnd.n1285 240.244
R5812 gnd.n2931 gnd.n1285 240.244
R5813 gnd.n2931 gnd.n1295 240.244
R5814 gnd.n2935 gnd.n1295 240.244
R5815 gnd.n2935 gnd.n1306 240.244
R5816 gnd.n2942 gnd.n1306 240.244
R5817 gnd.n2942 gnd.n1317 240.244
R5818 gnd.n3240 gnd.n1317 240.244
R5819 gnd.n3240 gnd.n1327 240.244
R5820 gnd.n1071 gnd.n1070 240.244
R5821 gnd.n4708 gnd.n1070 240.244
R5822 gnd.n4706 gnd.n4705 240.244
R5823 gnd.n4702 gnd.n4701 240.244
R5824 gnd.n4698 gnd.n4697 240.244
R5825 gnd.n4694 gnd.n4693 240.244
R5826 gnd.n4690 gnd.n4689 240.244
R5827 gnd.n4686 gnd.n4685 240.244
R5828 gnd.n4682 gnd.n4681 240.244
R5829 gnd.n4677 gnd.n4676 240.244
R5830 gnd.n4673 gnd.n4672 240.244
R5831 gnd.n4669 gnd.n4668 240.244
R5832 gnd.n4665 gnd.n4664 240.244
R5833 gnd.n4661 gnd.n4660 240.244
R5834 gnd.n4657 gnd.n4656 240.244
R5835 gnd.n4653 gnd.n4652 240.244
R5836 gnd.n4649 gnd.n4648 240.244
R5837 gnd.n4645 gnd.n4644 240.244
R5838 gnd.n1112 gnd.n1111 240.244
R5839 gnd.n2666 gnd.n1072 240.244
R5840 gnd.n2666 gnd.n1134 240.244
R5841 gnd.n4625 gnd.n1134 240.244
R5842 gnd.n4625 gnd.n1135 240.244
R5843 gnd.n4621 gnd.n1135 240.244
R5844 gnd.n4621 gnd.n1141 240.244
R5845 gnd.n4613 gnd.n1141 240.244
R5846 gnd.n4613 gnd.n1155 240.244
R5847 gnd.n4609 gnd.n1155 240.244
R5848 gnd.n4609 gnd.n1161 240.244
R5849 gnd.n4601 gnd.n1161 240.244
R5850 gnd.n4601 gnd.n1176 240.244
R5851 gnd.n4597 gnd.n1176 240.244
R5852 gnd.n4597 gnd.n1182 240.244
R5853 gnd.n4589 gnd.n1182 240.244
R5854 gnd.n4589 gnd.n1197 240.244
R5855 gnd.n1201 gnd.n1197 240.244
R5856 gnd.n4583 gnd.n1201 240.244
R5857 gnd.n4583 gnd.n1203 240.244
R5858 gnd.n4575 gnd.n1203 240.244
R5859 gnd.n4575 gnd.n1221 240.244
R5860 gnd.n4570 gnd.n1221 240.244
R5861 gnd.n4570 gnd.n1224 240.244
R5862 gnd.n4562 gnd.n1224 240.244
R5863 gnd.n4562 gnd.n1238 240.244
R5864 gnd.n4557 gnd.n1238 240.244
R5865 gnd.n4557 gnd.n1241 240.244
R5866 gnd.n4549 gnd.n1241 240.244
R5867 gnd.n4549 gnd.n1256 240.244
R5868 gnd.n4545 gnd.n1256 240.244
R5869 gnd.n4545 gnd.n1262 240.244
R5870 gnd.n4537 gnd.n1262 240.244
R5871 gnd.n4537 gnd.n1277 240.244
R5872 gnd.n4533 gnd.n1277 240.244
R5873 gnd.n4533 gnd.n1283 240.244
R5874 gnd.n4525 gnd.n1283 240.244
R5875 gnd.n4525 gnd.n1298 240.244
R5876 gnd.n4521 gnd.n1298 240.244
R5877 gnd.n4521 gnd.n1304 240.244
R5878 gnd.n4513 gnd.n1304 240.244
R5879 gnd.n4513 gnd.n1320 240.244
R5880 gnd.n4509 gnd.n1320 240.244
R5881 gnd.n4748 gnd.n4743 240.244
R5882 gnd.n6047 gnd.n6046 240.244
R5883 gnd.n6044 gnd.n4752 240.244
R5884 gnd.n6040 gnd.n6039 240.244
R5885 gnd.n6037 gnd.n4759 240.244
R5886 gnd.n6033 gnd.n6032 240.244
R5887 gnd.n6030 gnd.n4766 240.244
R5888 gnd.n6026 gnd.n6025 240.244
R5889 gnd.n5361 gnd.n5073 240.244
R5890 gnd.n5371 gnd.n5073 240.244
R5891 gnd.n5371 gnd.n5064 240.244
R5892 gnd.n5064 gnd.n5053 240.244
R5893 gnd.n5392 gnd.n5053 240.244
R5894 gnd.n5392 gnd.n5047 240.244
R5895 gnd.n5402 gnd.n5047 240.244
R5896 gnd.n5402 gnd.n5036 240.244
R5897 gnd.n5036 gnd.n5028 240.244
R5898 gnd.n5420 gnd.n5028 240.244
R5899 gnd.n5421 gnd.n5420 240.244
R5900 gnd.n5421 gnd.n5013 240.244
R5901 gnd.n5423 gnd.n5013 240.244
R5902 gnd.n5423 gnd.n4999 240.244
R5903 gnd.n5465 gnd.n4999 240.244
R5904 gnd.n5466 gnd.n5465 240.244
R5905 gnd.n5469 gnd.n5466 240.244
R5906 gnd.n5469 gnd.n4954 240.244
R5907 gnd.n4994 gnd.n4954 240.244
R5908 gnd.n4994 gnd.n4964 240.244
R5909 gnd.n5479 gnd.n4964 240.244
R5910 gnd.n5479 gnd.n4985 240.244
R5911 gnd.n5489 gnd.n4985 240.244
R5912 gnd.n5489 gnd.n4895 240.244
R5913 gnd.n5534 gnd.n4895 240.244
R5914 gnd.n5534 gnd.n4881 240.244
R5915 gnd.n5556 gnd.n4881 240.244
R5916 gnd.n5557 gnd.n5556 240.244
R5917 gnd.n5557 gnd.n4868 240.244
R5918 gnd.n4868 gnd.n4857 240.244
R5919 gnd.n5588 gnd.n4857 240.244
R5920 gnd.n5589 gnd.n5588 240.244
R5921 gnd.n5590 gnd.n5589 240.244
R5922 gnd.n5590 gnd.n4842 240.244
R5923 gnd.n4842 gnd.n4834 240.244
R5924 gnd.n5643 gnd.n4834 240.244
R5925 gnd.n5644 gnd.n5643 240.244
R5926 gnd.n5644 gnd.n943 240.244
R5927 gnd.n5621 gnd.n943 240.244
R5928 gnd.n5621 gnd.n953 240.244
R5929 gnd.n5656 gnd.n953 240.244
R5930 gnd.n5657 gnd.n5656 240.244
R5931 gnd.n5657 gnd.n966 240.244
R5932 gnd.n5946 gnd.n966 240.244
R5933 gnd.n5946 gnd.n978 240.244
R5934 gnd.n5942 gnd.n978 240.244
R5935 gnd.n5942 gnd.n5941 240.244
R5936 gnd.n5941 gnd.n991 240.244
R5937 gnd.n5937 gnd.n991 240.244
R5938 gnd.n5937 gnd.n1004 240.244
R5939 gnd.n5933 gnd.n1004 240.244
R5940 gnd.n5933 gnd.n5932 240.244
R5941 gnd.n5932 gnd.n1016 240.244
R5942 gnd.n5351 gnd.n5086 240.244
R5943 gnd.n5107 gnd.n5086 240.244
R5944 gnd.n5110 gnd.n5109 240.244
R5945 gnd.n5117 gnd.n5116 240.244
R5946 gnd.n5120 gnd.n5119 240.244
R5947 gnd.n5127 gnd.n5126 240.244
R5948 gnd.n5130 gnd.n5129 240.244
R5949 gnd.n5137 gnd.n5136 240.244
R5950 gnd.n5359 gnd.n5083 240.244
R5951 gnd.n5083 gnd.n5062 240.244
R5952 gnd.n5382 gnd.n5062 240.244
R5953 gnd.n5382 gnd.n5056 240.244
R5954 gnd.n5390 gnd.n5056 240.244
R5955 gnd.n5390 gnd.n5058 240.244
R5956 gnd.n5058 gnd.n5034 240.244
R5957 gnd.n5412 gnd.n5034 240.244
R5958 gnd.n5412 gnd.n5030 240.244
R5959 gnd.n5418 gnd.n5030 240.244
R5960 gnd.n5418 gnd.n5012 240.244
R5961 gnd.n5443 gnd.n5012 240.244
R5962 gnd.n5443 gnd.n5007 240.244
R5963 gnd.n5455 gnd.n5007 240.244
R5964 gnd.n5455 gnd.n5008 240.244
R5965 gnd.n5451 gnd.n5008 240.244
R5966 gnd.n5451 gnd.n4956 240.244
R5967 gnd.n5503 gnd.n4956 240.244
R5968 gnd.n5503 gnd.n4957 240.244
R5969 gnd.n5499 gnd.n4957 240.244
R5970 gnd.n5499 gnd.n4963 240.244
R5971 gnd.n4983 gnd.n4963 240.244
R5972 gnd.n4983 gnd.n4893 240.244
R5973 gnd.n5538 gnd.n4893 240.244
R5974 gnd.n5538 gnd.n4888 240.244
R5975 gnd.n5546 gnd.n4888 240.244
R5976 gnd.n5546 gnd.n4889 240.244
R5977 gnd.n4889 gnd.n4866 240.244
R5978 gnd.n5578 gnd.n4866 240.244
R5979 gnd.n5578 gnd.n4861 240.244
R5980 gnd.n5586 gnd.n4861 240.244
R5981 gnd.n5586 gnd.n4862 240.244
R5982 gnd.n4862 gnd.n4840 240.244
R5983 gnd.n5634 gnd.n4840 240.244
R5984 gnd.n5634 gnd.n4836 240.244
R5985 gnd.n5641 gnd.n4836 240.244
R5986 gnd.n5641 gnd.n944 240.244
R5987 gnd.n6096 gnd.n944 240.244
R5988 gnd.n6096 gnd.n945 240.244
R5989 gnd.n6092 gnd.n945 240.244
R5990 gnd.n6092 gnd.n951 240.244
R5991 gnd.n967 gnd.n951 240.244
R5992 gnd.n6082 gnd.n967 240.244
R5993 gnd.n6082 gnd.n968 240.244
R5994 gnd.n6078 gnd.n968 240.244
R5995 gnd.n6078 gnd.n976 240.244
R5996 gnd.n993 gnd.n976 240.244
R5997 gnd.n6068 gnd.n993 240.244
R5998 gnd.n6068 gnd.n994 240.244
R5999 gnd.n6064 gnd.n994 240.244
R6000 gnd.n6064 gnd.n1002 240.244
R6001 gnd.n4742 gnd.n1002 240.244
R6002 gnd.n6054 gnd.n4742 240.244
R6003 gnd.n4778 gnd.n1013 240.244
R6004 gnd.n6015 gnd.n6014 240.244
R6005 gnd.n6012 gnd.n4782 240.244
R6006 gnd.n6008 gnd.n6007 240.244
R6007 gnd.n6005 gnd.n4789 240.244
R6008 gnd.n6001 gnd.n6000 240.244
R6009 gnd.n5998 gnd.n4796 240.244
R6010 gnd.n5994 gnd.n5993 240.244
R6011 gnd.n5991 gnd.n4803 240.244
R6012 gnd.n5987 gnd.n5986 240.244
R6013 gnd.n5984 gnd.n4810 240.244
R6014 gnd.n5980 gnd.n5979 240.244
R6015 gnd.n5977 gnd.n4820 240.244
R6016 gnd.n5274 gnd.n5171 240.244
R6017 gnd.n5274 gnd.n5164 240.244
R6018 gnd.n5285 gnd.n5164 240.244
R6019 gnd.n5285 gnd.n5160 240.244
R6020 gnd.n5291 gnd.n5160 240.244
R6021 gnd.n5291 gnd.n5152 240.244
R6022 gnd.n5301 gnd.n5152 240.244
R6023 gnd.n5301 gnd.n5147 240.244
R6024 gnd.n5337 gnd.n5147 240.244
R6025 gnd.n5337 gnd.n5148 240.244
R6026 gnd.n5148 gnd.n5095 240.244
R6027 gnd.n5332 gnd.n5095 240.244
R6028 gnd.n5332 gnd.n5331 240.244
R6029 gnd.n5331 gnd.n5074 240.244
R6030 gnd.n5327 gnd.n5074 240.244
R6031 gnd.n5327 gnd.n5065 240.244
R6032 gnd.n5324 gnd.n5065 240.244
R6033 gnd.n5324 gnd.n5323 240.244
R6034 gnd.n5323 gnd.n5048 240.244
R6035 gnd.n5319 gnd.n5048 240.244
R6036 gnd.n5319 gnd.n5037 240.244
R6037 gnd.n5037 gnd.n5018 240.244
R6038 gnd.n5432 gnd.n5018 240.244
R6039 gnd.n5432 gnd.n5014 240.244
R6040 gnd.n5440 gnd.n5014 240.244
R6041 gnd.n5440 gnd.n5005 240.244
R6042 gnd.n5005 gnd.n4941 240.244
R6043 gnd.n5512 gnd.n4941 240.244
R6044 gnd.n5512 gnd.n4942 240.244
R6045 gnd.n4953 gnd.n4942 240.244
R6046 gnd.n4988 gnd.n4953 240.244
R6047 gnd.n4991 gnd.n4988 240.244
R6048 gnd.n4991 gnd.n4965 240.244
R6049 gnd.n4978 gnd.n4965 240.244
R6050 gnd.n4978 gnd.n4975 240.244
R6051 gnd.n4975 gnd.n4896 240.244
R6052 gnd.n5533 gnd.n4896 240.244
R6053 gnd.n5533 gnd.n4886 240.244
R6054 gnd.n5529 gnd.n4886 240.244
R6055 gnd.n5529 gnd.n4880 240.244
R6056 gnd.n5526 gnd.n4880 240.244
R6057 gnd.n5526 gnd.n4869 240.244
R6058 gnd.n5523 gnd.n4869 240.244
R6059 gnd.n5523 gnd.n4847 240.244
R6060 gnd.n5601 gnd.n4847 240.244
R6061 gnd.n5601 gnd.n4843 240.244
R6062 gnd.n5631 gnd.n4843 240.244
R6063 gnd.n5631 gnd.n932 240.244
R6064 gnd.n5627 gnd.n932 240.244
R6065 gnd.n5627 gnd.n942 240.244
R6066 gnd.n5624 gnd.n942 240.244
R6067 gnd.n5624 gnd.n5620 240.244
R6068 gnd.n5620 gnd.n954 240.244
R6069 gnd.n5616 gnd.n954 240.244
R6070 gnd.n5616 gnd.n965 240.244
R6071 gnd.n5949 gnd.n965 240.244
R6072 gnd.n5950 gnd.n5949 240.244
R6073 gnd.n5950 gnd.n979 240.244
R6074 gnd.n5956 gnd.n979 240.244
R6075 gnd.n5956 gnd.n990 240.244
R6076 gnd.n5960 gnd.n990 240.244
R6077 gnd.n5960 gnd.n5959 240.244
R6078 gnd.n5959 gnd.n1005 240.244
R6079 gnd.n5967 gnd.n1005 240.244
R6080 gnd.n5967 gnd.n1015 240.244
R6081 gnd.n5188 gnd.n5187 240.244
R6082 gnd.n5259 gnd.n5187 240.244
R6083 gnd.n5257 gnd.n5256 240.244
R6084 gnd.n5253 gnd.n5252 240.244
R6085 gnd.n5249 gnd.n5248 240.244
R6086 gnd.n5245 gnd.n5244 240.244
R6087 gnd.n5241 gnd.n5240 240.244
R6088 gnd.n5237 gnd.n5236 240.244
R6089 gnd.n5233 gnd.n5232 240.244
R6090 gnd.n5229 gnd.n5228 240.244
R6091 gnd.n5225 gnd.n5224 240.244
R6092 gnd.n5221 gnd.n5220 240.244
R6093 gnd.n5217 gnd.n5175 240.244
R6094 gnd.n5277 gnd.n5169 240.244
R6095 gnd.n5277 gnd.n5165 240.244
R6096 gnd.n5283 gnd.n5165 240.244
R6097 gnd.n5283 gnd.n5158 240.244
R6098 gnd.n5293 gnd.n5158 240.244
R6099 gnd.n5293 gnd.n5154 240.244
R6100 gnd.n5299 gnd.n5154 240.244
R6101 gnd.n5299 gnd.n5145 240.244
R6102 gnd.n5339 gnd.n5145 240.244
R6103 gnd.n5339 gnd.n5096 240.244
R6104 gnd.n5347 gnd.n5096 240.244
R6105 gnd.n5347 gnd.n5097 240.244
R6106 gnd.n5097 gnd.n5075 240.244
R6107 gnd.n5368 gnd.n5075 240.244
R6108 gnd.n5368 gnd.n5067 240.244
R6109 gnd.n5379 gnd.n5067 240.244
R6110 gnd.n5379 gnd.n5068 240.244
R6111 gnd.n5068 gnd.n5049 240.244
R6112 gnd.n5399 gnd.n5049 240.244
R6113 gnd.n5399 gnd.n5039 240.244
R6114 gnd.n5409 gnd.n5039 240.244
R6115 gnd.n5409 gnd.n5020 240.244
R6116 gnd.n5430 gnd.n5020 240.244
R6117 gnd.n5430 gnd.n5022 240.244
R6118 gnd.n5022 gnd.n5003 240.244
R6119 gnd.n5458 gnd.n5003 240.244
R6120 gnd.n5458 gnd.n4945 240.244
R6121 gnd.n5510 gnd.n4945 240.244
R6122 gnd.n5510 gnd.n4946 240.244
R6123 gnd.n5506 gnd.n4946 240.244
R6124 gnd.n5506 gnd.n4952 240.244
R6125 gnd.n4967 gnd.n4952 240.244
R6126 gnd.n5496 gnd.n4967 240.244
R6127 gnd.n5496 gnd.n4968 240.244
R6128 gnd.n5492 gnd.n4968 240.244
R6129 gnd.n5492 gnd.n4974 240.244
R6130 gnd.n4974 gnd.n4885 240.244
R6131 gnd.n5549 gnd.n4885 240.244
R6132 gnd.n5549 gnd.n4878 240.244
R6133 gnd.n5560 gnd.n4878 240.244
R6134 gnd.n5560 gnd.n4871 240.244
R6135 gnd.n5575 gnd.n4871 240.244
R6136 gnd.n5575 gnd.n4872 240.244
R6137 gnd.n4872 gnd.n4850 240.244
R6138 gnd.n5599 gnd.n4850 240.244
R6139 gnd.n5599 gnd.n4851 240.244
R6140 gnd.n4851 gnd.n933 240.244
R6141 gnd.n6103 gnd.n933 240.244
R6142 gnd.n6103 gnd.n934 240.244
R6143 gnd.n6099 gnd.n934 240.244
R6144 gnd.n6099 gnd.n940 240.244
R6145 gnd.n956 gnd.n940 240.244
R6146 gnd.n6089 gnd.n956 240.244
R6147 gnd.n6089 gnd.n957 240.244
R6148 gnd.n6085 gnd.n957 240.244
R6149 gnd.n6085 gnd.n963 240.244
R6150 gnd.n981 gnd.n963 240.244
R6151 gnd.n6075 gnd.n981 240.244
R6152 gnd.n6075 gnd.n982 240.244
R6153 gnd.n6071 gnd.n982 240.244
R6154 gnd.n6071 gnd.n988 240.244
R6155 gnd.n1007 gnd.n988 240.244
R6156 gnd.n6061 gnd.n1007 240.244
R6157 gnd.n6061 gnd.n1008 240.244
R6158 gnd.n6057 gnd.n1008 240.244
R6159 gnd.n7179 gnd.n7178 240.244
R6160 gnd.n7184 gnd.n7181 240.244
R6161 gnd.n7187 gnd.n7186 240.244
R6162 gnd.n7192 gnd.n7189 240.244
R6163 gnd.n7195 gnd.n7194 240.244
R6164 gnd.n7200 gnd.n7197 240.244
R6165 gnd.n7203 gnd.n7202 240.244
R6166 gnd.n7208 gnd.n7205 240.244
R6167 gnd.n7214 gnd.n7210 240.244
R6168 gnd.n4147 gnd.n1461 240.244
R6169 gnd.n4147 gnd.n1473 240.244
R6170 gnd.n4177 gnd.n1473 240.244
R6171 gnd.n4177 gnd.n1588 240.244
R6172 gnd.n4184 gnd.n1588 240.244
R6173 gnd.n4184 gnd.n1566 240.244
R6174 gnd.n1566 gnd.n1554 240.244
R6175 gnd.n4208 gnd.n1554 240.244
R6176 gnd.n4208 gnd.n1549 240.244
R6177 gnd.n4221 gnd.n1549 240.244
R6178 gnd.n4221 gnd.n1541 240.244
R6179 gnd.n4214 gnd.n1541 240.244
R6180 gnd.n4214 gnd.n1531 240.244
R6181 gnd.n1531 gnd.n1504 240.244
R6182 gnd.n4325 gnd.n1504 240.244
R6183 gnd.n4325 gnd.n1498 240.244
R6184 gnd.n1509 gnd.n1498 240.244
R6185 gnd.n1509 gnd.n235 240.244
R6186 gnd.n1510 gnd.n235 240.244
R6187 gnd.n4315 gnd.n1510 240.244
R6188 gnd.n4315 gnd.n1511 240.244
R6189 gnd.n1511 gnd.n54 240.244
R6190 gnd.n55 gnd.n54 240.244
R6191 gnd.n56 gnd.n55 240.244
R6192 gnd.n250 gnd.n56 240.244
R6193 gnd.n250 gnd.n59 240.244
R6194 gnd.n60 gnd.n59 240.244
R6195 gnd.n61 gnd.n60 240.244
R6196 gnd.n213 gnd.n61 240.244
R6197 gnd.n213 gnd.n64 240.244
R6198 gnd.n65 gnd.n64 240.244
R6199 gnd.n66 gnd.n65 240.244
R6200 gnd.n196 gnd.n66 240.244
R6201 gnd.n196 gnd.n69 240.244
R6202 gnd.n70 gnd.n69 240.244
R6203 gnd.n71 gnd.n70 240.244
R6204 gnd.n181 gnd.n71 240.244
R6205 gnd.n181 gnd.n74 240.244
R6206 gnd.n75 gnd.n74 240.244
R6207 gnd.n76 gnd.n75 240.244
R6208 gnd.n79 gnd.n76 240.244
R6209 gnd.n7327 gnd.n79 240.244
R6210 gnd.n1653 gnd.n1651 240.244
R6211 gnd.n1668 gnd.n1634 240.244
R6212 gnd.n1672 gnd.n1670 240.244
R6213 gnd.n1687 gnd.n1625 240.244
R6214 gnd.n1691 gnd.n1689 240.244
R6215 gnd.n1706 gnd.n1616 240.244
R6216 gnd.n1710 gnd.n1708 240.244
R6217 gnd.n1725 gnd.n1607 240.244
R6218 gnd.n1728 gnd.n1727 240.244
R6219 gnd.n1475 gnd.n1463 240.244
R6220 gnd.n4354 gnd.n1475 240.244
R6221 gnd.n4354 gnd.n1476 240.244
R6222 gnd.n1481 gnd.n1476 240.244
R6223 gnd.n1482 gnd.n1481 240.244
R6224 gnd.n1483 gnd.n1482 240.244
R6225 gnd.n1567 gnd.n1483 240.244
R6226 gnd.n1567 gnd.n1486 240.244
R6227 gnd.n1487 gnd.n1486 240.244
R6228 gnd.n1488 gnd.n1487 240.244
R6229 gnd.n4249 gnd.n1488 240.244
R6230 gnd.n4249 gnd.n1491 240.244
R6231 gnd.n1492 gnd.n1491 240.244
R6232 gnd.n1493 gnd.n1492 240.244
R6233 gnd.n1495 gnd.n1493 240.244
R6234 gnd.n4330 gnd.n1495 240.244
R6235 gnd.n4330 gnd.n237 240.244
R6236 gnd.n7112 gnd.n237 240.244
R6237 gnd.n7112 gnd.n238 240.244
R6238 gnd.n243 gnd.n238 240.244
R6239 gnd.n244 gnd.n243 240.244
R6240 gnd.n245 gnd.n244 240.244
R6241 gnd.n4289 gnd.n245 240.244
R6242 gnd.n4289 gnd.n248 240.244
R6243 gnd.n7099 gnd.n248 240.244
R6244 gnd.n7099 gnd.n219 240.244
R6245 gnd.n7123 gnd.n219 240.244
R6246 gnd.n7123 gnd.n215 240.244
R6247 gnd.n7129 gnd.n215 240.244
R6248 gnd.n7129 gnd.n202 240.244
R6249 gnd.n7139 gnd.n202 240.244
R6250 gnd.n7139 gnd.n198 240.244
R6251 gnd.n7145 gnd.n198 240.244
R6252 gnd.n7145 gnd.n187 240.244
R6253 gnd.n7155 gnd.n187 240.244
R6254 gnd.n7155 gnd.n183 240.244
R6255 gnd.n7161 gnd.n183 240.244
R6256 gnd.n7161 gnd.n168 240.244
R6257 gnd.n7173 gnd.n168 240.244
R6258 gnd.n7173 gnd.n163 240.244
R6259 gnd.n7246 gnd.n163 240.244
R6260 gnd.n7246 gnd.n84 240.244
R6261 gnd.n3018 gnd.n1330 240.244
R6262 gnd.n3021 gnd.n3020 240.244
R6263 gnd.n3031 gnd.n3023 240.244
R6264 gnd.n3034 gnd.n3033 240.244
R6265 gnd.n3043 gnd.n3042 240.244
R6266 gnd.n3054 gnd.n3045 240.244
R6267 gnd.n3057 gnd.n3056 240.244
R6268 gnd.n3066 gnd.n3065 240.244
R6269 gnd.n3077 gnd.n3068 240.244
R6270 gnd.n2669 gnd.n1120 240.244
R6271 gnd.n2752 gnd.n2669 240.244
R6272 gnd.n2752 gnd.n1132 240.244
R6273 gnd.n2748 gnd.n1132 240.244
R6274 gnd.n2748 gnd.n1144 240.244
R6275 gnd.n2655 gnd.n1144 240.244
R6276 gnd.n2655 gnd.n1153 240.244
R6277 gnd.n2809 gnd.n1153 240.244
R6278 gnd.n2809 gnd.n1164 240.244
R6279 gnd.n2815 gnd.n1164 240.244
R6280 gnd.n2815 gnd.n1174 240.244
R6281 gnd.n2826 gnd.n1174 240.244
R6282 gnd.n2826 gnd.n1185 240.244
R6283 gnd.n2835 gnd.n1185 240.244
R6284 gnd.n2835 gnd.n1195 240.244
R6285 gnd.n2613 gnd.n1195 240.244
R6286 gnd.n2892 gnd.n2613 240.244
R6287 gnd.n2892 gnd.n1206 240.244
R6288 gnd.n2888 gnd.n1206 240.244
R6289 gnd.n2888 gnd.n1219 240.244
R6290 gnd.n2853 gnd.n1219 240.244
R6291 gnd.n2853 gnd.n1227 240.244
R6292 gnd.n2875 gnd.n1227 240.244
R6293 gnd.n2875 gnd.n1236 240.244
R6294 gnd.n2869 gnd.n1236 240.244
R6295 gnd.n2869 gnd.n1244 240.244
R6296 gnd.n2908 gnd.n1244 240.244
R6297 gnd.n2908 gnd.n1254 240.244
R6298 gnd.n2914 gnd.n1254 240.244
R6299 gnd.n2914 gnd.n1265 240.244
R6300 gnd.n2959 gnd.n1265 240.244
R6301 gnd.n2959 gnd.n1275 240.244
R6302 gnd.n2582 gnd.n1275 240.244
R6303 gnd.n2582 gnd.n1286 240.244
R6304 gnd.n2583 gnd.n1286 240.244
R6305 gnd.n2583 gnd.n1296 240.244
R6306 gnd.n2586 gnd.n1296 240.244
R6307 gnd.n2586 gnd.n1307 240.244
R6308 gnd.n2944 gnd.n1307 240.244
R6309 gnd.n2944 gnd.n1318 240.244
R6310 gnd.n3238 gnd.n1318 240.244
R6311 gnd.n3238 gnd.n1328 240.244
R6312 gnd.n2689 gnd.n2688 240.244
R6313 gnd.n2695 gnd.n2694 240.244
R6314 gnd.n2699 gnd.n2698 240.244
R6315 gnd.n2705 gnd.n2704 240.244
R6316 gnd.n2709 gnd.n2708 240.244
R6317 gnd.n2715 gnd.n2714 240.244
R6318 gnd.n2719 gnd.n2718 240.244
R6319 gnd.n2677 gnd.n2676 240.244
R6320 gnd.n2672 gnd.n1068 240.244
R6321 gnd.n4634 gnd.n1123 240.244
R6322 gnd.n1128 gnd.n1123 240.244
R6323 gnd.n4627 gnd.n1128 240.244
R6324 gnd.n4627 gnd.n1129 240.244
R6325 gnd.n4619 gnd.n1129 240.244
R6326 gnd.n4619 gnd.n1146 240.244
R6327 gnd.n4615 gnd.n1146 240.244
R6328 gnd.n4615 gnd.n1151 240.244
R6329 gnd.n4607 gnd.n1151 240.244
R6330 gnd.n4607 gnd.n1165 240.244
R6331 gnd.n4603 gnd.n1165 240.244
R6332 gnd.n4603 gnd.n1171 240.244
R6333 gnd.n4595 gnd.n1171 240.244
R6334 gnd.n4595 gnd.n1187 240.244
R6335 gnd.n4591 gnd.n1187 240.244
R6336 gnd.n4591 gnd.n1193 240.244
R6337 gnd.n1208 gnd.n1193 240.244
R6338 gnd.n4581 gnd.n1208 240.244
R6339 gnd.n4581 gnd.n1209 240.244
R6340 gnd.n4577 gnd.n1209 240.244
R6341 gnd.n4577 gnd.n1217 240.244
R6342 gnd.n4568 gnd.n1217 240.244
R6343 gnd.n4568 gnd.n1228 240.244
R6344 gnd.n4564 gnd.n1228 240.244
R6345 gnd.n4564 gnd.n1233 240.244
R6346 gnd.n4555 gnd.n1233 240.244
R6347 gnd.n4555 gnd.n1246 240.244
R6348 gnd.n4551 gnd.n1246 240.244
R6349 gnd.n4551 gnd.n1252 240.244
R6350 gnd.n4543 gnd.n1252 240.244
R6351 gnd.n4543 gnd.n1266 240.244
R6352 gnd.n4539 gnd.n1266 240.244
R6353 gnd.n4539 gnd.n1272 240.244
R6354 gnd.n4531 gnd.n1272 240.244
R6355 gnd.n4531 gnd.n1288 240.244
R6356 gnd.n4527 gnd.n1288 240.244
R6357 gnd.n4527 gnd.n1294 240.244
R6358 gnd.n4519 gnd.n1294 240.244
R6359 gnd.n4519 gnd.n1309 240.244
R6360 gnd.n4515 gnd.n1309 240.244
R6361 gnd.n4515 gnd.n1315 240.244
R6362 gnd.n4507 gnd.n1315 240.244
R6363 gnd.n6275 gnd.n759 240.244
R6364 gnd.n6281 gnd.n759 240.244
R6365 gnd.n6281 gnd.n757 240.244
R6366 gnd.n6285 gnd.n757 240.244
R6367 gnd.n6285 gnd.n753 240.244
R6368 gnd.n6291 gnd.n753 240.244
R6369 gnd.n6291 gnd.n751 240.244
R6370 gnd.n6295 gnd.n751 240.244
R6371 gnd.n6295 gnd.n747 240.244
R6372 gnd.n6301 gnd.n747 240.244
R6373 gnd.n6301 gnd.n745 240.244
R6374 gnd.n6305 gnd.n745 240.244
R6375 gnd.n6305 gnd.n741 240.244
R6376 gnd.n6311 gnd.n741 240.244
R6377 gnd.n6311 gnd.n739 240.244
R6378 gnd.n6315 gnd.n739 240.244
R6379 gnd.n6315 gnd.n735 240.244
R6380 gnd.n6321 gnd.n735 240.244
R6381 gnd.n6321 gnd.n733 240.244
R6382 gnd.n6325 gnd.n733 240.244
R6383 gnd.n6325 gnd.n729 240.244
R6384 gnd.n6331 gnd.n729 240.244
R6385 gnd.n6331 gnd.n727 240.244
R6386 gnd.n6335 gnd.n727 240.244
R6387 gnd.n6335 gnd.n723 240.244
R6388 gnd.n6341 gnd.n723 240.244
R6389 gnd.n6341 gnd.n721 240.244
R6390 gnd.n6345 gnd.n721 240.244
R6391 gnd.n6345 gnd.n717 240.244
R6392 gnd.n6351 gnd.n717 240.244
R6393 gnd.n6351 gnd.n715 240.244
R6394 gnd.n6355 gnd.n715 240.244
R6395 gnd.n6355 gnd.n711 240.244
R6396 gnd.n6361 gnd.n711 240.244
R6397 gnd.n6361 gnd.n709 240.244
R6398 gnd.n6365 gnd.n709 240.244
R6399 gnd.n6365 gnd.n705 240.244
R6400 gnd.n6371 gnd.n705 240.244
R6401 gnd.n6371 gnd.n703 240.244
R6402 gnd.n6375 gnd.n703 240.244
R6403 gnd.n6375 gnd.n699 240.244
R6404 gnd.n6381 gnd.n699 240.244
R6405 gnd.n6381 gnd.n697 240.244
R6406 gnd.n6385 gnd.n697 240.244
R6407 gnd.n6385 gnd.n693 240.244
R6408 gnd.n6391 gnd.n693 240.244
R6409 gnd.n6391 gnd.n691 240.244
R6410 gnd.n6395 gnd.n691 240.244
R6411 gnd.n6395 gnd.n687 240.244
R6412 gnd.n6401 gnd.n687 240.244
R6413 gnd.n6401 gnd.n685 240.244
R6414 gnd.n6405 gnd.n685 240.244
R6415 gnd.n6405 gnd.n681 240.244
R6416 gnd.n6411 gnd.n681 240.244
R6417 gnd.n6411 gnd.n679 240.244
R6418 gnd.n6415 gnd.n679 240.244
R6419 gnd.n6415 gnd.n675 240.244
R6420 gnd.n6421 gnd.n675 240.244
R6421 gnd.n6421 gnd.n673 240.244
R6422 gnd.n6425 gnd.n673 240.244
R6423 gnd.n6425 gnd.n669 240.244
R6424 gnd.n6431 gnd.n669 240.244
R6425 gnd.n6431 gnd.n667 240.244
R6426 gnd.n6435 gnd.n667 240.244
R6427 gnd.n6435 gnd.n663 240.244
R6428 gnd.n6441 gnd.n663 240.244
R6429 gnd.n6441 gnd.n661 240.244
R6430 gnd.n6445 gnd.n661 240.244
R6431 gnd.n6445 gnd.n657 240.244
R6432 gnd.n6451 gnd.n657 240.244
R6433 gnd.n6451 gnd.n655 240.244
R6434 gnd.n6455 gnd.n655 240.244
R6435 gnd.n6455 gnd.n651 240.244
R6436 gnd.n6461 gnd.n651 240.244
R6437 gnd.n6461 gnd.n649 240.244
R6438 gnd.n6465 gnd.n649 240.244
R6439 gnd.n6465 gnd.n645 240.244
R6440 gnd.n6471 gnd.n645 240.244
R6441 gnd.n6471 gnd.n643 240.244
R6442 gnd.n6475 gnd.n643 240.244
R6443 gnd.n6475 gnd.n639 240.244
R6444 gnd.n6481 gnd.n639 240.244
R6445 gnd.n6481 gnd.n637 240.244
R6446 gnd.n6485 gnd.n637 240.244
R6447 gnd.n6485 gnd.n633 240.244
R6448 gnd.n6491 gnd.n633 240.244
R6449 gnd.n6491 gnd.n631 240.244
R6450 gnd.n6495 gnd.n631 240.244
R6451 gnd.n6495 gnd.n627 240.244
R6452 gnd.n6501 gnd.n627 240.244
R6453 gnd.n6501 gnd.n625 240.244
R6454 gnd.n6505 gnd.n625 240.244
R6455 gnd.n6505 gnd.n621 240.244
R6456 gnd.n6511 gnd.n621 240.244
R6457 gnd.n6511 gnd.n619 240.244
R6458 gnd.n6515 gnd.n619 240.244
R6459 gnd.n6515 gnd.n615 240.244
R6460 gnd.n6521 gnd.n615 240.244
R6461 gnd.n6521 gnd.n613 240.244
R6462 gnd.n6525 gnd.n613 240.244
R6463 gnd.n6525 gnd.n609 240.244
R6464 gnd.n6531 gnd.n609 240.244
R6465 gnd.n6531 gnd.n607 240.244
R6466 gnd.n6535 gnd.n607 240.244
R6467 gnd.n6535 gnd.n603 240.244
R6468 gnd.n6541 gnd.n603 240.244
R6469 gnd.n6541 gnd.n601 240.244
R6470 gnd.n6545 gnd.n601 240.244
R6471 gnd.n6545 gnd.n597 240.244
R6472 gnd.n6551 gnd.n597 240.244
R6473 gnd.n6551 gnd.n595 240.244
R6474 gnd.n6555 gnd.n595 240.244
R6475 gnd.n6555 gnd.n591 240.244
R6476 gnd.n6561 gnd.n591 240.244
R6477 gnd.n6561 gnd.n589 240.244
R6478 gnd.n6565 gnd.n589 240.244
R6479 gnd.n6565 gnd.n585 240.244
R6480 gnd.n6571 gnd.n585 240.244
R6481 gnd.n6571 gnd.n583 240.244
R6482 gnd.n6575 gnd.n583 240.244
R6483 gnd.n6575 gnd.n579 240.244
R6484 gnd.n6581 gnd.n579 240.244
R6485 gnd.n6581 gnd.n577 240.244
R6486 gnd.n6585 gnd.n577 240.244
R6487 gnd.n6585 gnd.n573 240.244
R6488 gnd.n6591 gnd.n573 240.244
R6489 gnd.n6591 gnd.n571 240.244
R6490 gnd.n6595 gnd.n571 240.244
R6491 gnd.n6595 gnd.n567 240.244
R6492 gnd.n6601 gnd.n567 240.244
R6493 gnd.n6601 gnd.n565 240.244
R6494 gnd.n6605 gnd.n565 240.244
R6495 gnd.n6605 gnd.n561 240.244
R6496 gnd.n6611 gnd.n561 240.244
R6497 gnd.n6611 gnd.n559 240.244
R6498 gnd.n6615 gnd.n559 240.244
R6499 gnd.n6615 gnd.n555 240.244
R6500 gnd.n6621 gnd.n555 240.244
R6501 gnd.n6621 gnd.n553 240.244
R6502 gnd.n6625 gnd.n553 240.244
R6503 gnd.n6625 gnd.n549 240.244
R6504 gnd.n6631 gnd.n549 240.244
R6505 gnd.n6631 gnd.n547 240.244
R6506 gnd.n6635 gnd.n547 240.244
R6507 gnd.n6635 gnd.n543 240.244
R6508 gnd.n6641 gnd.n543 240.244
R6509 gnd.n6641 gnd.n541 240.244
R6510 gnd.n6645 gnd.n541 240.244
R6511 gnd.n6645 gnd.n537 240.244
R6512 gnd.n6651 gnd.n537 240.244
R6513 gnd.n6651 gnd.n535 240.244
R6514 gnd.n6655 gnd.n535 240.244
R6515 gnd.n6655 gnd.n531 240.244
R6516 gnd.n6661 gnd.n531 240.244
R6517 gnd.n6661 gnd.n529 240.244
R6518 gnd.n6665 gnd.n529 240.244
R6519 gnd.n6665 gnd.n525 240.244
R6520 gnd.n6671 gnd.n525 240.244
R6521 gnd.n6671 gnd.n523 240.244
R6522 gnd.n6675 gnd.n523 240.244
R6523 gnd.n6675 gnd.n519 240.244
R6524 gnd.n6681 gnd.n519 240.244
R6525 gnd.n6681 gnd.n517 240.244
R6526 gnd.n6685 gnd.n517 240.244
R6527 gnd.n6685 gnd.n513 240.244
R6528 gnd.n6691 gnd.n513 240.244
R6529 gnd.n6691 gnd.n511 240.244
R6530 gnd.n6695 gnd.n511 240.244
R6531 gnd.n6695 gnd.n507 240.244
R6532 gnd.n6701 gnd.n507 240.244
R6533 gnd.n6701 gnd.n505 240.244
R6534 gnd.n6705 gnd.n505 240.244
R6535 gnd.n6705 gnd.n501 240.244
R6536 gnd.n6711 gnd.n501 240.244
R6537 gnd.n6711 gnd.n499 240.244
R6538 gnd.n6715 gnd.n499 240.244
R6539 gnd.n6715 gnd.n495 240.244
R6540 gnd.n6721 gnd.n495 240.244
R6541 gnd.n6721 gnd.n493 240.244
R6542 gnd.n6725 gnd.n493 240.244
R6543 gnd.n6725 gnd.n489 240.244
R6544 gnd.n6731 gnd.n489 240.244
R6545 gnd.n6731 gnd.n487 240.244
R6546 gnd.n6735 gnd.n487 240.244
R6547 gnd.n6735 gnd.n483 240.244
R6548 gnd.n6741 gnd.n483 240.244
R6549 gnd.n6741 gnd.n481 240.244
R6550 gnd.n6745 gnd.n481 240.244
R6551 gnd.n6745 gnd.n477 240.244
R6552 gnd.n6751 gnd.n477 240.244
R6553 gnd.n6751 gnd.n475 240.244
R6554 gnd.n6755 gnd.n475 240.244
R6555 gnd.n6755 gnd.n471 240.244
R6556 gnd.n6761 gnd.n471 240.244
R6557 gnd.n6761 gnd.n469 240.244
R6558 gnd.n6765 gnd.n469 240.244
R6559 gnd.n6765 gnd.n465 240.244
R6560 gnd.n6771 gnd.n465 240.244
R6561 gnd.n6771 gnd.n463 240.244
R6562 gnd.n6775 gnd.n463 240.244
R6563 gnd.n6775 gnd.n459 240.244
R6564 gnd.n6781 gnd.n459 240.244
R6565 gnd.n6781 gnd.n457 240.244
R6566 gnd.n6785 gnd.n457 240.244
R6567 gnd.n6785 gnd.n453 240.244
R6568 gnd.n6792 gnd.n453 240.244
R6569 gnd.n6792 gnd.n451 240.244
R6570 gnd.n6796 gnd.n448 240.244
R6571 gnd.n6802 gnd.n448 240.244
R6572 gnd.n6802 gnd.n446 240.244
R6573 gnd.n6806 gnd.n446 240.244
R6574 gnd.n6806 gnd.n442 240.244
R6575 gnd.n6812 gnd.n442 240.244
R6576 gnd.n6812 gnd.n440 240.244
R6577 gnd.n6816 gnd.n440 240.244
R6578 gnd.n6816 gnd.n436 240.244
R6579 gnd.n6822 gnd.n436 240.244
R6580 gnd.n6822 gnd.n434 240.244
R6581 gnd.n6826 gnd.n434 240.244
R6582 gnd.n6826 gnd.n430 240.244
R6583 gnd.n6832 gnd.n430 240.244
R6584 gnd.n6832 gnd.n428 240.244
R6585 gnd.n6836 gnd.n428 240.244
R6586 gnd.n6836 gnd.n424 240.244
R6587 gnd.n6842 gnd.n424 240.244
R6588 gnd.n6842 gnd.n422 240.244
R6589 gnd.n6846 gnd.n422 240.244
R6590 gnd.n6846 gnd.n418 240.244
R6591 gnd.n6852 gnd.n418 240.244
R6592 gnd.n6852 gnd.n416 240.244
R6593 gnd.n6856 gnd.n416 240.244
R6594 gnd.n6856 gnd.n412 240.244
R6595 gnd.n6862 gnd.n412 240.244
R6596 gnd.n6862 gnd.n410 240.244
R6597 gnd.n6866 gnd.n410 240.244
R6598 gnd.n6866 gnd.n406 240.244
R6599 gnd.n6872 gnd.n406 240.244
R6600 gnd.n6872 gnd.n404 240.244
R6601 gnd.n6876 gnd.n404 240.244
R6602 gnd.n6876 gnd.n400 240.244
R6603 gnd.n6882 gnd.n400 240.244
R6604 gnd.n6882 gnd.n398 240.244
R6605 gnd.n6886 gnd.n398 240.244
R6606 gnd.n6886 gnd.n394 240.244
R6607 gnd.n6892 gnd.n394 240.244
R6608 gnd.n6892 gnd.n392 240.244
R6609 gnd.n6896 gnd.n392 240.244
R6610 gnd.n6896 gnd.n388 240.244
R6611 gnd.n6902 gnd.n388 240.244
R6612 gnd.n6902 gnd.n386 240.244
R6613 gnd.n6906 gnd.n386 240.244
R6614 gnd.n6906 gnd.n382 240.244
R6615 gnd.n6912 gnd.n382 240.244
R6616 gnd.n6912 gnd.n380 240.244
R6617 gnd.n6916 gnd.n380 240.244
R6618 gnd.n6916 gnd.n376 240.244
R6619 gnd.n6922 gnd.n376 240.244
R6620 gnd.n6922 gnd.n374 240.244
R6621 gnd.n6926 gnd.n374 240.244
R6622 gnd.n6926 gnd.n370 240.244
R6623 gnd.n6932 gnd.n370 240.244
R6624 gnd.n6932 gnd.n368 240.244
R6625 gnd.n6936 gnd.n368 240.244
R6626 gnd.n6936 gnd.n364 240.244
R6627 gnd.n6942 gnd.n364 240.244
R6628 gnd.n6942 gnd.n362 240.244
R6629 gnd.n6946 gnd.n362 240.244
R6630 gnd.n6946 gnd.n358 240.244
R6631 gnd.n6952 gnd.n358 240.244
R6632 gnd.n6952 gnd.n356 240.244
R6633 gnd.n6956 gnd.n356 240.244
R6634 gnd.n6956 gnd.n352 240.244
R6635 gnd.n6962 gnd.n352 240.244
R6636 gnd.n6962 gnd.n350 240.244
R6637 gnd.n6966 gnd.n350 240.244
R6638 gnd.n6966 gnd.n346 240.244
R6639 gnd.n6972 gnd.n346 240.244
R6640 gnd.n6972 gnd.n344 240.244
R6641 gnd.n6976 gnd.n344 240.244
R6642 gnd.n6976 gnd.n340 240.244
R6643 gnd.n6982 gnd.n340 240.244
R6644 gnd.n6982 gnd.n338 240.244
R6645 gnd.n6986 gnd.n338 240.244
R6646 gnd.n6986 gnd.n334 240.244
R6647 gnd.n6992 gnd.n334 240.244
R6648 gnd.n6992 gnd.n332 240.244
R6649 gnd.n6996 gnd.n332 240.244
R6650 gnd.n6996 gnd.n328 240.244
R6651 gnd.n7002 gnd.n328 240.244
R6652 gnd.n7002 gnd.n326 240.244
R6653 gnd.n7006 gnd.n326 240.244
R6654 gnd.n4738 gnd.n1018 240.244
R6655 gnd.n4734 gnd.n1018 240.244
R6656 gnd.n4734 gnd.n1024 240.244
R6657 gnd.n4730 gnd.n1024 240.244
R6658 gnd.n4730 gnd.n1026 240.244
R6659 gnd.n4726 gnd.n1026 240.244
R6660 gnd.n4726 gnd.n1032 240.244
R6661 gnd.n4722 gnd.n1032 240.244
R6662 gnd.n4722 gnd.n1034 240.244
R6663 gnd.n4718 gnd.n1034 240.244
R6664 gnd.n4718 gnd.n1040 240.244
R6665 gnd.n2762 gnd.n1040 240.244
R6666 gnd.n2763 gnd.n2762 240.244
R6667 gnd.n2764 gnd.n2763 240.244
R6668 gnd.n2764 gnd.n2755 240.244
R6669 gnd.n2770 gnd.n2755 240.244
R6670 gnd.n2771 gnd.n2770 240.244
R6671 gnd.n2772 gnd.n2771 240.244
R6672 gnd.n2772 gnd.n2656 240.244
R6673 gnd.n2798 gnd.n2656 240.244
R6674 gnd.n2798 gnd.n2657 240.244
R6675 gnd.n2794 gnd.n2657 240.244
R6676 gnd.n2794 gnd.n2793 240.244
R6677 gnd.n2793 gnd.n2792 240.244
R6678 gnd.n2792 gnd.n2780 240.244
R6679 gnd.n2788 gnd.n2780 240.244
R6680 gnd.n2788 gnd.n2787 240.244
R6681 gnd.n2787 gnd.n2609 240.244
R6682 gnd.n2896 gnd.n2609 240.244
R6683 gnd.n2896 gnd.n2895 240.244
R6684 gnd.n2895 gnd.n2610 240.244
R6685 gnd.n2622 gnd.n2610 240.244
R6686 gnd.n2885 gnd.n2622 240.244
R6687 gnd.n2885 gnd.n2882 240.244
R6688 gnd.n2882 gnd.n2881 240.244
R6689 gnd.n2881 gnd.n2878 240.244
R6690 gnd.n2878 gnd.n2628 240.244
R6691 gnd.n2628 gnd.n2625 240.244
R6692 gnd.n2625 gnd.n2624 240.244
R6693 gnd.n2624 gnd.n2598 240.244
R6694 gnd.n2905 gnd.n2598 240.244
R6695 gnd.n2905 gnd.n2599 240.244
R6696 gnd.n2599 gnd.n2576 240.244
R6697 gnd.n2962 gnd.n2576 240.244
R6698 gnd.n2962 gnd.n2572 240.244
R6699 gnd.n2968 gnd.n2572 240.244
R6700 gnd.n2969 gnd.n2968 240.244
R6701 gnd.n2970 gnd.n2969 240.244
R6702 gnd.n2970 gnd.n2568 240.244
R6703 gnd.n2976 gnd.n2568 240.244
R6704 gnd.n2977 gnd.n2976 240.244
R6705 gnd.n2978 gnd.n2977 240.244
R6706 gnd.n2978 gnd.n2564 240.244
R6707 gnd.n2984 gnd.n2564 240.244
R6708 gnd.n2985 gnd.n2984 240.244
R6709 gnd.n2986 gnd.n2985 240.244
R6710 gnd.n2986 gnd.n2560 240.244
R6711 gnd.n2992 gnd.n2560 240.244
R6712 gnd.n2992 gnd.n2558 240.244
R6713 gnd.n3129 gnd.n2558 240.244
R6714 gnd.n3129 gnd.n2554 240.244
R6715 gnd.n3135 gnd.n2554 240.244
R6716 gnd.n3135 gnd.n2552 240.244
R6717 gnd.n3143 gnd.n2552 240.244
R6718 gnd.n3143 gnd.n2548 240.244
R6719 gnd.n3149 gnd.n2548 240.244
R6720 gnd.n3149 gnd.n2544 240.244
R6721 gnd.n3157 gnd.n2544 240.244
R6722 gnd.n3157 gnd.n2540 240.244
R6723 gnd.n3163 gnd.n2540 240.244
R6724 gnd.n3163 gnd.n2536 240.244
R6725 gnd.n3171 gnd.n2536 240.244
R6726 gnd.n3171 gnd.n2532 240.244
R6727 gnd.n3177 gnd.n2532 240.244
R6728 gnd.n3177 gnd.n2259 240.244
R6729 gnd.n3360 gnd.n2259 240.244
R6730 gnd.n3360 gnd.n2255 240.244
R6731 gnd.n3366 gnd.n2255 240.244
R6732 gnd.n3366 gnd.n2241 240.244
R6733 gnd.n3451 gnd.n2241 240.244
R6734 gnd.n3451 gnd.n2237 240.244
R6735 gnd.n3457 gnd.n2237 240.244
R6736 gnd.n3457 gnd.n2220 240.244
R6737 gnd.n3482 gnd.n2220 240.244
R6738 gnd.n3482 gnd.n2216 240.244
R6739 gnd.n3488 gnd.n2216 240.244
R6740 gnd.n3488 gnd.n2198 240.244
R6741 gnd.n3510 gnd.n2198 240.244
R6742 gnd.n3510 gnd.n2193 240.244
R6743 gnd.n3518 gnd.n2193 240.244
R6744 gnd.n3518 gnd.n2194 240.244
R6745 gnd.n2194 gnd.n2169 240.244
R6746 gnd.n3547 gnd.n2169 240.244
R6747 gnd.n3547 gnd.n2165 240.244
R6748 gnd.n3553 gnd.n2165 240.244
R6749 gnd.n3553 gnd.n2146 240.244
R6750 gnd.n3575 gnd.n2146 240.244
R6751 gnd.n3575 gnd.n2141 240.244
R6752 gnd.n3583 gnd.n2141 240.244
R6753 gnd.n3583 gnd.n2142 240.244
R6754 gnd.n2142 gnd.n2117 240.244
R6755 gnd.n3626 gnd.n2117 240.244
R6756 gnd.n3626 gnd.n2113 240.244
R6757 gnd.n3632 gnd.n2113 240.244
R6758 gnd.n3632 gnd.n2096 240.244
R6759 gnd.n3656 gnd.n2096 240.244
R6760 gnd.n3656 gnd.n2091 240.244
R6761 gnd.n3664 gnd.n2091 240.244
R6762 gnd.n3664 gnd.n2092 240.244
R6763 gnd.n2092 gnd.n2066 240.244
R6764 gnd.n3706 gnd.n2066 240.244
R6765 gnd.n3706 gnd.n2062 240.244
R6766 gnd.n3712 gnd.n2062 240.244
R6767 gnd.n3712 gnd.n2043 240.244
R6768 gnd.n3746 gnd.n2043 240.244
R6769 gnd.n3746 gnd.n2039 240.244
R6770 gnd.n3752 gnd.n2039 240.244
R6771 gnd.n3752 gnd.n2020 240.244
R6772 gnd.n3785 gnd.n2020 240.244
R6773 gnd.n3785 gnd.n2016 240.244
R6774 gnd.n3791 gnd.n2016 240.244
R6775 gnd.n3791 gnd.n1998 240.244
R6776 gnd.n3826 gnd.n1998 240.244
R6777 gnd.n3826 gnd.n1994 240.244
R6778 gnd.n3832 gnd.n1994 240.244
R6779 gnd.n3832 gnd.n1976 240.244
R6780 gnd.n3871 gnd.n1976 240.244
R6781 gnd.n3871 gnd.n1971 240.244
R6782 gnd.n3883 gnd.n1971 240.244
R6783 gnd.n3883 gnd.n1972 240.244
R6784 gnd.n3879 gnd.n1972 240.244
R6785 gnd.n3879 gnd.n1780 240.244
R6786 gnd.n4062 gnd.n1780 240.244
R6787 gnd.n4062 gnd.n1776 240.244
R6788 gnd.n4068 gnd.n1776 240.244
R6789 gnd.n4068 gnd.n1768 240.244
R6790 gnd.n4083 gnd.n1768 240.244
R6791 gnd.n4083 gnd.n1764 240.244
R6792 gnd.n4089 gnd.n1764 240.244
R6793 gnd.n4089 gnd.n1756 240.244
R6794 gnd.n4106 gnd.n1756 240.244
R6795 gnd.n4106 gnd.n1752 240.244
R6796 gnd.n4113 gnd.n1752 240.244
R6797 gnd.n4113 gnd.n1442 240.244
R6798 gnd.n4375 gnd.n1442 240.244
R6799 gnd.n4375 gnd.n1443 240.244
R6800 gnd.n4371 gnd.n1443 240.244
R6801 gnd.n4371 gnd.n1449 240.244
R6802 gnd.n4367 gnd.n1449 240.244
R6803 gnd.n4367 gnd.n1452 240.244
R6804 gnd.n4363 gnd.n1452 240.244
R6805 gnd.n4363 gnd.n1458 240.244
R6806 gnd.n1574 gnd.n1458 240.244
R6807 gnd.n1580 gnd.n1574 240.244
R6808 gnd.n1581 gnd.n1580 240.244
R6809 gnd.n4187 gnd.n1581 240.244
R6810 gnd.n4187 gnd.n1569 240.244
R6811 gnd.n4195 gnd.n1569 240.244
R6812 gnd.n4195 gnd.n1570 240.244
R6813 gnd.n1570 gnd.n1547 240.244
R6814 gnd.n4224 gnd.n1547 240.244
R6815 gnd.n4224 gnd.n1542 240.244
R6816 gnd.n4247 gnd.n1542 240.244
R6817 gnd.n4247 gnd.n1543 240.244
R6818 gnd.n4243 gnd.n1543 240.244
R6819 gnd.n4243 gnd.n4242 240.244
R6820 gnd.n4242 gnd.n4241 240.244
R6821 gnd.n4241 gnd.n4232 240.244
R6822 gnd.n4236 gnd.n4232 240.244
R6823 gnd.n4236 gnd.n1522 240.244
R6824 gnd.n4300 gnd.n1522 240.244
R6825 gnd.n4300 gnd.n1519 240.244
R6826 gnd.n4307 gnd.n1519 240.244
R6827 gnd.n4307 gnd.n1520 240.244
R6828 gnd.n1520 gnd.n257 240.244
R6829 gnd.n7092 gnd.n257 240.244
R6830 gnd.n7092 gnd.n258 240.244
R6831 gnd.n7087 gnd.n258 240.244
R6832 gnd.n7087 gnd.n7086 240.244
R6833 gnd.n7086 gnd.n262 240.244
R6834 gnd.n278 gnd.n262 240.244
R6835 gnd.n279 gnd.n278 240.244
R6836 gnd.n279 gnd.n270 240.244
R6837 gnd.n7072 gnd.n270 240.244
R6838 gnd.n7072 gnd.n271 240.244
R6839 gnd.n7068 gnd.n271 240.244
R6840 gnd.n7068 gnd.n7067 240.244
R6841 gnd.n7067 gnd.n7045 240.244
R6842 gnd.n7045 gnd.n287 240.244
R6843 gnd.n7041 gnd.n287 240.244
R6844 gnd.n7041 gnd.n7040 240.244
R6845 gnd.n7040 gnd.n7039 240.244
R6846 gnd.n7039 gnd.n293 240.244
R6847 gnd.n7035 gnd.n293 240.244
R6848 gnd.n7035 gnd.n7034 240.244
R6849 gnd.n7034 gnd.n7032 240.244
R6850 gnd.n7032 gnd.n299 240.244
R6851 gnd.n7028 gnd.n299 240.244
R6852 gnd.n7028 gnd.n302 240.244
R6853 gnd.n7024 gnd.n302 240.244
R6854 gnd.n7024 gnd.n311 240.244
R6855 gnd.n7020 gnd.n311 240.244
R6856 gnd.n7020 gnd.n313 240.244
R6857 gnd.n7016 gnd.n313 240.244
R6858 gnd.n7016 gnd.n319 240.244
R6859 gnd.n7012 gnd.n319 240.244
R6860 gnd.n7012 gnd.n321 240.244
R6861 gnd.n6271 gnd.n762 240.244
R6862 gnd.n6271 gnd.n764 240.244
R6863 gnd.n6267 gnd.n764 240.244
R6864 gnd.n6267 gnd.n770 240.244
R6865 gnd.n6263 gnd.n770 240.244
R6866 gnd.n6263 gnd.n772 240.244
R6867 gnd.n6259 gnd.n772 240.244
R6868 gnd.n6259 gnd.n778 240.244
R6869 gnd.n6255 gnd.n778 240.244
R6870 gnd.n6255 gnd.n780 240.244
R6871 gnd.n6251 gnd.n780 240.244
R6872 gnd.n6251 gnd.n786 240.244
R6873 gnd.n6247 gnd.n786 240.244
R6874 gnd.n6247 gnd.n788 240.244
R6875 gnd.n6243 gnd.n788 240.244
R6876 gnd.n6243 gnd.n794 240.244
R6877 gnd.n6239 gnd.n794 240.244
R6878 gnd.n6239 gnd.n796 240.244
R6879 gnd.n6235 gnd.n796 240.244
R6880 gnd.n6235 gnd.n802 240.244
R6881 gnd.n6231 gnd.n802 240.244
R6882 gnd.n6231 gnd.n804 240.244
R6883 gnd.n6227 gnd.n804 240.244
R6884 gnd.n6227 gnd.n810 240.244
R6885 gnd.n6223 gnd.n810 240.244
R6886 gnd.n6223 gnd.n812 240.244
R6887 gnd.n6219 gnd.n812 240.244
R6888 gnd.n6219 gnd.n818 240.244
R6889 gnd.n6215 gnd.n818 240.244
R6890 gnd.n6215 gnd.n820 240.244
R6891 gnd.n6211 gnd.n820 240.244
R6892 gnd.n6211 gnd.n826 240.244
R6893 gnd.n6207 gnd.n826 240.244
R6894 gnd.n6207 gnd.n828 240.244
R6895 gnd.n6203 gnd.n828 240.244
R6896 gnd.n6203 gnd.n834 240.244
R6897 gnd.n6199 gnd.n834 240.244
R6898 gnd.n6199 gnd.n836 240.244
R6899 gnd.n6195 gnd.n836 240.244
R6900 gnd.n6195 gnd.n842 240.244
R6901 gnd.n6191 gnd.n842 240.244
R6902 gnd.n6191 gnd.n844 240.244
R6903 gnd.n6187 gnd.n844 240.244
R6904 gnd.n6187 gnd.n850 240.244
R6905 gnd.n6183 gnd.n850 240.244
R6906 gnd.n6183 gnd.n852 240.244
R6907 gnd.n6179 gnd.n852 240.244
R6908 gnd.n6179 gnd.n858 240.244
R6909 gnd.n6175 gnd.n858 240.244
R6910 gnd.n6175 gnd.n860 240.244
R6911 gnd.n6171 gnd.n860 240.244
R6912 gnd.n6171 gnd.n866 240.244
R6913 gnd.n6167 gnd.n866 240.244
R6914 gnd.n6167 gnd.n868 240.244
R6915 gnd.n6163 gnd.n868 240.244
R6916 gnd.n6163 gnd.n874 240.244
R6917 gnd.n6159 gnd.n874 240.244
R6918 gnd.n6159 gnd.n876 240.244
R6919 gnd.n6155 gnd.n876 240.244
R6920 gnd.n6155 gnd.n882 240.244
R6921 gnd.n6151 gnd.n882 240.244
R6922 gnd.n6151 gnd.n884 240.244
R6923 gnd.n6147 gnd.n884 240.244
R6924 gnd.n6147 gnd.n890 240.244
R6925 gnd.n6143 gnd.n890 240.244
R6926 gnd.n6143 gnd.n892 240.244
R6927 gnd.n6139 gnd.n892 240.244
R6928 gnd.n6139 gnd.n898 240.244
R6929 gnd.n6135 gnd.n898 240.244
R6930 gnd.n6135 gnd.n900 240.244
R6931 gnd.n6131 gnd.n900 240.244
R6932 gnd.n6131 gnd.n906 240.244
R6933 gnd.n6127 gnd.n906 240.244
R6934 gnd.n6127 gnd.n908 240.244
R6935 gnd.n6123 gnd.n908 240.244
R6936 gnd.n6123 gnd.n914 240.244
R6937 gnd.n6119 gnd.n914 240.244
R6938 gnd.n6119 gnd.n916 240.244
R6939 gnd.n6115 gnd.n916 240.244
R6940 gnd.n6115 gnd.n922 240.244
R6941 gnd.n6111 gnd.n922 240.244
R6942 gnd.n6111 gnd.n924 240.244
R6943 gnd.n6107 gnd.n924 240.244
R6944 gnd.n6107 gnd.n930 240.244
R6945 gnd.n1336 gnd.n1335 240.244
R6946 gnd.n1337 gnd.n1336 240.244
R6947 gnd.n2546 gnd.n1337 240.244
R6948 gnd.n2546 gnd.n1340 240.244
R6949 gnd.n1341 gnd.n1340 240.244
R6950 gnd.n1342 gnd.n1341 240.244
R6951 gnd.n2538 gnd.n1342 240.244
R6952 gnd.n2538 gnd.n1345 240.244
R6953 gnd.n1346 gnd.n1345 240.244
R6954 gnd.n1347 gnd.n1346 240.244
R6955 gnd.n3179 gnd.n1347 240.244
R6956 gnd.n3179 gnd.n1350 240.244
R6957 gnd.n1351 gnd.n1350 240.244
R6958 gnd.n1352 gnd.n1351 240.244
R6959 gnd.n2253 gnd.n1352 240.244
R6960 gnd.n2253 gnd.n1355 240.244
R6961 gnd.n1356 gnd.n1355 240.244
R6962 gnd.n1357 gnd.n1356 240.244
R6963 gnd.n3459 gnd.n1357 240.244
R6964 gnd.n3459 gnd.n1360 240.244
R6965 gnd.n1361 gnd.n1360 240.244
R6966 gnd.n1362 gnd.n1361 240.244
R6967 gnd.n3490 gnd.n1362 240.244
R6968 gnd.n3490 gnd.n1365 240.244
R6969 gnd.n1366 gnd.n1365 240.244
R6970 gnd.n1367 gnd.n1366 240.244
R6971 gnd.n2190 gnd.n1367 240.244
R6972 gnd.n2190 gnd.n1370 240.244
R6973 gnd.n1371 gnd.n1370 240.244
R6974 gnd.n1372 gnd.n1371 240.244
R6975 gnd.n3544 gnd.n1372 240.244
R6976 gnd.n3544 gnd.n1375 240.244
R6977 gnd.n1376 gnd.n1375 240.244
R6978 gnd.n1377 gnd.n1376 240.244
R6979 gnd.n2148 gnd.n1377 240.244
R6980 gnd.n2148 gnd.n1380 240.244
R6981 gnd.n1381 gnd.n1380 240.244
R6982 gnd.n1382 gnd.n1381 240.244
R6983 gnd.n3616 gnd.n1382 240.244
R6984 gnd.n3616 gnd.n1385 240.244
R6985 gnd.n1386 gnd.n1385 240.244
R6986 gnd.n1387 gnd.n1386 240.244
R6987 gnd.n2103 gnd.n1387 240.244
R6988 gnd.n2103 gnd.n1390 240.244
R6989 gnd.n1391 gnd.n1390 240.244
R6990 gnd.n1392 gnd.n1391 240.244
R6991 gnd.n2073 gnd.n1392 240.244
R6992 gnd.n2073 gnd.n1395 240.244
R6993 gnd.n1396 gnd.n1395 240.244
R6994 gnd.n1397 gnd.n1396 240.244
R6995 gnd.n3714 gnd.n1397 240.244
R6996 gnd.n3714 gnd.n1400 240.244
R6997 gnd.n1401 gnd.n1400 240.244
R6998 gnd.n1402 gnd.n1401 240.244
R6999 gnd.n3754 gnd.n1402 240.244
R7000 gnd.n3754 gnd.n1405 240.244
R7001 gnd.n1406 gnd.n1405 240.244
R7002 gnd.n1407 gnd.n1406 240.244
R7003 gnd.n3793 gnd.n1407 240.244
R7004 gnd.n3793 gnd.n1410 240.244
R7005 gnd.n1411 gnd.n1410 240.244
R7006 gnd.n1412 gnd.n1411 240.244
R7007 gnd.n3834 gnd.n1412 240.244
R7008 gnd.n3834 gnd.n1415 240.244
R7009 gnd.n1416 gnd.n1415 240.244
R7010 gnd.n1417 gnd.n1416 240.244
R7011 gnd.n3851 gnd.n1417 240.244
R7012 gnd.n3851 gnd.n1420 240.244
R7013 gnd.n1421 gnd.n1420 240.244
R7014 gnd.n1422 gnd.n1421 240.244
R7015 gnd.n4059 gnd.n1422 240.244
R7016 gnd.n4059 gnd.n1425 240.244
R7017 gnd.n1426 gnd.n1425 240.244
R7018 gnd.n1427 gnd.n1426 240.244
R7019 gnd.n4080 gnd.n1427 240.244
R7020 gnd.n4080 gnd.n1430 240.244
R7021 gnd.n1431 gnd.n1430 240.244
R7022 gnd.n1432 gnd.n1431 240.244
R7023 gnd.n4103 gnd.n1432 240.244
R7024 gnd.n4103 gnd.n1435 240.244
R7025 gnd.n1436 gnd.n1435 240.244
R7026 gnd.n4378 gnd.n1436 240.244
R7027 gnd.n3011 gnd.n3010 240.244
R7028 gnd.n3026 gnd.n3010 240.244
R7029 gnd.n3028 gnd.n3027 240.244
R7030 gnd.n3038 gnd.n3037 240.244
R7031 gnd.n3049 gnd.n3048 240.244
R7032 gnd.n3051 gnd.n3050 240.244
R7033 gnd.n3061 gnd.n3060 240.244
R7034 gnd.n3074 gnd.n3073 240.244
R7035 gnd.n3076 gnd.n3075 240.244
R7036 gnd.n2501 gnd.n2500 240.244
R7037 gnd.n3004 gnd.n2502 240.244
R7038 gnd.n2506 gnd.n2505 240.244
R7039 gnd.n2512 gnd.n2507 240.244
R7040 gnd.n2514 gnd.n2513 240.244
R7041 gnd.n2518 gnd.n2517 240.244
R7042 gnd.n2519 gnd.n2518 240.244
R7043 gnd.n2545 gnd.n2519 240.244
R7044 gnd.n2545 gnd.n2522 240.244
R7045 gnd.n2523 gnd.n2522 240.244
R7046 gnd.n2524 gnd.n2523 240.244
R7047 gnd.n2537 gnd.n2524 240.244
R7048 gnd.n2537 gnd.n2527 240.244
R7049 gnd.n2528 gnd.n2527 240.244
R7050 gnd.n2529 gnd.n2528 240.244
R7051 gnd.n3181 gnd.n2529 240.244
R7052 gnd.n3182 gnd.n3181 240.244
R7053 gnd.n3184 gnd.n3182 240.244
R7054 gnd.n3184 gnd.n2261 240.244
R7055 gnd.n3187 gnd.n2261 240.244
R7056 gnd.n3188 gnd.n3187 240.244
R7057 gnd.n3189 gnd.n3188 240.244
R7058 gnd.n3189 gnd.n2233 240.244
R7059 gnd.n3461 gnd.n2233 240.244
R7060 gnd.n3461 gnd.n2229 240.244
R7061 gnd.n3467 gnd.n2229 240.244
R7062 gnd.n3467 gnd.n2213 240.244
R7063 gnd.n3492 gnd.n2213 240.244
R7064 gnd.n3492 gnd.n2207 240.244
R7065 gnd.n3499 gnd.n2207 240.244
R7066 gnd.n3499 gnd.n2208 240.244
R7067 gnd.n2208 gnd.n2183 240.244
R7068 gnd.n3528 gnd.n2183 240.244
R7069 gnd.n3528 gnd.n2179 240.244
R7070 gnd.n3534 gnd.n2179 240.244
R7071 gnd.n3534 gnd.n2162 240.244
R7072 gnd.n3556 gnd.n2162 240.244
R7073 gnd.n3556 gnd.n2156 240.244
R7074 gnd.n3563 gnd.n2156 240.244
R7075 gnd.n3563 gnd.n2157 240.244
R7076 gnd.n2157 gnd.n2132 240.244
R7077 gnd.n3594 gnd.n2132 240.244
R7078 gnd.n3594 gnd.n2126 240.244
R7079 gnd.n3615 gnd.n2126 240.244
R7080 gnd.n3615 gnd.n2127 240.244
R7081 gnd.n3599 gnd.n2127 240.244
R7082 gnd.n3600 gnd.n3599 240.244
R7083 gnd.n3601 gnd.n3600 240.244
R7084 gnd.n3601 gnd.n2098 240.244
R7085 gnd.n2098 gnd.n2082 240.244
R7086 gnd.n3676 gnd.n2082 240.244
R7087 gnd.n3677 gnd.n3676 240.244
R7088 gnd.n3677 gnd.n2076 240.244
R7089 gnd.n2078 gnd.n2076 240.244
R7090 gnd.n3684 gnd.n2078 240.244
R7091 gnd.n3684 gnd.n2053 240.244
R7092 gnd.n3733 gnd.n2053 240.244
R7093 gnd.n3733 gnd.n2054 240.244
R7094 gnd.n3727 gnd.n2054 240.244
R7095 gnd.n3727 gnd.n2030 240.244
R7096 gnd.n3773 gnd.n2030 240.244
R7097 gnd.n3773 gnd.n2031 240.244
R7098 gnd.n3767 gnd.n2031 240.244
R7099 gnd.n3767 gnd.n2009 240.244
R7100 gnd.n3812 gnd.n2009 240.244
R7101 gnd.n3812 gnd.n2000 240.244
R7102 gnd.n3806 gnd.n2000 240.244
R7103 gnd.n3806 gnd.n1985 240.244
R7104 gnd.n3860 gnd.n1985 240.244
R7105 gnd.n3860 gnd.n1978 240.244
R7106 gnd.n3849 gnd.n1978 240.244
R7107 gnd.n3853 gnd.n3849 240.244
R7108 gnd.n3853 gnd.n1785 240.244
R7109 gnd.n4051 gnd.n1785 240.244
R7110 gnd.n4051 gnd.n1781 240.244
R7111 gnd.n4057 gnd.n1781 240.244
R7112 gnd.n4057 gnd.n1774 240.244
R7113 gnd.n4072 gnd.n1774 240.244
R7114 gnd.n4072 gnd.n1770 240.244
R7115 gnd.n4078 gnd.n1770 240.244
R7116 gnd.n4078 gnd.n1762 240.244
R7117 gnd.n4093 gnd.n1762 240.244
R7118 gnd.n4093 gnd.n1758 240.244
R7119 gnd.n4100 gnd.n1758 240.244
R7120 gnd.n4100 gnd.n1751 240.244
R7121 gnd.n4116 gnd.n1751 240.244
R7122 gnd.n4116 gnd.n1440 240.244
R7123 gnd.n1660 gnd.n1659 240.244
R7124 gnd.n1663 gnd.n1662 240.244
R7125 gnd.n1679 gnd.n1678 240.244
R7126 gnd.n1682 gnd.n1681 240.244
R7127 gnd.n1698 gnd.n1697 240.244
R7128 gnd.n1701 gnd.n1700 240.244
R7129 gnd.n1717 gnd.n1716 240.244
R7130 gnd.n1720 gnd.n1719 240.244
R7131 gnd.n1734 gnd.n1733 240.244
R7132 gnd.n1737 gnd.n1736 240.244
R7133 gnd.n1742 gnd.n1739 240.244
R7134 gnd.n1745 gnd.n1744 240.244
R7135 gnd.n4121 gnd.n1747 240.244
R7136 gnd.n4124 gnd.n4123 240.244
R7137 gnd.n2273 gnd.n2272 240.132
R7138 gnd.n3899 gnd.n3898 240.132
R7139 gnd.n6274 gnd.n758 225.874
R7140 gnd.n6282 gnd.n758 225.874
R7141 gnd.n6283 gnd.n6282 225.874
R7142 gnd.n6284 gnd.n6283 225.874
R7143 gnd.n6284 gnd.n752 225.874
R7144 gnd.n6292 gnd.n752 225.874
R7145 gnd.n6293 gnd.n6292 225.874
R7146 gnd.n6294 gnd.n6293 225.874
R7147 gnd.n6294 gnd.n746 225.874
R7148 gnd.n6302 gnd.n746 225.874
R7149 gnd.n6303 gnd.n6302 225.874
R7150 gnd.n6304 gnd.n6303 225.874
R7151 gnd.n6304 gnd.n740 225.874
R7152 gnd.n6312 gnd.n740 225.874
R7153 gnd.n6313 gnd.n6312 225.874
R7154 gnd.n6314 gnd.n6313 225.874
R7155 gnd.n6314 gnd.n734 225.874
R7156 gnd.n6322 gnd.n734 225.874
R7157 gnd.n6323 gnd.n6322 225.874
R7158 gnd.n6324 gnd.n6323 225.874
R7159 gnd.n6324 gnd.n728 225.874
R7160 gnd.n6332 gnd.n728 225.874
R7161 gnd.n6333 gnd.n6332 225.874
R7162 gnd.n6334 gnd.n6333 225.874
R7163 gnd.n6334 gnd.n722 225.874
R7164 gnd.n6342 gnd.n722 225.874
R7165 gnd.n6343 gnd.n6342 225.874
R7166 gnd.n6344 gnd.n6343 225.874
R7167 gnd.n6344 gnd.n716 225.874
R7168 gnd.n6352 gnd.n716 225.874
R7169 gnd.n6353 gnd.n6352 225.874
R7170 gnd.n6354 gnd.n6353 225.874
R7171 gnd.n6354 gnd.n710 225.874
R7172 gnd.n6362 gnd.n710 225.874
R7173 gnd.n6363 gnd.n6362 225.874
R7174 gnd.n6364 gnd.n6363 225.874
R7175 gnd.n6364 gnd.n704 225.874
R7176 gnd.n6372 gnd.n704 225.874
R7177 gnd.n6373 gnd.n6372 225.874
R7178 gnd.n6374 gnd.n6373 225.874
R7179 gnd.n6374 gnd.n698 225.874
R7180 gnd.n6382 gnd.n698 225.874
R7181 gnd.n6383 gnd.n6382 225.874
R7182 gnd.n6384 gnd.n6383 225.874
R7183 gnd.n6384 gnd.n692 225.874
R7184 gnd.n6392 gnd.n692 225.874
R7185 gnd.n6393 gnd.n6392 225.874
R7186 gnd.n6394 gnd.n6393 225.874
R7187 gnd.n6394 gnd.n686 225.874
R7188 gnd.n6402 gnd.n686 225.874
R7189 gnd.n6403 gnd.n6402 225.874
R7190 gnd.n6404 gnd.n6403 225.874
R7191 gnd.n6404 gnd.n680 225.874
R7192 gnd.n6412 gnd.n680 225.874
R7193 gnd.n6413 gnd.n6412 225.874
R7194 gnd.n6414 gnd.n6413 225.874
R7195 gnd.n6414 gnd.n674 225.874
R7196 gnd.n6422 gnd.n674 225.874
R7197 gnd.n6423 gnd.n6422 225.874
R7198 gnd.n6424 gnd.n6423 225.874
R7199 gnd.n6424 gnd.n668 225.874
R7200 gnd.n6432 gnd.n668 225.874
R7201 gnd.n6433 gnd.n6432 225.874
R7202 gnd.n6434 gnd.n6433 225.874
R7203 gnd.n6434 gnd.n662 225.874
R7204 gnd.n6442 gnd.n662 225.874
R7205 gnd.n6443 gnd.n6442 225.874
R7206 gnd.n6444 gnd.n6443 225.874
R7207 gnd.n6444 gnd.n656 225.874
R7208 gnd.n6452 gnd.n656 225.874
R7209 gnd.n6453 gnd.n6452 225.874
R7210 gnd.n6454 gnd.n6453 225.874
R7211 gnd.n6454 gnd.n650 225.874
R7212 gnd.n6462 gnd.n650 225.874
R7213 gnd.n6463 gnd.n6462 225.874
R7214 gnd.n6464 gnd.n6463 225.874
R7215 gnd.n6464 gnd.n644 225.874
R7216 gnd.n6472 gnd.n644 225.874
R7217 gnd.n6473 gnd.n6472 225.874
R7218 gnd.n6474 gnd.n6473 225.874
R7219 gnd.n6474 gnd.n638 225.874
R7220 gnd.n6482 gnd.n638 225.874
R7221 gnd.n6483 gnd.n6482 225.874
R7222 gnd.n6484 gnd.n6483 225.874
R7223 gnd.n6484 gnd.n632 225.874
R7224 gnd.n6492 gnd.n632 225.874
R7225 gnd.n6493 gnd.n6492 225.874
R7226 gnd.n6494 gnd.n6493 225.874
R7227 gnd.n6494 gnd.n626 225.874
R7228 gnd.n6502 gnd.n626 225.874
R7229 gnd.n6503 gnd.n6502 225.874
R7230 gnd.n6504 gnd.n6503 225.874
R7231 gnd.n6504 gnd.n620 225.874
R7232 gnd.n6512 gnd.n620 225.874
R7233 gnd.n6513 gnd.n6512 225.874
R7234 gnd.n6514 gnd.n6513 225.874
R7235 gnd.n6514 gnd.n614 225.874
R7236 gnd.n6522 gnd.n614 225.874
R7237 gnd.n6523 gnd.n6522 225.874
R7238 gnd.n6524 gnd.n6523 225.874
R7239 gnd.n6524 gnd.n608 225.874
R7240 gnd.n6532 gnd.n608 225.874
R7241 gnd.n6533 gnd.n6532 225.874
R7242 gnd.n6534 gnd.n6533 225.874
R7243 gnd.n6534 gnd.n602 225.874
R7244 gnd.n6542 gnd.n602 225.874
R7245 gnd.n6543 gnd.n6542 225.874
R7246 gnd.n6544 gnd.n6543 225.874
R7247 gnd.n6544 gnd.n596 225.874
R7248 gnd.n6552 gnd.n596 225.874
R7249 gnd.n6553 gnd.n6552 225.874
R7250 gnd.n6554 gnd.n6553 225.874
R7251 gnd.n6554 gnd.n590 225.874
R7252 gnd.n6562 gnd.n590 225.874
R7253 gnd.n6563 gnd.n6562 225.874
R7254 gnd.n6564 gnd.n6563 225.874
R7255 gnd.n6564 gnd.n584 225.874
R7256 gnd.n6572 gnd.n584 225.874
R7257 gnd.n6573 gnd.n6572 225.874
R7258 gnd.n6574 gnd.n6573 225.874
R7259 gnd.n6574 gnd.n578 225.874
R7260 gnd.n6582 gnd.n578 225.874
R7261 gnd.n6583 gnd.n6582 225.874
R7262 gnd.n6584 gnd.n6583 225.874
R7263 gnd.n6584 gnd.n572 225.874
R7264 gnd.n6592 gnd.n572 225.874
R7265 gnd.n6593 gnd.n6592 225.874
R7266 gnd.n6594 gnd.n6593 225.874
R7267 gnd.n6594 gnd.n566 225.874
R7268 gnd.n6602 gnd.n566 225.874
R7269 gnd.n6603 gnd.n6602 225.874
R7270 gnd.n6604 gnd.n6603 225.874
R7271 gnd.n6604 gnd.n560 225.874
R7272 gnd.n6612 gnd.n560 225.874
R7273 gnd.n6613 gnd.n6612 225.874
R7274 gnd.n6614 gnd.n6613 225.874
R7275 gnd.n6614 gnd.n554 225.874
R7276 gnd.n6622 gnd.n554 225.874
R7277 gnd.n6623 gnd.n6622 225.874
R7278 gnd.n6624 gnd.n6623 225.874
R7279 gnd.n6624 gnd.n548 225.874
R7280 gnd.n6632 gnd.n548 225.874
R7281 gnd.n6633 gnd.n6632 225.874
R7282 gnd.n6634 gnd.n6633 225.874
R7283 gnd.n6634 gnd.n542 225.874
R7284 gnd.n6642 gnd.n542 225.874
R7285 gnd.n6643 gnd.n6642 225.874
R7286 gnd.n6644 gnd.n6643 225.874
R7287 gnd.n6644 gnd.n536 225.874
R7288 gnd.n6652 gnd.n536 225.874
R7289 gnd.n6653 gnd.n6652 225.874
R7290 gnd.n6654 gnd.n6653 225.874
R7291 gnd.n6654 gnd.n530 225.874
R7292 gnd.n6662 gnd.n530 225.874
R7293 gnd.n6663 gnd.n6662 225.874
R7294 gnd.n6664 gnd.n6663 225.874
R7295 gnd.n6664 gnd.n524 225.874
R7296 gnd.n6672 gnd.n524 225.874
R7297 gnd.n6673 gnd.n6672 225.874
R7298 gnd.n6674 gnd.n6673 225.874
R7299 gnd.n6674 gnd.n518 225.874
R7300 gnd.n6682 gnd.n518 225.874
R7301 gnd.n6683 gnd.n6682 225.874
R7302 gnd.n6684 gnd.n6683 225.874
R7303 gnd.n6684 gnd.n512 225.874
R7304 gnd.n6692 gnd.n512 225.874
R7305 gnd.n6693 gnd.n6692 225.874
R7306 gnd.n6694 gnd.n6693 225.874
R7307 gnd.n6694 gnd.n506 225.874
R7308 gnd.n6702 gnd.n506 225.874
R7309 gnd.n6703 gnd.n6702 225.874
R7310 gnd.n6704 gnd.n6703 225.874
R7311 gnd.n6704 gnd.n500 225.874
R7312 gnd.n6712 gnd.n500 225.874
R7313 gnd.n6713 gnd.n6712 225.874
R7314 gnd.n6714 gnd.n6713 225.874
R7315 gnd.n6714 gnd.n494 225.874
R7316 gnd.n6722 gnd.n494 225.874
R7317 gnd.n6723 gnd.n6722 225.874
R7318 gnd.n6724 gnd.n6723 225.874
R7319 gnd.n6724 gnd.n488 225.874
R7320 gnd.n6732 gnd.n488 225.874
R7321 gnd.n6733 gnd.n6732 225.874
R7322 gnd.n6734 gnd.n6733 225.874
R7323 gnd.n6734 gnd.n482 225.874
R7324 gnd.n6742 gnd.n482 225.874
R7325 gnd.n6743 gnd.n6742 225.874
R7326 gnd.n6744 gnd.n6743 225.874
R7327 gnd.n6744 gnd.n476 225.874
R7328 gnd.n6752 gnd.n476 225.874
R7329 gnd.n6753 gnd.n6752 225.874
R7330 gnd.n6754 gnd.n6753 225.874
R7331 gnd.n6754 gnd.n470 225.874
R7332 gnd.n6762 gnd.n470 225.874
R7333 gnd.n6763 gnd.n6762 225.874
R7334 gnd.n6764 gnd.n6763 225.874
R7335 gnd.n6764 gnd.n464 225.874
R7336 gnd.n6772 gnd.n464 225.874
R7337 gnd.n6773 gnd.n6772 225.874
R7338 gnd.n6774 gnd.n6773 225.874
R7339 gnd.n6774 gnd.n458 225.874
R7340 gnd.n6782 gnd.n458 225.874
R7341 gnd.n6783 gnd.n6782 225.874
R7342 gnd.n6784 gnd.n6783 225.874
R7343 gnd.n6784 gnd.n452 225.874
R7344 gnd.n6793 gnd.n452 225.874
R7345 gnd.n6794 gnd.n6793 225.874
R7346 gnd.n5212 gnd.t125 224.174
R7347 gnd.n4815 gnd.t37 224.174
R7348 gnd.n1826 gnd.n1823 199.319
R7349 gnd.n1954 gnd.n1823 199.319
R7350 gnd.n2406 gnd.n2400 199.319
R7351 gnd.n2405 gnd.n2400 199.319
R7352 gnd.n2274 gnd.n2271 186.49
R7353 gnd.n3900 gnd.n3897 186.49
R7354 gnd.n5917 gnd.n5916 185
R7355 gnd.n5915 gnd.n5914 185
R7356 gnd.n5894 gnd.n5893 185
R7357 gnd.n5909 gnd.n5908 185
R7358 gnd.n5907 gnd.n5906 185
R7359 gnd.n5898 gnd.n5897 185
R7360 gnd.n5901 gnd.n5900 185
R7361 gnd.n5885 gnd.n5884 185
R7362 gnd.n5883 gnd.n5882 185
R7363 gnd.n5862 gnd.n5861 185
R7364 gnd.n5877 gnd.n5876 185
R7365 gnd.n5875 gnd.n5874 185
R7366 gnd.n5866 gnd.n5865 185
R7367 gnd.n5869 gnd.n5868 185
R7368 gnd.n5853 gnd.n5852 185
R7369 gnd.n5851 gnd.n5850 185
R7370 gnd.n5830 gnd.n5829 185
R7371 gnd.n5845 gnd.n5844 185
R7372 gnd.n5843 gnd.n5842 185
R7373 gnd.n5834 gnd.n5833 185
R7374 gnd.n5837 gnd.n5836 185
R7375 gnd.n5822 gnd.n5821 185
R7376 gnd.n5820 gnd.n5819 185
R7377 gnd.n5799 gnd.n5798 185
R7378 gnd.n5814 gnd.n5813 185
R7379 gnd.n5812 gnd.n5811 185
R7380 gnd.n5803 gnd.n5802 185
R7381 gnd.n5806 gnd.n5805 185
R7382 gnd.n5790 gnd.n5789 185
R7383 gnd.n5788 gnd.n5787 185
R7384 gnd.n5767 gnd.n5766 185
R7385 gnd.n5782 gnd.n5781 185
R7386 gnd.n5780 gnd.n5779 185
R7387 gnd.n5771 gnd.n5770 185
R7388 gnd.n5774 gnd.n5773 185
R7389 gnd.n5758 gnd.n5757 185
R7390 gnd.n5756 gnd.n5755 185
R7391 gnd.n5735 gnd.n5734 185
R7392 gnd.n5750 gnd.n5749 185
R7393 gnd.n5748 gnd.n5747 185
R7394 gnd.n5739 gnd.n5738 185
R7395 gnd.n5742 gnd.n5741 185
R7396 gnd.n5726 gnd.n5725 185
R7397 gnd.n5724 gnd.n5723 185
R7398 gnd.n5703 gnd.n5702 185
R7399 gnd.n5718 gnd.n5717 185
R7400 gnd.n5716 gnd.n5715 185
R7401 gnd.n5707 gnd.n5706 185
R7402 gnd.n5710 gnd.n5709 185
R7403 gnd.n5695 gnd.n5694 185
R7404 gnd.n5693 gnd.n5692 185
R7405 gnd.n5672 gnd.n5671 185
R7406 gnd.n5687 gnd.n5686 185
R7407 gnd.n5685 gnd.n5684 185
R7408 gnd.n5676 gnd.n5675 185
R7409 gnd.n5679 gnd.n5678 185
R7410 gnd.n5213 gnd.t124 178.987
R7411 gnd.n4816 gnd.t38 178.987
R7412 gnd.n1 gnd.t273 170.774
R7413 gnd.n7 gnd.t172 170.103
R7414 gnd.n6 gnd.t275 170.103
R7415 gnd.n5 gnd.t281 170.103
R7416 gnd.n4 gnd.t279 170.103
R7417 gnd.n3 gnd.t160 170.103
R7418 gnd.n2 gnd.t144 170.103
R7419 gnd.n1 gnd.t141 170.103
R7420 gnd.n3971 gnd.n3970 163.367
R7421 gnd.n3967 gnd.n3966 163.367
R7422 gnd.n3963 gnd.n3962 163.367
R7423 gnd.n3959 gnd.n3958 163.367
R7424 gnd.n3955 gnd.n3954 163.367
R7425 gnd.n3951 gnd.n3950 163.367
R7426 gnd.n3947 gnd.n3946 163.367
R7427 gnd.n3943 gnd.n3942 163.367
R7428 gnd.n3939 gnd.n3938 163.367
R7429 gnd.n3935 gnd.n3934 163.367
R7430 gnd.n3931 gnd.n3930 163.367
R7431 gnd.n3927 gnd.n3926 163.367
R7432 gnd.n3923 gnd.n3922 163.367
R7433 gnd.n3919 gnd.n3918 163.367
R7434 gnd.n3914 gnd.n3913 163.367
R7435 gnd.n3910 gnd.n3909 163.367
R7436 gnd.n4047 gnd.n4046 163.367
R7437 gnd.n4043 gnd.n4042 163.367
R7438 gnd.n4038 gnd.n4037 163.367
R7439 gnd.n4034 gnd.n4033 163.367
R7440 gnd.n4030 gnd.n4029 163.367
R7441 gnd.n4026 gnd.n4025 163.367
R7442 gnd.n4022 gnd.n4021 163.367
R7443 gnd.n4018 gnd.n4017 163.367
R7444 gnd.n4014 gnd.n4013 163.367
R7445 gnd.n4010 gnd.n4009 163.367
R7446 gnd.n4006 gnd.n4005 163.367
R7447 gnd.n4002 gnd.n4001 163.367
R7448 gnd.n3998 gnd.n3997 163.367
R7449 gnd.n3994 gnd.n3993 163.367
R7450 gnd.n3990 gnd.n3989 163.367
R7451 gnd.n3986 gnd.n3985 163.367
R7452 gnd.n2331 gnd.n2262 163.367
R7453 gnd.n2262 gnd.n2252 163.367
R7454 gnd.n3368 gnd.n2252 163.367
R7455 gnd.n3368 gnd.n2250 163.367
R7456 gnd.n3437 gnd.n2250 163.367
R7457 gnd.n3437 gnd.n2243 163.367
R7458 gnd.n3433 gnd.n2243 163.367
R7459 gnd.n3433 gnd.n3430 163.367
R7460 gnd.n3430 gnd.n3429 163.367
R7461 gnd.n3429 gnd.n2227 163.367
R7462 gnd.n2228 gnd.n2227 163.367
R7463 gnd.n2228 gnd.n2221 163.367
R7464 gnd.n3423 gnd.n2221 163.367
R7465 gnd.n3423 gnd.n3420 163.367
R7466 gnd.n3420 gnd.n3419 163.367
R7467 gnd.n3419 gnd.n2206 163.367
R7468 gnd.n3415 gnd.n2206 163.367
R7469 gnd.n3415 gnd.n2200 163.367
R7470 gnd.n3412 gnd.n2200 163.367
R7471 gnd.n3412 gnd.n2192 163.367
R7472 gnd.n3408 gnd.n2192 163.367
R7473 gnd.n3408 gnd.n2185 163.367
R7474 gnd.n3405 gnd.n2185 163.367
R7475 gnd.n3405 gnd.n2178 163.367
R7476 gnd.n3400 gnd.n2178 163.367
R7477 gnd.n3400 gnd.n2171 163.367
R7478 gnd.n3397 gnd.n2171 163.367
R7479 gnd.n3397 gnd.n2164 163.367
R7480 gnd.n2164 gnd.n2154 163.367
R7481 gnd.n2155 gnd.n2154 163.367
R7482 gnd.n2155 gnd.n2147 163.367
R7483 gnd.n3391 gnd.n2147 163.367
R7484 gnd.n3391 gnd.n2140 163.367
R7485 gnd.n3387 gnd.n2140 163.367
R7486 gnd.n3387 gnd.n2134 163.367
R7487 gnd.n3384 gnd.n2134 163.367
R7488 gnd.n3384 gnd.n2125 163.367
R7489 gnd.n3379 gnd.n2125 163.367
R7490 gnd.n3379 gnd.n2119 163.367
R7491 gnd.n3376 gnd.n2119 163.367
R7492 gnd.n3376 gnd.n2110 163.367
R7493 gnd.n2110 gnd.n2101 163.367
R7494 gnd.n3642 gnd.n2101 163.367
R7495 gnd.n3642 gnd.n2099 163.367
R7496 gnd.n3652 gnd.n2099 163.367
R7497 gnd.n3652 gnd.n2089 163.367
R7498 gnd.n2090 gnd.n2089 163.367
R7499 gnd.n2090 gnd.n2083 163.367
R7500 gnd.n3646 gnd.n2083 163.367
R7501 gnd.n3646 gnd.n2075 163.367
R7502 gnd.n3691 gnd.n2075 163.367
R7503 gnd.n3691 gnd.n2067 163.367
R7504 gnd.n3687 gnd.n2067 163.367
R7505 gnd.n3687 gnd.n2060 163.367
R7506 gnd.n3717 gnd.n2060 163.367
R7507 gnd.n3717 gnd.n2052 163.367
R7508 gnd.n3720 gnd.n2052 163.367
R7509 gnd.n3720 gnd.n2045 163.367
R7510 gnd.n3724 gnd.n2045 163.367
R7511 gnd.n3724 gnd.n2037 163.367
R7512 gnd.n3757 gnd.n2037 163.367
R7513 gnd.n3757 gnd.n2029 163.367
R7514 gnd.n3760 gnd.n2029 163.367
R7515 gnd.n3760 gnd.n2022 163.367
R7516 gnd.n3764 gnd.n2022 163.367
R7517 gnd.n3764 gnd.n2014 163.367
R7518 gnd.n3796 gnd.n2014 163.367
R7519 gnd.n3796 gnd.n2008 163.367
R7520 gnd.n3799 gnd.n2008 163.367
R7521 gnd.n3799 gnd.n2001 163.367
R7522 gnd.n3803 gnd.n2001 163.367
R7523 gnd.n3803 gnd.n1992 163.367
R7524 gnd.n3837 gnd.n1992 163.367
R7525 gnd.n3837 gnd.n1984 163.367
R7526 gnd.n3840 gnd.n1984 163.367
R7527 gnd.n3840 gnd.n1979 163.367
R7528 gnd.n3846 gnd.n1979 163.367
R7529 gnd.n3846 gnd.n1970 163.367
R7530 gnd.n1970 gnd.n1962 163.367
R7531 gnd.n3980 gnd.n1962 163.367
R7532 gnd.n3981 gnd.n3980 163.367
R7533 gnd.n3347 gnd.n2288 163.367
R7534 gnd.n3347 gnd.n2323 163.367
R7535 gnd.n3343 gnd.n3342 163.367
R7536 gnd.n3339 gnd.n3338 163.367
R7537 gnd.n3335 gnd.n3334 163.367
R7538 gnd.n3331 gnd.n3330 163.367
R7539 gnd.n3327 gnd.n3326 163.367
R7540 gnd.n3323 gnd.n3322 163.367
R7541 gnd.n3319 gnd.n3318 163.367
R7542 gnd.n3315 gnd.n3314 163.367
R7543 gnd.n3311 gnd.n3310 163.367
R7544 gnd.n3307 gnd.n3306 163.367
R7545 gnd.n3303 gnd.n3302 163.367
R7546 gnd.n3299 gnd.n3298 163.367
R7547 gnd.n3295 gnd.n3294 163.367
R7548 gnd.n3291 gnd.n3290 163.367
R7549 gnd.n3287 gnd.n3286 163.367
R7550 gnd.n2393 gnd.n2392 163.367
R7551 gnd.n2388 gnd.n2387 163.367
R7552 gnd.n2384 gnd.n2383 163.367
R7553 gnd.n2380 gnd.n2379 163.367
R7554 gnd.n2376 gnd.n2375 163.367
R7555 gnd.n2372 gnd.n2371 163.367
R7556 gnd.n2368 gnd.n2367 163.367
R7557 gnd.n2364 gnd.n2363 163.367
R7558 gnd.n2360 gnd.n2359 163.367
R7559 gnd.n2356 gnd.n2355 163.367
R7560 gnd.n2352 gnd.n2351 163.367
R7561 gnd.n2348 gnd.n2347 163.367
R7562 gnd.n2344 gnd.n2343 163.367
R7563 gnd.n2340 gnd.n2339 163.367
R7564 gnd.n2336 gnd.n2335 163.367
R7565 gnd.n3356 gnd.n2264 163.367
R7566 gnd.n3356 gnd.n2266 163.367
R7567 gnd.n2266 gnd.n2248 163.367
R7568 gnd.n3441 gnd.n2248 163.367
R7569 gnd.n3441 gnd.n2245 163.367
R7570 gnd.n3448 gnd.n2245 163.367
R7571 gnd.n3448 gnd.n2246 163.367
R7572 gnd.n3444 gnd.n2246 163.367
R7573 gnd.n3444 gnd.n2226 163.367
R7574 gnd.n3472 gnd.n2226 163.367
R7575 gnd.n3472 gnd.n2223 163.367
R7576 gnd.n3479 gnd.n2223 163.367
R7577 gnd.n3479 gnd.n2224 163.367
R7578 gnd.n3475 gnd.n2224 163.367
R7579 gnd.n3475 gnd.n2204 163.367
R7580 gnd.n3503 gnd.n2204 163.367
R7581 gnd.n3503 gnd.n2202 163.367
R7582 gnd.n3507 gnd.n2202 163.367
R7583 gnd.n3507 gnd.n2189 163.367
R7584 gnd.n3521 gnd.n2189 163.367
R7585 gnd.n3521 gnd.n2187 163.367
R7586 gnd.n3525 gnd.n2187 163.367
R7587 gnd.n3525 gnd.n2176 163.367
R7588 gnd.n3537 gnd.n2176 163.367
R7589 gnd.n3537 gnd.n2173 163.367
R7590 gnd.n3542 gnd.n2173 163.367
R7591 gnd.n3542 gnd.n2174 163.367
R7592 gnd.n2174 gnd.n2152 163.367
R7593 gnd.n3568 gnd.n2152 163.367
R7594 gnd.n3568 gnd.n2150 163.367
R7595 gnd.n3572 gnd.n2150 163.367
R7596 gnd.n3572 gnd.n2138 163.367
R7597 gnd.n3587 gnd.n2138 163.367
R7598 gnd.n3587 gnd.n2136 163.367
R7599 gnd.n3591 gnd.n2136 163.367
R7600 gnd.n3591 gnd.n2123 163.367
R7601 gnd.n3619 gnd.n2123 163.367
R7602 gnd.n3619 gnd.n2121 163.367
R7603 gnd.n3623 gnd.n2121 163.367
R7604 gnd.n3623 gnd.n2108 163.367
R7605 gnd.n3635 gnd.n2108 163.367
R7606 gnd.n3635 gnd.n2105 163.367
R7607 gnd.n3640 gnd.n2105 163.367
R7608 gnd.n3640 gnd.n2106 163.367
R7609 gnd.n2106 gnd.n2087 163.367
R7610 gnd.n3669 gnd.n2087 163.367
R7611 gnd.n3669 gnd.n2085 163.367
R7612 gnd.n3673 gnd.n2085 163.367
R7613 gnd.n3673 gnd.n2072 163.367
R7614 gnd.n3696 gnd.n2072 163.367
R7615 gnd.n3696 gnd.n2069 163.367
R7616 gnd.n3703 gnd.n2069 163.367
R7617 gnd.n3703 gnd.n2070 163.367
R7618 gnd.n3699 gnd.n2070 163.367
R7619 gnd.n3699 gnd.n2050 163.367
R7620 gnd.n3736 gnd.n2050 163.367
R7621 gnd.n3736 gnd.n2047 163.367
R7622 gnd.n3743 gnd.n2047 163.367
R7623 gnd.n3743 gnd.n2048 163.367
R7624 gnd.n3739 gnd.n2048 163.367
R7625 gnd.n3739 gnd.n2027 163.367
R7626 gnd.n3775 gnd.n2027 163.367
R7627 gnd.n3775 gnd.n2024 163.367
R7628 gnd.n3782 gnd.n2024 163.367
R7629 gnd.n3782 gnd.n2025 163.367
R7630 gnd.n3778 gnd.n2025 163.367
R7631 gnd.n3778 gnd.n2006 163.367
R7632 gnd.n3815 gnd.n2006 163.367
R7633 gnd.n3815 gnd.n2003 163.367
R7634 gnd.n3822 gnd.n2003 163.367
R7635 gnd.n3822 gnd.n2004 163.367
R7636 gnd.n3818 gnd.n2004 163.367
R7637 gnd.n3818 gnd.n1982 163.367
R7638 gnd.n3863 gnd.n1982 163.367
R7639 gnd.n3863 gnd.n1980 163.367
R7640 gnd.n3867 gnd.n1980 163.367
R7641 gnd.n3867 gnd.n1969 163.367
R7642 gnd.n3885 gnd.n1969 163.367
R7643 gnd.n3885 gnd.n1966 163.367
R7644 gnd.n3978 gnd.n1966 163.367
R7645 gnd.n3978 gnd.n1967 163.367
R7646 gnd.n3906 gnd.n3905 156.462
R7647 gnd.n5857 gnd.n5825 153.042
R7648 gnd.n5921 gnd.n5920 152.079
R7649 gnd.n5889 gnd.n5888 152.079
R7650 gnd.n5857 gnd.n5856 152.079
R7651 gnd.n2279 gnd.n2278 152
R7652 gnd.n2280 gnd.n2269 152
R7653 gnd.n2282 gnd.n2281 152
R7654 gnd.n2284 gnd.n2267 152
R7655 gnd.n2286 gnd.n2285 152
R7656 gnd.n3904 gnd.n3888 152
R7657 gnd.n3896 gnd.n3889 152
R7658 gnd.n3895 gnd.n3894 152
R7659 gnd.n3893 gnd.n3890 152
R7660 gnd.n3891 gnd.t77 150.546
R7661 gnd.t166 gnd.n5899 147.661
R7662 gnd.t1 gnd.n5867 147.661
R7663 gnd.t146 gnd.n5835 147.661
R7664 gnd.t164 gnd.n5804 147.661
R7665 gnd.t24 gnd.n5772 147.661
R7666 gnd.t158 gnd.n5740 147.661
R7667 gnd.t168 gnd.n5708 147.661
R7668 gnd.t170 gnd.n5677 147.661
R7669 gnd.n1821 gnd.n1803 143.351
R7670 gnd.n3285 gnd.n2304 143.351
R7671 gnd.n3285 gnd.n2305 143.351
R7672 gnd.n2276 gnd.t126 130.484
R7673 gnd.n2285 gnd.t42 126.766
R7674 gnd.n2283 gnd.t103 126.766
R7675 gnd.n2269 gnd.t53 126.766
R7676 gnd.n2277 gnd.t80 126.766
R7677 gnd.n3892 gnd.t129 126.766
R7678 gnd.n3894 gnd.t100 126.766
R7679 gnd.n3903 gnd.t39 126.766
R7680 gnd.n3905 gnd.t112 126.766
R7681 gnd.n1958 gnd.n1957 108.609
R7682 gnd.n3288 gnd.n3284 108.609
R7683 gnd.n5916 gnd.n5915 104.615
R7684 gnd.n5915 gnd.n5893 104.615
R7685 gnd.n5908 gnd.n5893 104.615
R7686 gnd.n5908 gnd.n5907 104.615
R7687 gnd.n5907 gnd.n5897 104.615
R7688 gnd.n5900 gnd.n5897 104.615
R7689 gnd.n5884 gnd.n5883 104.615
R7690 gnd.n5883 gnd.n5861 104.615
R7691 gnd.n5876 gnd.n5861 104.615
R7692 gnd.n5876 gnd.n5875 104.615
R7693 gnd.n5875 gnd.n5865 104.615
R7694 gnd.n5868 gnd.n5865 104.615
R7695 gnd.n5852 gnd.n5851 104.615
R7696 gnd.n5851 gnd.n5829 104.615
R7697 gnd.n5844 gnd.n5829 104.615
R7698 gnd.n5844 gnd.n5843 104.615
R7699 gnd.n5843 gnd.n5833 104.615
R7700 gnd.n5836 gnd.n5833 104.615
R7701 gnd.n5821 gnd.n5820 104.615
R7702 gnd.n5820 gnd.n5798 104.615
R7703 gnd.n5813 gnd.n5798 104.615
R7704 gnd.n5813 gnd.n5812 104.615
R7705 gnd.n5812 gnd.n5802 104.615
R7706 gnd.n5805 gnd.n5802 104.615
R7707 gnd.n5789 gnd.n5788 104.615
R7708 gnd.n5788 gnd.n5766 104.615
R7709 gnd.n5781 gnd.n5766 104.615
R7710 gnd.n5781 gnd.n5780 104.615
R7711 gnd.n5780 gnd.n5770 104.615
R7712 gnd.n5773 gnd.n5770 104.615
R7713 gnd.n5757 gnd.n5756 104.615
R7714 gnd.n5756 gnd.n5734 104.615
R7715 gnd.n5749 gnd.n5734 104.615
R7716 gnd.n5749 gnd.n5748 104.615
R7717 gnd.n5748 gnd.n5738 104.615
R7718 gnd.n5741 gnd.n5738 104.615
R7719 gnd.n5725 gnd.n5724 104.615
R7720 gnd.n5724 gnd.n5702 104.615
R7721 gnd.n5717 gnd.n5702 104.615
R7722 gnd.n5717 gnd.n5716 104.615
R7723 gnd.n5716 gnd.n5706 104.615
R7724 gnd.n5709 gnd.n5706 104.615
R7725 gnd.n5694 gnd.n5693 104.615
R7726 gnd.n5693 gnd.n5671 104.615
R7727 gnd.n5686 gnd.n5671 104.615
R7728 gnd.n5686 gnd.n5685 104.615
R7729 gnd.n5685 gnd.n5675 104.615
R7730 gnd.n5678 gnd.n5675 104.615
R7731 gnd.n5138 gnd.t52 100.632
R7732 gnd.n4771 gnd.t91 100.632
R7733 gnd.n7318 gnd.n93 99.6594
R7734 gnd.n7316 gnd.n7315 99.6594
R7735 gnd.n7311 gnd.n101 99.6594
R7736 gnd.n7309 gnd.n7308 99.6594
R7737 gnd.n7304 gnd.n108 99.6594
R7738 gnd.n7302 gnd.n7301 99.6594
R7739 gnd.n7297 gnd.n115 99.6594
R7740 gnd.n7295 gnd.n7294 99.6594
R7741 gnd.n7287 gnd.n122 99.6594
R7742 gnd.n7285 gnd.n7284 99.6594
R7743 gnd.n7280 gnd.n129 99.6594
R7744 gnd.n7278 gnd.n7277 99.6594
R7745 gnd.n7273 gnd.n136 99.6594
R7746 gnd.n7271 gnd.n7270 99.6594
R7747 gnd.n7266 gnd.n143 99.6594
R7748 gnd.n7264 gnd.n7263 99.6594
R7749 gnd.n7259 gnd.n150 99.6594
R7750 gnd.n7257 gnd.n7256 99.6594
R7751 gnd.n155 gnd.n154 99.6594
R7752 gnd.n1841 gnd.n1464 99.6594
R7753 gnd.n1849 gnd.n1848 99.6594
R7754 gnd.n1852 gnd.n1851 99.6594
R7755 gnd.n1859 gnd.n1858 99.6594
R7756 gnd.n1862 gnd.n1861 99.6594
R7757 gnd.n1870 gnd.n1869 99.6594
R7758 gnd.n1873 gnd.n1872 99.6594
R7759 gnd.n1827 gnd.n1826 99.6594
R7760 gnd.n1953 gnd.n1952 99.6594
R7761 gnd.n1946 gnd.n1883 99.6594
R7762 gnd.n1945 gnd.n1944 99.6594
R7763 gnd.n1938 gnd.n1889 99.6594
R7764 gnd.n1937 gnd.n1936 99.6594
R7765 gnd.n1930 gnd.n1895 99.6594
R7766 gnd.n1929 gnd.n1928 99.6594
R7767 gnd.n1922 gnd.n1901 99.6594
R7768 gnd.n1921 gnd.n1920 99.6594
R7769 gnd.n1912 gnd.n1907 99.6594
R7770 gnd.n2458 gnd.n2457 99.6594
R7771 gnd.n2453 gnd.n2412 99.6594
R7772 gnd.n2449 gnd.n2411 99.6594
R7773 gnd.n2445 gnd.n2410 99.6594
R7774 gnd.n2441 gnd.n2409 99.6594
R7775 gnd.n2437 gnd.n2408 99.6594
R7776 gnd.n2433 gnd.n2407 99.6594
R7777 gnd.n2405 gnd.n2404 99.6594
R7778 gnd.n3278 gnd.n3277 99.6594
R7779 gnd.n3275 gnd.n3274 99.6594
R7780 gnd.n3270 gnd.n2467 99.6594
R7781 gnd.n3268 gnd.n3267 99.6594
R7782 gnd.n3263 gnd.n2474 99.6594
R7783 gnd.n3261 gnd.n3260 99.6594
R7784 gnd.n3256 gnd.n2481 99.6594
R7785 gnd.n3254 gnd.n3253 99.6594
R7786 gnd.n3249 gnd.n2490 99.6594
R7787 gnd.n3247 gnd.n3246 99.6594
R7788 gnd.n4714 gnd.n4713 99.6594
R7789 gnd.n4708 gnd.n1041 99.6594
R7790 gnd.n4705 gnd.n1042 99.6594
R7791 gnd.n4701 gnd.n1043 99.6594
R7792 gnd.n4697 gnd.n1044 99.6594
R7793 gnd.n4693 gnd.n1045 99.6594
R7794 gnd.n4689 gnd.n1046 99.6594
R7795 gnd.n4685 gnd.n1047 99.6594
R7796 gnd.n4681 gnd.n1048 99.6594
R7797 gnd.n4676 gnd.n1049 99.6594
R7798 gnd.n4672 gnd.n1050 99.6594
R7799 gnd.n4668 gnd.n1051 99.6594
R7800 gnd.n4664 gnd.n1052 99.6594
R7801 gnd.n4660 gnd.n1053 99.6594
R7802 gnd.n4656 gnd.n1054 99.6594
R7803 gnd.n4652 gnd.n1055 99.6594
R7804 gnd.n4648 gnd.n1056 99.6594
R7805 gnd.n4644 gnd.n1057 99.6594
R7806 gnd.n1112 gnd.n1058 99.6594
R7807 gnd.n6047 gnd.n4751 99.6594
R7808 gnd.n6045 gnd.n6044 99.6594
R7809 gnd.n6040 gnd.n4758 99.6594
R7810 gnd.n6038 gnd.n6037 99.6594
R7811 gnd.n6033 gnd.n4765 99.6594
R7812 gnd.n6031 gnd.n6030 99.6594
R7813 gnd.n6026 gnd.n4774 99.6594
R7814 gnd.n6024 gnd.n6023 99.6594
R7815 gnd.n5350 gnd.n5081 99.6594
R7816 gnd.n5107 gnd.n5088 99.6594
R7817 gnd.n5109 gnd.n5089 99.6594
R7818 gnd.n5117 gnd.n5090 99.6594
R7819 gnd.n5119 gnd.n5091 99.6594
R7820 gnd.n5127 gnd.n5092 99.6594
R7821 gnd.n5129 gnd.n5093 99.6594
R7822 gnd.n5137 gnd.n5094 99.6594
R7823 gnd.n6015 gnd.n4781 99.6594
R7824 gnd.n6013 gnd.n6012 99.6594
R7825 gnd.n6008 gnd.n4788 99.6594
R7826 gnd.n6006 gnd.n6005 99.6594
R7827 gnd.n6001 gnd.n4795 99.6594
R7828 gnd.n5999 gnd.n5998 99.6594
R7829 gnd.n5994 gnd.n4802 99.6594
R7830 gnd.n5992 gnd.n5991 99.6594
R7831 gnd.n5987 gnd.n4809 99.6594
R7832 gnd.n5985 gnd.n5984 99.6594
R7833 gnd.n5980 gnd.n4818 99.6594
R7834 gnd.n5978 gnd.n5977 99.6594
R7835 gnd.n5973 gnd.n5972 99.6594
R7836 gnd.n5265 gnd.n5264 99.6594
R7837 gnd.n5259 gnd.n5176 99.6594
R7838 gnd.n5256 gnd.n5177 99.6594
R7839 gnd.n5252 gnd.n5178 99.6594
R7840 gnd.n5248 gnd.n5179 99.6594
R7841 gnd.n5244 gnd.n5180 99.6594
R7842 gnd.n5240 gnd.n5181 99.6594
R7843 gnd.n5236 gnd.n5182 99.6594
R7844 gnd.n5232 gnd.n5183 99.6594
R7845 gnd.n5228 gnd.n5184 99.6594
R7846 gnd.n5224 gnd.n5185 99.6594
R7847 gnd.n5220 gnd.n5186 99.6594
R7848 gnd.n5267 gnd.n5175 99.6594
R7849 gnd.n7181 gnd.n7180 99.6594
R7850 gnd.n7186 gnd.n7185 99.6594
R7851 gnd.n7189 gnd.n7188 99.6594
R7852 gnd.n7194 gnd.n7193 99.6594
R7853 gnd.n7197 gnd.n7196 99.6594
R7854 gnd.n7202 gnd.n7201 99.6594
R7855 gnd.n7205 gnd.n7204 99.6594
R7856 gnd.n7210 gnd.n7209 99.6594
R7857 gnd.n7213 gnd.n80 99.6594
R7858 gnd.n1650 gnd.n1649 99.6594
R7859 gnd.n1653 gnd.n1652 99.6594
R7860 gnd.n1669 gnd.n1668 99.6594
R7861 gnd.n1672 gnd.n1671 99.6594
R7862 gnd.n1688 gnd.n1687 99.6594
R7863 gnd.n1691 gnd.n1690 99.6594
R7864 gnd.n1707 gnd.n1706 99.6594
R7865 gnd.n1710 gnd.n1709 99.6594
R7866 gnd.n1726 gnd.n1725 99.6594
R7867 gnd.n3020 gnd.n3019 99.6594
R7868 gnd.n3023 gnd.n3022 99.6594
R7869 gnd.n3033 gnd.n3032 99.6594
R7870 gnd.n3042 gnd.n3041 99.6594
R7871 gnd.n3045 gnd.n3044 99.6594
R7872 gnd.n3056 gnd.n3055 99.6594
R7873 gnd.n3065 gnd.n3064 99.6594
R7874 gnd.n3068 gnd.n3067 99.6594
R7875 gnd.n3079 gnd.n3078 99.6594
R7876 gnd.n1122 gnd.n1059 99.6594
R7877 gnd.n2689 gnd.n1060 99.6594
R7878 gnd.n2695 gnd.n1061 99.6594
R7879 gnd.n2699 gnd.n1062 99.6594
R7880 gnd.n2705 gnd.n1063 99.6594
R7881 gnd.n2709 gnd.n1064 99.6594
R7882 gnd.n2715 gnd.n1065 99.6594
R7883 gnd.n2719 gnd.n1066 99.6594
R7884 gnd.n2677 gnd.n1067 99.6594
R7885 gnd.n2688 gnd.n1059 99.6594
R7886 gnd.n2694 gnd.n1060 99.6594
R7887 gnd.n2698 gnd.n1061 99.6594
R7888 gnd.n2704 gnd.n1062 99.6594
R7889 gnd.n2708 gnd.n1063 99.6594
R7890 gnd.n2714 gnd.n1064 99.6594
R7891 gnd.n2718 gnd.n1065 99.6594
R7892 gnd.n2676 gnd.n1066 99.6594
R7893 gnd.n2672 gnd.n1067 99.6594
R7894 gnd.n3078 gnd.n3077 99.6594
R7895 gnd.n3067 gnd.n3066 99.6594
R7896 gnd.n3064 gnd.n3057 99.6594
R7897 gnd.n3055 gnd.n3054 99.6594
R7898 gnd.n3044 gnd.n3043 99.6594
R7899 gnd.n3041 gnd.n3034 99.6594
R7900 gnd.n3032 gnd.n3031 99.6594
R7901 gnd.n3022 gnd.n3021 99.6594
R7902 gnd.n3019 gnd.n3018 99.6594
R7903 gnd.n1651 gnd.n1650 99.6594
R7904 gnd.n1652 gnd.n1634 99.6594
R7905 gnd.n1670 gnd.n1669 99.6594
R7906 gnd.n1671 gnd.n1625 99.6594
R7907 gnd.n1689 gnd.n1688 99.6594
R7908 gnd.n1690 gnd.n1616 99.6594
R7909 gnd.n1708 gnd.n1707 99.6594
R7910 gnd.n1709 gnd.n1607 99.6594
R7911 gnd.n1727 gnd.n1726 99.6594
R7912 gnd.n7214 gnd.n7213 99.6594
R7913 gnd.n7209 gnd.n7208 99.6594
R7914 gnd.n7204 gnd.n7203 99.6594
R7915 gnd.n7201 gnd.n7200 99.6594
R7916 gnd.n7196 gnd.n7195 99.6594
R7917 gnd.n7193 gnd.n7192 99.6594
R7918 gnd.n7188 gnd.n7187 99.6594
R7919 gnd.n7185 gnd.n7184 99.6594
R7920 gnd.n7180 gnd.n7179 99.6594
R7921 gnd.n5265 gnd.n5188 99.6594
R7922 gnd.n5257 gnd.n5176 99.6594
R7923 gnd.n5253 gnd.n5177 99.6594
R7924 gnd.n5249 gnd.n5178 99.6594
R7925 gnd.n5245 gnd.n5179 99.6594
R7926 gnd.n5241 gnd.n5180 99.6594
R7927 gnd.n5237 gnd.n5181 99.6594
R7928 gnd.n5233 gnd.n5182 99.6594
R7929 gnd.n5229 gnd.n5183 99.6594
R7930 gnd.n5225 gnd.n5184 99.6594
R7931 gnd.n5221 gnd.n5185 99.6594
R7932 gnd.n5217 gnd.n5186 99.6594
R7933 gnd.n5268 gnd.n5267 99.6594
R7934 gnd.n5972 gnd.n4820 99.6594
R7935 gnd.n5979 gnd.n5978 99.6594
R7936 gnd.n4818 gnd.n4810 99.6594
R7937 gnd.n5986 gnd.n5985 99.6594
R7938 gnd.n4809 gnd.n4803 99.6594
R7939 gnd.n5993 gnd.n5992 99.6594
R7940 gnd.n4802 gnd.n4796 99.6594
R7941 gnd.n6000 gnd.n5999 99.6594
R7942 gnd.n4795 gnd.n4789 99.6594
R7943 gnd.n6007 gnd.n6006 99.6594
R7944 gnd.n4788 gnd.n4782 99.6594
R7945 gnd.n6014 gnd.n6013 99.6594
R7946 gnd.n4781 gnd.n4778 99.6594
R7947 gnd.n5351 gnd.n5350 99.6594
R7948 gnd.n5110 gnd.n5088 99.6594
R7949 gnd.n5116 gnd.n5089 99.6594
R7950 gnd.n5120 gnd.n5090 99.6594
R7951 gnd.n5126 gnd.n5091 99.6594
R7952 gnd.n5130 gnd.n5092 99.6594
R7953 gnd.n5136 gnd.n5093 99.6594
R7954 gnd.n5094 gnd.n5078 99.6594
R7955 gnd.n6025 gnd.n6024 99.6594
R7956 gnd.n4774 gnd.n4766 99.6594
R7957 gnd.n6032 gnd.n6031 99.6594
R7958 gnd.n4765 gnd.n4759 99.6594
R7959 gnd.n6039 gnd.n6038 99.6594
R7960 gnd.n4758 gnd.n4752 99.6594
R7961 gnd.n6046 gnd.n6045 99.6594
R7962 gnd.n4751 gnd.n4748 99.6594
R7963 gnd.n4714 gnd.n1071 99.6594
R7964 gnd.n4706 gnd.n1041 99.6594
R7965 gnd.n4702 gnd.n1042 99.6594
R7966 gnd.n4698 gnd.n1043 99.6594
R7967 gnd.n4694 gnd.n1044 99.6594
R7968 gnd.n4690 gnd.n1045 99.6594
R7969 gnd.n4686 gnd.n1046 99.6594
R7970 gnd.n4682 gnd.n1047 99.6594
R7971 gnd.n4677 gnd.n1048 99.6594
R7972 gnd.n4673 gnd.n1049 99.6594
R7973 gnd.n4669 gnd.n1050 99.6594
R7974 gnd.n4665 gnd.n1051 99.6594
R7975 gnd.n4661 gnd.n1052 99.6594
R7976 gnd.n4657 gnd.n1053 99.6594
R7977 gnd.n4653 gnd.n1054 99.6594
R7978 gnd.n4649 gnd.n1055 99.6594
R7979 gnd.n4645 gnd.n1056 99.6594
R7980 gnd.n1111 gnd.n1057 99.6594
R7981 gnd.n4637 gnd.n1058 99.6594
R7982 gnd.n3248 gnd.n3247 99.6594
R7983 gnd.n2490 gnd.n2482 99.6594
R7984 gnd.n3255 gnd.n3254 99.6594
R7985 gnd.n2481 gnd.n2475 99.6594
R7986 gnd.n3262 gnd.n3261 99.6594
R7987 gnd.n2474 gnd.n2468 99.6594
R7988 gnd.n3269 gnd.n3268 99.6594
R7989 gnd.n2467 gnd.n2461 99.6594
R7990 gnd.n3276 gnd.n3275 99.6594
R7991 gnd.n3279 gnd.n3278 99.6594
R7992 gnd.n2432 gnd.n2406 99.6594
R7993 gnd.n2436 gnd.n2407 99.6594
R7994 gnd.n2440 gnd.n2408 99.6594
R7995 gnd.n2444 gnd.n2409 99.6594
R7996 gnd.n2448 gnd.n2410 99.6594
R7997 gnd.n2452 gnd.n2411 99.6594
R7998 gnd.n2414 gnd.n2412 99.6594
R7999 gnd.n2458 gnd.n2413 99.6594
R8000 gnd.n1842 gnd.n1841 99.6594
R8001 gnd.n1850 gnd.n1849 99.6594
R8002 gnd.n1851 gnd.n1833 99.6594
R8003 gnd.n1860 gnd.n1859 99.6594
R8004 gnd.n1861 gnd.n1829 99.6594
R8005 gnd.n1871 gnd.n1870 99.6594
R8006 gnd.n1874 gnd.n1873 99.6594
R8007 gnd.n1955 gnd.n1954 99.6594
R8008 gnd.n1952 gnd.n1951 99.6594
R8009 gnd.n1947 gnd.n1946 99.6594
R8010 gnd.n1944 gnd.n1943 99.6594
R8011 gnd.n1939 gnd.n1938 99.6594
R8012 gnd.n1936 gnd.n1935 99.6594
R8013 gnd.n1931 gnd.n1930 99.6594
R8014 gnd.n1928 gnd.n1927 99.6594
R8015 gnd.n1923 gnd.n1922 99.6594
R8016 gnd.n1920 gnd.n1919 99.6594
R8017 gnd.n1913 gnd.n1912 99.6594
R8018 gnd.n154 gnd.n151 99.6594
R8019 gnd.n7258 gnd.n7257 99.6594
R8020 gnd.n150 gnd.n144 99.6594
R8021 gnd.n7265 gnd.n7264 99.6594
R8022 gnd.n143 gnd.n137 99.6594
R8023 gnd.n7272 gnd.n7271 99.6594
R8024 gnd.n136 gnd.n130 99.6594
R8025 gnd.n7279 gnd.n7278 99.6594
R8026 gnd.n129 gnd.n123 99.6594
R8027 gnd.n7286 gnd.n7285 99.6594
R8028 gnd.n122 gnd.n116 99.6594
R8029 gnd.n7296 gnd.n7295 99.6594
R8030 gnd.n115 gnd.n109 99.6594
R8031 gnd.n7303 gnd.n7302 99.6594
R8032 gnd.n108 gnd.n102 99.6594
R8033 gnd.n7310 gnd.n7309 99.6594
R8034 gnd.n101 gnd.n95 99.6594
R8035 gnd.n7317 gnd.n7316 99.6594
R8036 gnd.n93 gnd.n90 99.6594
R8037 gnd.n3126 gnd.n3125 99.6594
R8038 gnd.n3026 gnd.n2995 99.6594
R8039 gnd.n3028 gnd.n2996 99.6594
R8040 gnd.n3038 gnd.n2997 99.6594
R8041 gnd.n3049 gnd.n2998 99.6594
R8042 gnd.n3051 gnd.n2999 99.6594
R8043 gnd.n3061 gnd.n3000 99.6594
R8044 gnd.n3074 gnd.n3001 99.6594
R8045 gnd.n3075 gnd.n3002 99.6594
R8046 gnd.n3003 gnd.n2501 99.6594
R8047 gnd.n3005 gnd.n3004 99.6594
R8048 gnd.n3006 gnd.n2506 99.6594
R8049 gnd.n3007 gnd.n2512 99.6594
R8050 gnd.n3009 gnd.n2514 99.6594
R8051 gnd.n3126 gnd.n3011 99.6594
R8052 gnd.n3027 gnd.n2995 99.6594
R8053 gnd.n3037 gnd.n2996 99.6594
R8054 gnd.n3048 gnd.n2997 99.6594
R8055 gnd.n3050 gnd.n2998 99.6594
R8056 gnd.n3060 gnd.n2999 99.6594
R8057 gnd.n3073 gnd.n3000 99.6594
R8058 gnd.n3076 gnd.n3001 99.6594
R8059 gnd.n3002 gnd.n2500 99.6594
R8060 gnd.n3003 gnd.n2502 99.6594
R8061 gnd.n3005 gnd.n2505 99.6594
R8062 gnd.n3006 gnd.n2507 99.6594
R8063 gnd.n3007 gnd.n2513 99.6594
R8064 gnd.n3009 gnd.n3008 99.6594
R8065 gnd.n1659 gnd.n1639 99.6594
R8066 gnd.n1663 gnd.n1661 99.6594
R8067 gnd.n1678 gnd.n1630 99.6594
R8068 gnd.n1682 gnd.n1680 99.6594
R8069 gnd.n1697 gnd.n1621 99.6594
R8070 gnd.n1701 gnd.n1699 99.6594
R8071 gnd.n1716 gnd.n1612 99.6594
R8072 gnd.n1720 gnd.n1718 99.6594
R8073 gnd.n1733 gnd.n1601 99.6594
R8074 gnd.n1736 gnd.n1735 99.6594
R8075 gnd.n1739 gnd.n1738 99.6594
R8076 gnd.n1744 gnd.n1743 99.6594
R8077 gnd.n1747 gnd.n1746 99.6594
R8078 gnd.n4123 gnd.n4122 99.6594
R8079 gnd.n4122 gnd.n4121 99.6594
R8080 gnd.n1746 gnd.n1745 99.6594
R8081 gnd.n1743 gnd.n1742 99.6594
R8082 gnd.n1738 gnd.n1737 99.6594
R8083 gnd.n1735 gnd.n1734 99.6594
R8084 gnd.n1719 gnd.n1601 99.6594
R8085 gnd.n1718 gnd.n1717 99.6594
R8086 gnd.n1700 gnd.n1612 99.6594
R8087 gnd.n1699 gnd.n1698 99.6594
R8088 gnd.n1681 gnd.n1621 99.6594
R8089 gnd.n1680 gnd.n1679 99.6594
R8090 gnd.n1662 gnd.n1630 99.6594
R8091 gnd.n1661 gnd.n1660 99.6594
R8092 gnd.n1639 gnd.n1438 99.6594
R8093 gnd.n2508 gnd.t99 98.63
R8094 gnd.n7211 gnd.t87 98.63
R8095 gnd.n1604 gnd.t72 98.63
R8096 gnd.n3069 gnd.t94 98.63
R8097 gnd.n1879 gnd.t69 98.63
R8098 gnd.n1908 gnd.t48 98.63
R8099 gnd.n157 gnd.t33 98.63
R8100 gnd.n7289 gnd.t61 98.63
R8101 gnd.n1091 gnd.t134 98.63
R8102 gnd.n1113 gnd.t121 98.63
R8103 gnd.n2673 gnd.t118 98.63
R8104 gnd.n2487 gnd.t65 98.63
R8105 gnd.n2398 gnd.t84 98.63
R8106 gnd.n4131 gnd.t75 98.63
R8107 gnd.n2327 gnd.t108 96.6984
R8108 gnd.n1959 gnd.t58 96.6984
R8109 gnd.n2324 gnd.t30 96.6906
R8110 gnd.n3907 gnd.t110 96.6906
R8111 gnd.n2276 gnd.n2275 81.8399
R8112 gnd.n5139 gnd.t51 74.8376
R8113 gnd.n4772 gnd.t92 74.8376
R8114 gnd.n2328 gnd.t107 72.8438
R8115 gnd.n1960 gnd.t59 72.8438
R8116 gnd.n2277 gnd.n2270 72.8411
R8117 gnd.n2283 gnd.n2268 72.8411
R8118 gnd.n3903 gnd.n3902 72.8411
R8119 gnd.n2509 gnd.t98 72.836
R8120 gnd.n2325 gnd.t29 72.836
R8121 gnd.n3908 gnd.t111 72.836
R8122 gnd.n7212 gnd.t88 72.836
R8123 gnd.n1605 gnd.t71 72.836
R8124 gnd.n3070 gnd.t95 72.836
R8125 gnd.n1880 gnd.t68 72.836
R8126 gnd.n1909 gnd.t47 72.836
R8127 gnd.n158 gnd.t34 72.836
R8128 gnd.n7290 gnd.t62 72.836
R8129 gnd.n1092 gnd.t133 72.836
R8130 gnd.n1114 gnd.t120 72.836
R8131 gnd.n2674 gnd.t117 72.836
R8132 gnd.n2488 gnd.t66 72.836
R8133 gnd.n2399 gnd.t85 72.836
R8134 gnd.n4132 gnd.t76 72.836
R8135 gnd.n3971 gnd.n1787 71.676
R8136 gnd.n3967 gnd.n1788 71.676
R8137 gnd.n3963 gnd.n1789 71.676
R8138 gnd.n3959 gnd.n1790 71.676
R8139 gnd.n3955 gnd.n1791 71.676
R8140 gnd.n3951 gnd.n1792 71.676
R8141 gnd.n3947 gnd.n1793 71.676
R8142 gnd.n3943 gnd.n1794 71.676
R8143 gnd.n3939 gnd.n1795 71.676
R8144 gnd.n3935 gnd.n1796 71.676
R8145 gnd.n3931 gnd.n1797 71.676
R8146 gnd.n3927 gnd.n1798 71.676
R8147 gnd.n3923 gnd.n1799 71.676
R8148 gnd.n3919 gnd.n1800 71.676
R8149 gnd.n3914 gnd.n1801 71.676
R8150 gnd.n3910 gnd.n1802 71.676
R8151 gnd.n4047 gnd.n1821 71.676
R8152 gnd.n4043 gnd.n1820 71.676
R8153 gnd.n4038 gnd.n1819 71.676
R8154 gnd.n4034 gnd.n1818 71.676
R8155 gnd.n4030 gnd.n1817 71.676
R8156 gnd.n4026 gnd.n1816 71.676
R8157 gnd.n4022 gnd.n1815 71.676
R8158 gnd.n4018 gnd.n1814 71.676
R8159 gnd.n4014 gnd.n1813 71.676
R8160 gnd.n4010 gnd.n1812 71.676
R8161 gnd.n4006 gnd.n1811 71.676
R8162 gnd.n4002 gnd.n1810 71.676
R8163 gnd.n3998 gnd.n1809 71.676
R8164 gnd.n3994 gnd.n1808 71.676
R8165 gnd.n3990 gnd.n1807 71.676
R8166 gnd.n3986 gnd.n1806 71.676
R8167 gnd.n3982 gnd.n1805 71.676
R8168 gnd.n3350 gnd.n3349 71.676
R8169 gnd.n2323 gnd.n2290 71.676
R8170 gnd.n3342 gnd.n2291 71.676
R8171 gnd.n3338 gnd.n2292 71.676
R8172 gnd.n3334 gnd.n2293 71.676
R8173 gnd.n3330 gnd.n2294 71.676
R8174 gnd.n3326 gnd.n2295 71.676
R8175 gnd.n3322 gnd.n2296 71.676
R8176 gnd.n3318 gnd.n2297 71.676
R8177 gnd.n3314 gnd.n2298 71.676
R8178 gnd.n3310 gnd.n2299 71.676
R8179 gnd.n3306 gnd.n2300 71.676
R8180 gnd.n3302 gnd.n2301 71.676
R8181 gnd.n3298 gnd.n2302 71.676
R8182 gnd.n3294 gnd.n2303 71.676
R8183 gnd.n3290 gnd.n2304 71.676
R8184 gnd.n3286 gnd.n2306 71.676
R8185 gnd.n2392 gnd.n2307 71.676
R8186 gnd.n2387 gnd.n2308 71.676
R8187 gnd.n2383 gnd.n2309 71.676
R8188 gnd.n2379 gnd.n2310 71.676
R8189 gnd.n2375 gnd.n2311 71.676
R8190 gnd.n2371 gnd.n2312 71.676
R8191 gnd.n2367 gnd.n2313 71.676
R8192 gnd.n2363 gnd.n2314 71.676
R8193 gnd.n2359 gnd.n2315 71.676
R8194 gnd.n2355 gnd.n2316 71.676
R8195 gnd.n2351 gnd.n2317 71.676
R8196 gnd.n2347 gnd.n2318 71.676
R8197 gnd.n2343 gnd.n2319 71.676
R8198 gnd.n2339 gnd.n2320 71.676
R8199 gnd.n2335 gnd.n2321 71.676
R8200 gnd.n3349 gnd.n2288 71.676
R8201 gnd.n3343 gnd.n2290 71.676
R8202 gnd.n3339 gnd.n2291 71.676
R8203 gnd.n3335 gnd.n2292 71.676
R8204 gnd.n3331 gnd.n2293 71.676
R8205 gnd.n3327 gnd.n2294 71.676
R8206 gnd.n3323 gnd.n2295 71.676
R8207 gnd.n3319 gnd.n2296 71.676
R8208 gnd.n3315 gnd.n2297 71.676
R8209 gnd.n3311 gnd.n2298 71.676
R8210 gnd.n3307 gnd.n2299 71.676
R8211 gnd.n3303 gnd.n2300 71.676
R8212 gnd.n3299 gnd.n2301 71.676
R8213 gnd.n3295 gnd.n2302 71.676
R8214 gnd.n3291 gnd.n2303 71.676
R8215 gnd.n3287 gnd.n2305 71.676
R8216 gnd.n2393 gnd.n2306 71.676
R8217 gnd.n2388 gnd.n2307 71.676
R8218 gnd.n2384 gnd.n2308 71.676
R8219 gnd.n2380 gnd.n2309 71.676
R8220 gnd.n2376 gnd.n2310 71.676
R8221 gnd.n2372 gnd.n2311 71.676
R8222 gnd.n2368 gnd.n2312 71.676
R8223 gnd.n2364 gnd.n2313 71.676
R8224 gnd.n2360 gnd.n2314 71.676
R8225 gnd.n2356 gnd.n2315 71.676
R8226 gnd.n2352 gnd.n2316 71.676
R8227 gnd.n2348 gnd.n2317 71.676
R8228 gnd.n2344 gnd.n2318 71.676
R8229 gnd.n2340 gnd.n2319 71.676
R8230 gnd.n2336 gnd.n2320 71.676
R8231 gnd.n2332 gnd.n2321 71.676
R8232 gnd.n3985 gnd.n1805 71.676
R8233 gnd.n3989 gnd.n1806 71.676
R8234 gnd.n3993 gnd.n1807 71.676
R8235 gnd.n3997 gnd.n1808 71.676
R8236 gnd.n4001 gnd.n1809 71.676
R8237 gnd.n4005 gnd.n1810 71.676
R8238 gnd.n4009 gnd.n1811 71.676
R8239 gnd.n4013 gnd.n1812 71.676
R8240 gnd.n4017 gnd.n1813 71.676
R8241 gnd.n4021 gnd.n1814 71.676
R8242 gnd.n4025 gnd.n1815 71.676
R8243 gnd.n4029 gnd.n1816 71.676
R8244 gnd.n4033 gnd.n1817 71.676
R8245 gnd.n4037 gnd.n1818 71.676
R8246 gnd.n4042 gnd.n1819 71.676
R8247 gnd.n4046 gnd.n1820 71.676
R8248 gnd.n3909 gnd.n1803 71.676
R8249 gnd.n3913 gnd.n1802 71.676
R8250 gnd.n3918 gnd.n1801 71.676
R8251 gnd.n3922 gnd.n1800 71.676
R8252 gnd.n3926 gnd.n1799 71.676
R8253 gnd.n3930 gnd.n1798 71.676
R8254 gnd.n3934 gnd.n1797 71.676
R8255 gnd.n3938 gnd.n1796 71.676
R8256 gnd.n3942 gnd.n1795 71.676
R8257 gnd.n3946 gnd.n1794 71.676
R8258 gnd.n3950 gnd.n1793 71.676
R8259 gnd.n3954 gnd.n1792 71.676
R8260 gnd.n3958 gnd.n1791 71.676
R8261 gnd.n3962 gnd.n1790 71.676
R8262 gnd.n3966 gnd.n1789 71.676
R8263 gnd.n3970 gnd.n1788 71.676
R8264 gnd.n3973 gnd.n1787 71.676
R8265 gnd.n8 gnd.t271 69.1507
R8266 gnd.n14 gnd.t148 68.4792
R8267 gnd.n13 gnd.t138 68.4792
R8268 gnd.n12 gnd.t277 68.4792
R8269 gnd.n11 gnd.t162 68.4792
R8270 gnd.n10 gnd.t283 68.4792
R8271 gnd.n9 gnd.t152 68.4792
R8272 gnd.n8 gnd.t154 68.4792
R8273 gnd.n5266 gnd.n5170 64.369
R8274 gnd.n4740 gnd.n4739 59.5891
R8275 gnd.n7005 gnd.n320 59.5891
R8276 gnd.n2390 gnd.n2328 59.5399
R8277 gnd.n4040 gnd.n1960 59.5399
R8278 gnd.n2326 gnd.n2325 59.5399
R8279 gnd.n3916 gnd.n3908 59.5399
R8280 gnd.n3352 gnd.n2286 59.1804
R8281 gnd.n6055 gnd.n4741 57.3586
R8282 gnd.n4925 gnd.t177 56.607
R8283 gnd.n40 gnd.t252 56.607
R8284 gnd.n4902 gnd.t225 56.407
R8285 gnd.n4913 gnd.t210 56.407
R8286 gnd.n17 gnd.t243 56.407
R8287 gnd.n28 gnd.t229 56.407
R8288 gnd.n4934 gnd.t209 55.8337
R8289 gnd.n4911 gnd.t239 55.8337
R8290 gnd.n4922 gnd.t223 55.8337
R8291 gnd.n49 gnd.t268 55.8337
R8292 gnd.n26 gnd.t259 55.8337
R8293 gnd.n37 gnd.t246 55.8337
R8294 gnd.n2274 gnd.n2273 54.358
R8295 gnd.n3900 gnd.n3899 54.358
R8296 gnd.n4925 gnd.n4924 53.0052
R8297 gnd.n4927 gnd.n4926 53.0052
R8298 gnd.n4929 gnd.n4928 53.0052
R8299 gnd.n4931 gnd.n4930 53.0052
R8300 gnd.n4933 gnd.n4932 53.0052
R8301 gnd.n4902 gnd.n4901 53.0052
R8302 gnd.n4904 gnd.n4903 53.0052
R8303 gnd.n4906 gnd.n4905 53.0052
R8304 gnd.n4908 gnd.n4907 53.0052
R8305 gnd.n4910 gnd.n4909 53.0052
R8306 gnd.n4913 gnd.n4912 53.0052
R8307 gnd.n4915 gnd.n4914 53.0052
R8308 gnd.n4917 gnd.n4916 53.0052
R8309 gnd.n4919 gnd.n4918 53.0052
R8310 gnd.n4921 gnd.n4920 53.0052
R8311 gnd.n48 gnd.n47 53.0052
R8312 gnd.n46 gnd.n45 53.0052
R8313 gnd.n44 gnd.n43 53.0052
R8314 gnd.n42 gnd.n41 53.0052
R8315 gnd.n40 gnd.n39 53.0052
R8316 gnd.n25 gnd.n24 53.0052
R8317 gnd.n23 gnd.n22 53.0052
R8318 gnd.n21 gnd.n20 53.0052
R8319 gnd.n19 gnd.n18 53.0052
R8320 gnd.n17 gnd.n16 53.0052
R8321 gnd.n36 gnd.n35 53.0052
R8322 gnd.n34 gnd.n33 53.0052
R8323 gnd.n32 gnd.n31 53.0052
R8324 gnd.n30 gnd.n29 53.0052
R8325 gnd.n28 gnd.n27 53.0052
R8326 gnd.n3891 gnd.n3890 52.4801
R8327 gnd.n5900 gnd.t166 52.3082
R8328 gnd.n5868 gnd.t1 52.3082
R8329 gnd.n5836 gnd.t146 52.3082
R8330 gnd.n5805 gnd.t164 52.3082
R8331 gnd.n5773 gnd.t24 52.3082
R8332 gnd.n5741 gnd.t158 52.3082
R8333 gnd.n5709 gnd.t168 52.3082
R8334 gnd.n5678 gnd.t170 52.3082
R8335 gnd.n5730 gnd.n5698 51.4173
R8336 gnd.n5794 gnd.n5793 50.455
R8337 gnd.n5762 gnd.n5761 50.455
R8338 gnd.n5730 gnd.n5729 50.455
R8339 gnd.n5213 gnd.n5212 45.1884
R8340 gnd.n4816 gnd.n4815 45.1884
R8341 gnd.n3975 gnd.n3906 44.3322
R8342 gnd.n2277 gnd.n2276 44.3189
R8343 gnd.n6273 gnd.n6272 43.8952
R8344 gnd.n6272 gnd.n763 43.8952
R8345 gnd.n6266 gnd.n763 43.8952
R8346 gnd.n6266 gnd.n6265 43.8952
R8347 gnd.n6265 gnd.n6264 43.8952
R8348 gnd.n6264 gnd.n771 43.8952
R8349 gnd.n6258 gnd.n771 43.8952
R8350 gnd.n6258 gnd.n6257 43.8952
R8351 gnd.n6257 gnd.n6256 43.8952
R8352 gnd.n6256 gnd.n779 43.8952
R8353 gnd.n6250 gnd.n779 43.8952
R8354 gnd.n6250 gnd.n6249 43.8952
R8355 gnd.n6249 gnd.n6248 43.8952
R8356 gnd.n6248 gnd.n787 43.8952
R8357 gnd.n6242 gnd.n787 43.8952
R8358 gnd.n6242 gnd.n6241 43.8952
R8359 gnd.n6241 gnd.n6240 43.8952
R8360 gnd.n6240 gnd.n795 43.8952
R8361 gnd.n6234 gnd.n795 43.8952
R8362 gnd.n6234 gnd.n6233 43.8952
R8363 gnd.n6233 gnd.n6232 43.8952
R8364 gnd.n6232 gnd.n803 43.8952
R8365 gnd.n6226 gnd.n803 43.8952
R8366 gnd.n6226 gnd.n6225 43.8952
R8367 gnd.n6225 gnd.n6224 43.8952
R8368 gnd.n6224 gnd.n811 43.8952
R8369 gnd.n6218 gnd.n811 43.8952
R8370 gnd.n6218 gnd.n6217 43.8952
R8371 gnd.n6217 gnd.n6216 43.8952
R8372 gnd.n6216 gnd.n819 43.8952
R8373 gnd.n6210 gnd.n819 43.8952
R8374 gnd.n6210 gnd.n6209 43.8952
R8375 gnd.n6209 gnd.n6208 43.8952
R8376 gnd.n6208 gnd.n827 43.8952
R8377 gnd.n6202 gnd.n827 43.8952
R8378 gnd.n6202 gnd.n6201 43.8952
R8379 gnd.n6201 gnd.n6200 43.8952
R8380 gnd.n6200 gnd.n835 43.8952
R8381 gnd.n6194 gnd.n835 43.8952
R8382 gnd.n6194 gnd.n6193 43.8952
R8383 gnd.n6193 gnd.n6192 43.8952
R8384 gnd.n6192 gnd.n843 43.8952
R8385 gnd.n6186 gnd.n843 43.8952
R8386 gnd.n6186 gnd.n6185 43.8952
R8387 gnd.n6185 gnd.n6184 43.8952
R8388 gnd.n6184 gnd.n851 43.8952
R8389 gnd.n6178 gnd.n851 43.8952
R8390 gnd.n6178 gnd.n6177 43.8952
R8391 gnd.n6177 gnd.n6176 43.8952
R8392 gnd.n6176 gnd.n859 43.8952
R8393 gnd.n6170 gnd.n859 43.8952
R8394 gnd.n6170 gnd.n6169 43.8952
R8395 gnd.n6169 gnd.n6168 43.8952
R8396 gnd.n6168 gnd.n867 43.8952
R8397 gnd.n6162 gnd.n867 43.8952
R8398 gnd.n6162 gnd.n6161 43.8952
R8399 gnd.n6161 gnd.n6160 43.8952
R8400 gnd.n6160 gnd.n875 43.8952
R8401 gnd.n6154 gnd.n875 43.8952
R8402 gnd.n6154 gnd.n6153 43.8952
R8403 gnd.n6153 gnd.n6152 43.8952
R8404 gnd.n6152 gnd.n883 43.8952
R8405 gnd.n6146 gnd.n883 43.8952
R8406 gnd.n6146 gnd.n6145 43.8952
R8407 gnd.n6145 gnd.n6144 43.8952
R8408 gnd.n6144 gnd.n891 43.8952
R8409 gnd.n6138 gnd.n891 43.8952
R8410 gnd.n6138 gnd.n6137 43.8952
R8411 gnd.n6137 gnd.n6136 43.8952
R8412 gnd.n6136 gnd.n899 43.8952
R8413 gnd.n6130 gnd.n899 43.8952
R8414 gnd.n6130 gnd.n6129 43.8952
R8415 gnd.n6129 gnd.n6128 43.8952
R8416 gnd.n6128 gnd.n907 43.8952
R8417 gnd.n6122 gnd.n907 43.8952
R8418 gnd.n6122 gnd.n6121 43.8952
R8419 gnd.n6121 gnd.n6120 43.8952
R8420 gnd.n6120 gnd.n915 43.8952
R8421 gnd.n6114 gnd.n915 43.8952
R8422 gnd.n6114 gnd.n6113 43.8952
R8423 gnd.n6113 gnd.n6112 43.8952
R8424 gnd.n6112 gnd.n923 43.8952
R8425 gnd.n6106 gnd.n923 43.8952
R8426 gnd.n2510 gnd.n2509 42.2793
R8427 gnd.n5214 gnd.n5213 42.2793
R8428 gnd.n4817 gnd.n4816 42.2793
R8429 gnd.n5140 gnd.n5139 42.2793
R8430 gnd.n4773 gnd.n4772 42.2793
R8431 gnd.n7216 gnd.n7212 42.2793
R8432 gnd.n1606 gnd.n1605 42.2793
R8433 gnd.n3071 gnd.n3070 42.2793
R8434 gnd.n1910 gnd.n1909 42.2793
R8435 gnd.n7254 gnd.n158 42.2793
R8436 gnd.n7291 gnd.n7290 42.2793
R8437 gnd.n4679 gnd.n1092 42.2793
R8438 gnd.n1115 gnd.n1114 42.2793
R8439 gnd.n2725 gnd.n2674 42.2793
R8440 gnd.n2489 gnd.n2488 42.2793
R8441 gnd.n4133 gnd.n4132 42.2793
R8442 gnd.n2275 gnd.n2274 41.6274
R8443 gnd.n3901 gnd.n3900 41.6274
R8444 gnd.n2284 gnd.n2283 40.8975
R8445 gnd.n3904 gnd.n3903 40.8975
R8446 gnd.n1957 gnd.n1880 36.9518
R8447 gnd.n3284 gnd.n2399 36.9518
R8448 gnd.n2283 gnd.n2282 35.055
R8449 gnd.n2278 gnd.n2277 35.055
R8450 gnd.n3893 gnd.n3892 35.055
R8451 gnd.n3903 gnd.n3889 35.055
R8452 gnd.n3983 gnd.n1961 33.2493
R8453 gnd.n2333 gnd.n2330 33.2493
R8454 gnd.n5276 gnd.n5170 31.8661
R8455 gnd.n5276 gnd.n5275 31.8661
R8456 gnd.n5284 gnd.n5159 31.8661
R8457 gnd.n5292 gnd.n5159 31.8661
R8458 gnd.n5292 gnd.n5153 31.8661
R8459 gnd.n5300 gnd.n5153 31.8661
R8460 gnd.n5300 gnd.n5146 31.8661
R8461 gnd.n5338 gnd.n5146 31.8661
R8462 gnd.n5348 gnd.n5079 31.8661
R8463 gnd.n4739 gnd.n1017 31.8661
R8464 gnd.n4733 gnd.n1017 31.8661
R8465 gnd.n4733 gnd.n4732 31.8661
R8466 gnd.n4732 gnd.n4731 31.8661
R8467 gnd.n4731 gnd.n1025 31.8661
R8468 gnd.n4725 gnd.n1025 31.8661
R8469 gnd.n4725 gnd.n4724 31.8661
R8470 gnd.n4724 gnd.n4723 31.8661
R8471 gnd.n4723 gnd.n1033 31.8661
R8472 gnd.n4717 gnd.n1033 31.8661
R8473 gnd.n4717 gnd.n4716 31.8661
R8474 gnd.n1119 gnd.n1069 31.8661
R8475 gnd.n2559 gnd.n1329 31.8661
R8476 gnd.n2994 gnd.n2993 31.8661
R8477 gnd.n3128 gnd.n2994 31.8661
R8478 gnd.n3136 gnd.n2553 31.8661
R8479 gnd.n4376 gnd.n1441 31.8661
R8480 gnd.n4370 gnd.n4369 31.8661
R8481 gnd.n4369 gnd.n4368 31.8661
R8482 gnd.n4362 gnd.n1459 31.8661
R8483 gnd.n7033 gnd.n83 31.8661
R8484 gnd.n7031 gnd.n7030 31.8661
R8485 gnd.n7030 gnd.n7029 31.8661
R8486 gnd.n7029 gnd.n301 31.8661
R8487 gnd.n7023 gnd.n301 31.8661
R8488 gnd.n7023 gnd.n7022 31.8661
R8489 gnd.n7022 gnd.n7021 31.8661
R8490 gnd.n7021 gnd.n312 31.8661
R8491 gnd.n7015 gnd.n312 31.8661
R8492 gnd.n7015 gnd.n7014 31.8661
R8493 gnd.n7014 gnd.n7013 31.8661
R8494 gnd.n7013 gnd.n320 31.8661
R8495 gnd.n6106 gnd.n6105 26.3373
R8496 gnd.n2509 gnd.n2508 25.7944
R8497 gnd.n5139 gnd.n5138 25.7944
R8498 gnd.n4772 gnd.n4771 25.7944
R8499 gnd.n7212 gnd.n7211 25.7944
R8500 gnd.n1605 gnd.n1604 25.7944
R8501 gnd.n3070 gnd.n3069 25.7944
R8502 gnd.n1880 gnd.n1879 25.7944
R8503 gnd.n1909 gnd.n1908 25.7944
R8504 gnd.n158 gnd.n157 25.7944
R8505 gnd.n7290 gnd.n7289 25.7944
R8506 gnd.n1092 gnd.n1091 25.7944
R8507 gnd.n1114 gnd.n1113 25.7944
R8508 gnd.n2674 gnd.n2673 25.7944
R8509 gnd.n2488 gnd.n2487 25.7944
R8510 gnd.n2399 gnd.n2398 25.7944
R8511 gnd.n4132 gnd.n4131 25.7944
R8512 gnd.n5360 gnd.n5080 24.8557
R8513 gnd.n5370 gnd.n5063 24.8557
R8514 gnd.n5066 gnd.n5054 24.8557
R8515 gnd.n5391 gnd.n5055 24.8557
R8516 gnd.n5401 gnd.n5035 24.8557
R8517 gnd.n5411 gnd.n5410 24.8557
R8518 gnd.n5021 gnd.n5019 24.8557
R8519 gnd.n5442 gnd.n5441 24.8557
R8520 gnd.n5457 gnd.n5004 24.8557
R8521 gnd.n5511 gnd.n4943 24.8557
R8522 gnd.n5467 gnd.n4944 24.8557
R8523 gnd.n5504 gnd.n4955 24.8557
R8524 gnd.n4993 gnd.n4992 24.8557
R8525 gnd.n5498 gnd.n5497 24.8557
R8526 gnd.n4979 gnd.n4966 24.8557
R8527 gnd.n5537 gnd.n5536 24.8557
R8528 gnd.n5547 gnd.n4887 24.8557
R8529 gnd.n5559 gnd.n4879 24.8557
R8530 gnd.n5558 gnd.n4867 24.8557
R8531 gnd.n5577 gnd.n5576 24.8557
R8532 gnd.n5587 gnd.n4860 24.8557
R8533 gnd.n5600 gnd.n4848 24.8557
R8534 gnd.n5633 gnd.n5632 24.8557
R8535 gnd.n5642 gnd.n4835 24.8557
R8536 gnd.n6098 gnd.n941 24.8557
R8537 gnd.n5622 gnd.n952 24.8557
R8538 gnd.n6091 gnd.n6090 24.8557
R8539 gnd.n6084 gnd.n964 24.8557
R8540 gnd.n5947 gnd.n977 24.8557
R8541 gnd.n6077 gnd.n6076 24.8557
R8542 gnd.n6070 gnd.n989 24.8557
R8543 gnd.n6069 gnd.n992 24.8557
R8544 gnd.n5936 gnd.n1003 24.8557
R8545 gnd.n6056 gnd.n1014 24.8557
R8546 gnd.n2328 gnd.n2327 23.855
R8547 gnd.n1960 gnd.n1959 23.855
R8548 gnd.n2325 gnd.n2324 23.855
R8549 gnd.n3908 gnd.n3907 23.855
R8550 gnd.n5381 gnd.t169 23.2624
R8551 gnd.n5082 gnd.t50 22.6251
R8552 gnd.n4716 gnd.n4715 21.6691
R8553 gnd.n7031 gnd.n94 21.6691
R8554 gnd.t163 gnd.n5087 21.3504
R8555 gnd.n3353 gnd.n3352 21.0737
R8556 gnd.n3976 gnd.n3975 21.0737
R8557 gnd.n4635 gnd.n1119 21.0318
R8558 gnd.n2667 gnd.n1121 21.0318
R8559 gnd.n4626 gnd.n1130 21.0318
R8560 gnd.n2747 gnd.n1133 21.0318
R8561 gnd.n4620 gnd.n1142 21.0318
R8562 gnd.n2800 gnd.n1145 21.0318
R8563 gnd.n2808 gnd.n1154 21.0318
R8564 gnd.n4608 gnd.n1162 21.0318
R8565 gnd.n2816 gnd.n2648 21.0318
R8566 gnd.n4602 gnd.n1172 21.0318
R8567 gnd.n4596 gnd.n1183 21.0318
R8568 gnd.n2837 gnd.n1186 21.0318
R8569 gnd.n2611 gnd.n1196 21.0318
R8570 gnd.n2894 gnd.n2893 21.0318
R8571 gnd.n4582 gnd.n1204 21.0318
R8572 gnd.n2887 gnd.n1207 21.0318
R8573 gnd.n2854 gnd.n1220 21.0318
R8574 gnd.n4569 gnd.n1225 21.0318
R8575 gnd.n2877 gnd.n2876 21.0318
R8576 gnd.n4563 gnd.n1234 21.0318
R8577 gnd.n4556 gnd.n1242 21.0318
R8578 gnd.n2907 gnd.n1245 21.0318
R8579 gnd.n2915 gnd.n1255 21.0318
R8580 gnd.n4544 gnd.n1263 21.0318
R8581 gnd.n2961 gnd.n2960 21.0318
R8582 gnd.n4538 gnd.n1273 21.0318
R8583 gnd.n4532 gnd.n1284 21.0318
R8584 gnd.n2930 gnd.n1287 21.0318
R8585 gnd.n2934 gnd.n1297 21.0318
R8586 gnd.n4520 gnd.n1305 21.0318
R8587 gnd.n2943 gnd.n1308 21.0318
R8588 gnd.n4514 gnd.n1316 21.0318
R8589 gnd.n4508 gnd.n1326 21.0318
R8590 gnd.n4361 gnd.n1462 21.0318
R8591 gnd.n4355 gnd.n1474 21.0318
R8592 gnd.n4176 gnd.n4175 21.0318
R8593 gnd.n4186 gnd.n1586 21.0318
R8594 gnd.n4185 gnd.n1564 21.0318
R8595 gnd.n1568 gnd.n1555 21.0318
R8596 gnd.n4207 gnd.n1557 21.0318
R8597 gnd.n4222 gnd.n1539 21.0318
R8598 gnd.n4250 gnd.n4248 21.0318
R8599 gnd.n4213 gnd.n1530 21.0318
R8600 gnd.n4260 gnd.n1533 21.0318
R8601 gnd.n4326 gnd.n1496 21.0318
R8602 gnd.n4329 gnd.n1499 21.0318
R8603 gnd.n7113 gnd.n236 21.0318
R8604 gnd.n4299 gnd.n4298 21.0318
R8605 gnd.n4314 gnd.n1513 21.0318
R8606 gnd.n4309 gnd.n4308 21.0318
R8607 gnd.n4290 gnd.n255 21.0318
R8608 gnd.n7094 gnd.n7093 21.0318
R8609 gnd.n7098 gnd.n251 21.0318
R8610 gnd.n4282 gnd.n220 21.0318
R8611 gnd.n7084 gnd.n211 21.0318
R8612 gnd.n7130 gnd.n214 21.0318
R8613 gnd.n7138 gnd.n205 21.0318
R8614 gnd.n7074 gnd.n7073 21.0318
R8615 gnd.n7146 gnd.n197 21.0318
R8616 gnd.n7048 gnd.n188 21.0318
R8617 gnd.n7065 gnd.n179 21.0318
R8618 gnd.n7162 gnd.n182 21.0318
R8619 gnd.n7059 gnd.n169 21.0318
R8620 gnd.n7172 gnd.n171 21.0318
R8621 gnd.n7247 gnd.n81 21.0318
R8622 gnd.n7326 gnd.n83 21.0318
R8623 gnd.n5615 gnd.t10 20.7131
R8624 gnd.n4590 gnd.t178 20.7131
R8625 gnd.t202 gnd.n1237 20.7131
R8626 gnd.t220 gnd.n233 20.7131
R8627 gnd.n7122 gnd.t234 20.7131
R8628 gnd.n2559 gnd.n2459 20.3945
R8629 gnd.n1459 gnd.n1451 20.3945
R8630 gnd.t12 gnd.n4841 20.0758
R8631 gnd.n4614 gnd.t208 20.0758
R8632 gnd.t190 gnd.n1276 20.0758
R8633 gnd.n4223 gnd.t200 20.0758
R8634 gnd.n7154 gnd.t245 20.0758
R8635 gnd.n2271 gnd.t82 19.8005
R8636 gnd.n2271 gnd.t128 19.8005
R8637 gnd.n2272 gnd.t105 19.8005
R8638 gnd.n2272 gnd.t55 19.8005
R8639 gnd.n3897 gnd.t41 19.8005
R8640 gnd.n3897 gnd.t114 19.8005
R8641 gnd.n3898 gnd.t131 19.8005
R8642 gnd.n3898 gnd.t102 19.8005
R8643 gnd.n2268 gnd.n2267 19.5087
R8644 gnd.n2281 gnd.n2268 19.5087
R8645 gnd.n2279 gnd.n2270 19.5087
R8646 gnd.n3902 gnd.n3896 19.5087
R8647 gnd.n5548 gnd.t15 19.4385
R8648 gnd.n3215 gnd.n3214 19.3944
R8649 gnd.n3214 gnd.n3213 19.3944
R8650 gnd.n3213 gnd.n2520 19.3944
R8651 gnd.n3209 gnd.n2520 19.3944
R8652 gnd.n3209 gnd.n3208 19.3944
R8653 gnd.n3208 gnd.n3207 19.3944
R8654 gnd.n3207 gnd.n2525 19.3944
R8655 gnd.n3203 gnd.n2525 19.3944
R8656 gnd.n3203 gnd.n3202 19.3944
R8657 gnd.n3202 gnd.n3201 19.3944
R8658 gnd.n3201 gnd.n2530 19.3944
R8659 gnd.n3197 gnd.n2530 19.3944
R8660 gnd.n3197 gnd.n3196 19.3944
R8661 gnd.n3196 gnd.n3195 19.3944
R8662 gnd.n3195 gnd.n3185 19.3944
R8663 gnd.n3191 gnd.n3185 19.3944
R8664 gnd.n3191 gnd.n3190 19.3944
R8665 gnd.n3190 gnd.n2232 19.3944
R8666 gnd.n3462 gnd.n2232 19.3944
R8667 gnd.n3462 gnd.n2230 19.3944
R8668 gnd.n3466 gnd.n2230 19.3944
R8669 gnd.n3466 gnd.n2212 19.3944
R8670 gnd.n3493 gnd.n2212 19.3944
R8671 gnd.n3493 gnd.n2209 19.3944
R8672 gnd.n3498 gnd.n2209 19.3944
R8673 gnd.n3498 gnd.n2210 19.3944
R8674 gnd.n2210 gnd.n2182 19.3944
R8675 gnd.n3529 gnd.n2182 19.3944
R8676 gnd.n3529 gnd.n2180 19.3944
R8677 gnd.n3533 gnd.n2180 19.3944
R8678 gnd.n3533 gnd.n2161 19.3944
R8679 gnd.n3557 gnd.n2161 19.3944
R8680 gnd.n3557 gnd.n2158 19.3944
R8681 gnd.n3562 gnd.n2158 19.3944
R8682 gnd.n3562 gnd.n2159 19.3944
R8683 gnd.n2159 gnd.n2131 19.3944
R8684 gnd.n3595 gnd.n2131 19.3944
R8685 gnd.n3595 gnd.n2128 19.3944
R8686 gnd.n3614 gnd.n2128 19.3944
R8687 gnd.n3614 gnd.n2129 19.3944
R8688 gnd.n3610 gnd.n2129 19.3944
R8689 gnd.n3610 gnd.n3609 19.3944
R8690 gnd.n3609 gnd.n3608 19.3944
R8691 gnd.n3608 gnd.n3602 19.3944
R8692 gnd.n3604 gnd.n3602 19.3944
R8693 gnd.n3604 gnd.n2081 19.3944
R8694 gnd.n3678 gnd.n2081 19.3944
R8695 gnd.n3679 gnd.n3678 19.3944
R8696 gnd.n3679 gnd.n2079 19.3944
R8697 gnd.n3683 gnd.n2079 19.3944
R8698 gnd.n3683 gnd.n2055 19.3944
R8699 gnd.n3732 gnd.n2055 19.3944
R8700 gnd.n3732 gnd.n2056 19.3944
R8701 gnd.n3728 gnd.n2056 19.3944
R8702 gnd.n3728 gnd.n2032 19.3944
R8703 gnd.n3772 gnd.n2032 19.3944
R8704 gnd.n3772 gnd.n2033 19.3944
R8705 gnd.n3768 gnd.n2033 19.3944
R8706 gnd.n3768 gnd.n2010 19.3944
R8707 gnd.n3811 gnd.n2010 19.3944
R8708 gnd.n3811 gnd.n2011 19.3944
R8709 gnd.n3807 gnd.n2011 19.3944
R8710 gnd.n3807 gnd.n1986 19.3944
R8711 gnd.n3859 gnd.n1986 19.3944
R8712 gnd.n3859 gnd.n1987 19.3944
R8713 gnd.n3855 gnd.n1987 19.3944
R8714 gnd.n3855 gnd.n3854 19.3944
R8715 gnd.n3854 gnd.n1784 19.3944
R8716 gnd.n4052 gnd.n1784 19.3944
R8717 gnd.n4052 gnd.n1782 19.3944
R8718 gnd.n4056 gnd.n1782 19.3944
R8719 gnd.n4056 gnd.n1773 19.3944
R8720 gnd.n4073 gnd.n1773 19.3944
R8721 gnd.n4073 gnd.n1771 19.3944
R8722 gnd.n4077 gnd.n1771 19.3944
R8723 gnd.n4077 gnd.n1761 19.3944
R8724 gnd.n4094 gnd.n1761 19.3944
R8725 gnd.n4094 gnd.n1759 19.3944
R8726 gnd.n4099 gnd.n1759 19.3944
R8727 gnd.n4099 gnd.n1750 19.3944
R8728 gnd.n4117 gnd.n1750 19.3944
R8729 gnd.n4118 gnd.n4117 19.3944
R8730 gnd.n3221 gnd.n3220 19.3944
R8731 gnd.n3220 gnd.n3219 19.3944
R8732 gnd.n3219 gnd.n2515 19.3944
R8733 gnd.n3124 gnd.n3123 19.3944
R8734 gnd.n3123 gnd.n3013 19.3944
R8735 gnd.n3116 gnd.n3013 19.3944
R8736 gnd.n3116 gnd.n3115 19.3944
R8737 gnd.n3115 gnd.n3029 19.3944
R8738 gnd.n3108 gnd.n3029 19.3944
R8739 gnd.n3108 gnd.n3107 19.3944
R8740 gnd.n3107 gnd.n3039 19.3944
R8741 gnd.n3100 gnd.n3039 19.3944
R8742 gnd.n3100 gnd.n3099 19.3944
R8743 gnd.n3099 gnd.n3052 19.3944
R8744 gnd.n3092 gnd.n3052 19.3944
R8745 gnd.n3092 gnd.n3091 19.3944
R8746 gnd.n3091 gnd.n3062 19.3944
R8747 gnd.n3084 gnd.n3062 19.3944
R8748 gnd.n3084 gnd.n3083 19.3944
R8749 gnd.n3083 gnd.n2499 19.3944
R8750 gnd.n3232 gnd.n2499 19.3944
R8751 gnd.n3232 gnd.n3231 19.3944
R8752 gnd.n3231 gnd.n3230 19.3944
R8753 gnd.n3230 gnd.n2503 19.3944
R8754 gnd.n3226 gnd.n2503 19.3944
R8755 gnd.n3226 gnd.n3225 19.3944
R8756 gnd.n3225 gnd.n3224 19.3944
R8757 gnd.n5263 gnd.n5262 19.3944
R8758 gnd.n5262 gnd.n5261 19.3944
R8759 gnd.n5261 gnd.n5260 19.3944
R8760 gnd.n5260 gnd.n5258 19.3944
R8761 gnd.n5258 gnd.n5255 19.3944
R8762 gnd.n5255 gnd.n5254 19.3944
R8763 gnd.n5254 gnd.n5251 19.3944
R8764 gnd.n5251 gnd.n5250 19.3944
R8765 gnd.n5250 gnd.n5247 19.3944
R8766 gnd.n5247 gnd.n5246 19.3944
R8767 gnd.n5246 gnd.n5243 19.3944
R8768 gnd.n5243 gnd.n5242 19.3944
R8769 gnd.n5242 gnd.n5239 19.3944
R8770 gnd.n5239 gnd.n5238 19.3944
R8771 gnd.n5238 gnd.n5235 19.3944
R8772 gnd.n5235 gnd.n5234 19.3944
R8773 gnd.n5234 gnd.n5231 19.3944
R8774 gnd.n5231 gnd.n5230 19.3944
R8775 gnd.n5230 gnd.n5227 19.3944
R8776 gnd.n5227 gnd.n5226 19.3944
R8777 gnd.n5226 gnd.n5223 19.3944
R8778 gnd.n5223 gnd.n5222 19.3944
R8779 gnd.n5219 gnd.n5218 19.3944
R8780 gnd.n5218 gnd.n5174 19.3944
R8781 gnd.n5269 gnd.n5174 19.3944
R8782 gnd.n5976 gnd.n4819 19.3944
R8783 gnd.n5976 gnd.n5975 19.3944
R8784 gnd.n5975 gnd.n5974 19.3944
R8785 gnd.n6018 gnd.n6017 19.3944
R8786 gnd.n6017 gnd.n6016 19.3944
R8787 gnd.n6016 gnd.n4780 19.3944
R8788 gnd.n6011 gnd.n4780 19.3944
R8789 gnd.n6011 gnd.n6010 19.3944
R8790 gnd.n6010 gnd.n6009 19.3944
R8791 gnd.n6009 gnd.n4787 19.3944
R8792 gnd.n6004 gnd.n4787 19.3944
R8793 gnd.n6004 gnd.n6003 19.3944
R8794 gnd.n6003 gnd.n6002 19.3944
R8795 gnd.n6002 gnd.n4794 19.3944
R8796 gnd.n5997 gnd.n4794 19.3944
R8797 gnd.n5997 gnd.n5996 19.3944
R8798 gnd.n5996 gnd.n5995 19.3944
R8799 gnd.n5995 gnd.n4801 19.3944
R8800 gnd.n5990 gnd.n4801 19.3944
R8801 gnd.n5990 gnd.n5989 19.3944
R8802 gnd.n5989 gnd.n5988 19.3944
R8803 gnd.n5988 gnd.n4808 19.3944
R8804 gnd.n5983 gnd.n4808 19.3944
R8805 gnd.n5983 gnd.n5982 19.3944
R8806 gnd.n5982 gnd.n5981 19.3944
R8807 gnd.n5362 gnd.n5071 19.3944
R8808 gnd.n5372 gnd.n5071 19.3944
R8809 gnd.n5373 gnd.n5372 19.3944
R8810 gnd.n5373 gnd.n5052 19.3944
R8811 gnd.n5393 gnd.n5052 19.3944
R8812 gnd.n5393 gnd.n5044 19.3944
R8813 gnd.n5403 gnd.n5044 19.3944
R8814 gnd.n5404 gnd.n5403 19.3944
R8815 gnd.n5405 gnd.n5404 19.3944
R8816 gnd.n5405 gnd.n5027 19.3944
R8817 gnd.n5422 gnd.n5027 19.3944
R8818 gnd.n5425 gnd.n5422 19.3944
R8819 gnd.n5425 gnd.n5424 19.3944
R8820 gnd.n5424 gnd.n5000 19.3944
R8821 gnd.n5464 gnd.n5000 19.3944
R8822 gnd.n5464 gnd.n4997 19.3944
R8823 gnd.n5470 gnd.n4997 19.3944
R8824 gnd.n5471 gnd.n5470 19.3944
R8825 gnd.n5471 gnd.n4995 19.3944
R8826 gnd.n5477 gnd.n4995 19.3944
R8827 gnd.n5480 gnd.n5477 19.3944
R8828 gnd.n5482 gnd.n5480 19.3944
R8829 gnd.n5488 gnd.n5482 19.3944
R8830 gnd.n5488 gnd.n5487 19.3944
R8831 gnd.n5487 gnd.n4882 19.3944
R8832 gnd.n5554 gnd.n4882 19.3944
R8833 gnd.n5555 gnd.n5554 19.3944
R8834 gnd.n5555 gnd.n4875 19.3944
R8835 gnd.n5566 gnd.n4875 19.3944
R8836 gnd.n5567 gnd.n5566 19.3944
R8837 gnd.n5567 gnd.n4858 19.3944
R8838 gnd.n4858 gnd.n4856 19.3944
R8839 gnd.n5591 gnd.n4856 19.3944
R8840 gnd.n5594 gnd.n5591 19.3944
R8841 gnd.n5594 gnd.n5593 19.3944
R8842 gnd.n5593 gnd.n4832 19.3944
R8843 gnd.n5645 gnd.n4832 19.3944
R8844 gnd.n5646 gnd.n5645 19.3944
R8845 gnd.n5646 gnd.n4830 19.3944
R8846 gnd.n5652 gnd.n4830 19.3944
R8847 gnd.n5654 gnd.n5652 19.3944
R8848 gnd.n5658 gnd.n5654 19.3944
R8849 gnd.n5659 gnd.n5658 19.3944
R8850 gnd.n5945 gnd.n5659 19.3944
R8851 gnd.n5945 gnd.n5944 19.3944
R8852 gnd.n5944 gnd.n5943 19.3944
R8853 gnd.n5943 gnd.n5940 19.3944
R8854 gnd.n5940 gnd.n5939 19.3944
R8855 gnd.n5939 gnd.n5938 19.3944
R8856 gnd.n5938 gnd.n5935 19.3944
R8857 gnd.n5935 gnd.n5934 19.3944
R8858 gnd.n5934 gnd.n5931 19.3944
R8859 gnd.n5931 gnd.n5930 19.3944
R8860 gnd.n5353 gnd.n5352 19.3944
R8861 gnd.n5352 gnd.n5085 19.3944
R8862 gnd.n5108 gnd.n5085 19.3944
R8863 gnd.n5111 gnd.n5108 19.3944
R8864 gnd.n5111 gnd.n5104 19.3944
R8865 gnd.n5115 gnd.n5104 19.3944
R8866 gnd.n5118 gnd.n5115 19.3944
R8867 gnd.n5121 gnd.n5118 19.3944
R8868 gnd.n5121 gnd.n5102 19.3944
R8869 gnd.n5125 gnd.n5102 19.3944
R8870 gnd.n5128 gnd.n5125 19.3944
R8871 gnd.n5131 gnd.n5128 19.3944
R8872 gnd.n5131 gnd.n5100 19.3944
R8873 gnd.n5135 gnd.n5100 19.3944
R8874 gnd.n5358 gnd.n5357 19.3944
R8875 gnd.n5357 gnd.n5061 19.3944
R8876 gnd.n5383 gnd.n5061 19.3944
R8877 gnd.n5383 gnd.n5059 19.3944
R8878 gnd.n5389 gnd.n5059 19.3944
R8879 gnd.n5389 gnd.n5388 19.3944
R8880 gnd.n5388 gnd.n5033 19.3944
R8881 gnd.n5413 gnd.n5033 19.3944
R8882 gnd.n5413 gnd.n5031 19.3944
R8883 gnd.n5417 gnd.n5031 19.3944
R8884 gnd.n5417 gnd.n5011 19.3944
R8885 gnd.n5444 gnd.n5011 19.3944
R8886 gnd.n5444 gnd.n5009 19.3944
R8887 gnd.n5454 gnd.n5009 19.3944
R8888 gnd.n5454 gnd.n5453 19.3944
R8889 gnd.n5453 gnd.n5452 19.3944
R8890 gnd.n5452 gnd.n4958 19.3944
R8891 gnd.n5502 gnd.n4958 19.3944
R8892 gnd.n5502 gnd.n5501 19.3944
R8893 gnd.n5501 gnd.n5500 19.3944
R8894 gnd.n5500 gnd.n4962 19.3944
R8895 gnd.n4982 gnd.n4962 19.3944
R8896 gnd.n4982 gnd.n4892 19.3944
R8897 gnd.n5539 gnd.n4892 19.3944
R8898 gnd.n5539 gnd.n4890 19.3944
R8899 gnd.n5545 gnd.n4890 19.3944
R8900 gnd.n5545 gnd.n5544 19.3944
R8901 gnd.n5544 gnd.n4865 19.3944
R8902 gnd.n5579 gnd.n4865 19.3944
R8903 gnd.n5579 gnd.n4863 19.3944
R8904 gnd.n5585 gnd.n4863 19.3944
R8905 gnd.n5585 gnd.n5584 19.3944
R8906 gnd.n5584 gnd.n4839 19.3944
R8907 gnd.n5635 gnd.n4839 19.3944
R8908 gnd.n5635 gnd.n4837 19.3944
R8909 gnd.n5640 gnd.n4837 19.3944
R8910 gnd.n5640 gnd.n946 19.3944
R8911 gnd.n6095 gnd.n946 19.3944
R8912 gnd.n6095 gnd.n6094 19.3944
R8913 gnd.n6094 gnd.n6093 19.3944
R8914 gnd.n6093 gnd.n950 19.3944
R8915 gnd.n969 gnd.n950 19.3944
R8916 gnd.n6081 gnd.n969 19.3944
R8917 gnd.n6081 gnd.n6080 19.3944
R8918 gnd.n6080 gnd.n6079 19.3944
R8919 gnd.n6079 gnd.n975 19.3944
R8920 gnd.n995 gnd.n975 19.3944
R8921 gnd.n6067 gnd.n995 19.3944
R8922 gnd.n6067 gnd.n6066 19.3944
R8923 gnd.n6066 gnd.n6065 19.3944
R8924 gnd.n6065 gnd.n1001 19.3944
R8925 gnd.n4744 gnd.n1001 19.3944
R8926 gnd.n6053 gnd.n4744 19.3944
R8927 gnd.n6050 gnd.n6049 19.3944
R8928 gnd.n6049 gnd.n6048 19.3944
R8929 gnd.n6048 gnd.n4750 19.3944
R8930 gnd.n6043 gnd.n4750 19.3944
R8931 gnd.n6043 gnd.n6042 19.3944
R8932 gnd.n6042 gnd.n6041 19.3944
R8933 gnd.n6041 gnd.n4757 19.3944
R8934 gnd.n6036 gnd.n4757 19.3944
R8935 gnd.n6036 gnd.n6035 19.3944
R8936 gnd.n6035 gnd.n6034 19.3944
R8937 gnd.n6034 gnd.n4764 19.3944
R8938 gnd.n6029 gnd.n4764 19.3944
R8939 gnd.n6029 gnd.n6028 19.3944
R8940 gnd.n6028 gnd.n6027 19.3944
R8941 gnd.n5273 gnd.n5172 19.3944
R8942 gnd.n5273 gnd.n5163 19.3944
R8943 gnd.n5286 gnd.n5163 19.3944
R8944 gnd.n5286 gnd.n5161 19.3944
R8945 gnd.n5290 gnd.n5161 19.3944
R8946 gnd.n5290 gnd.n5151 19.3944
R8947 gnd.n5302 gnd.n5151 19.3944
R8948 gnd.n5302 gnd.n5149 19.3944
R8949 gnd.n5336 gnd.n5149 19.3944
R8950 gnd.n5336 gnd.n5335 19.3944
R8951 gnd.n5335 gnd.n5334 19.3944
R8952 gnd.n5334 gnd.n5333 19.3944
R8953 gnd.n5333 gnd.n5330 19.3944
R8954 gnd.n5330 gnd.n5329 19.3944
R8955 gnd.n5329 gnd.n5328 19.3944
R8956 gnd.n5328 gnd.n5326 19.3944
R8957 gnd.n5326 gnd.n5325 19.3944
R8958 gnd.n5325 gnd.n5322 19.3944
R8959 gnd.n5322 gnd.n5321 19.3944
R8960 gnd.n5321 gnd.n5320 19.3944
R8961 gnd.n5320 gnd.n5318 19.3944
R8962 gnd.n5318 gnd.n5017 19.3944
R8963 gnd.n5433 gnd.n5017 19.3944
R8964 gnd.n5433 gnd.n5015 19.3944
R8965 gnd.n5439 gnd.n5015 19.3944
R8966 gnd.n5439 gnd.n5438 19.3944
R8967 gnd.n5438 gnd.n4939 19.3944
R8968 gnd.n5513 gnd.n4939 19.3944
R8969 gnd.n5513 gnd.n4940 19.3944
R8970 gnd.n4987 gnd.n4986 19.3944
R8971 gnd.n4990 gnd.n4989 19.3944
R8972 gnd.n4977 gnd.n4976 19.3944
R8973 gnd.n5532 gnd.n4897 19.3944
R8974 gnd.n5532 gnd.n5531 19.3944
R8975 gnd.n5531 gnd.n5530 19.3944
R8976 gnd.n5530 gnd.n5528 19.3944
R8977 gnd.n5528 gnd.n5527 19.3944
R8978 gnd.n5527 gnd.n5525 19.3944
R8979 gnd.n5525 gnd.n5524 19.3944
R8980 gnd.n5524 gnd.n4846 19.3944
R8981 gnd.n5602 gnd.n4846 19.3944
R8982 gnd.n5602 gnd.n4844 19.3944
R8983 gnd.n5630 gnd.n4844 19.3944
R8984 gnd.n5630 gnd.n5629 19.3944
R8985 gnd.n5629 gnd.n5628 19.3944
R8986 gnd.n5628 gnd.n5626 19.3944
R8987 gnd.n5626 gnd.n5625 19.3944
R8988 gnd.n5625 gnd.n5619 19.3944
R8989 gnd.n5619 gnd.n5618 19.3944
R8990 gnd.n5618 gnd.n5617 19.3944
R8991 gnd.n5617 gnd.n5614 19.3944
R8992 gnd.n5614 gnd.n4829 19.3944
R8993 gnd.n5951 gnd.n4829 19.3944
R8994 gnd.n5951 gnd.n4827 19.3944
R8995 gnd.n5957 gnd.n4827 19.3944
R8996 gnd.n5958 gnd.n5957 19.3944
R8997 gnd.n5961 gnd.n5958 19.3944
R8998 gnd.n5961 gnd.n4825 19.3944
R8999 gnd.n5965 gnd.n4825 19.3944
R9000 gnd.n5968 gnd.n5965 19.3944
R9001 gnd.n5969 gnd.n5968 19.3944
R9002 gnd.n5278 gnd.n5168 19.3944
R9003 gnd.n5278 gnd.n5166 19.3944
R9004 gnd.n5282 gnd.n5166 19.3944
R9005 gnd.n5282 gnd.n5157 19.3944
R9006 gnd.n5294 gnd.n5157 19.3944
R9007 gnd.n5294 gnd.n5155 19.3944
R9008 gnd.n5298 gnd.n5155 19.3944
R9009 gnd.n5298 gnd.n5144 19.3944
R9010 gnd.n5340 gnd.n5144 19.3944
R9011 gnd.n5340 gnd.n5098 19.3944
R9012 gnd.n5346 gnd.n5098 19.3944
R9013 gnd.n5346 gnd.n5345 19.3944
R9014 gnd.n5345 gnd.n5076 19.3944
R9015 gnd.n5367 gnd.n5076 19.3944
R9016 gnd.n5367 gnd.n5069 19.3944
R9017 gnd.n5378 gnd.n5069 19.3944
R9018 gnd.n5378 gnd.n5377 19.3944
R9019 gnd.n5377 gnd.n5050 19.3944
R9020 gnd.n5398 gnd.n5050 19.3944
R9021 gnd.n5398 gnd.n5040 19.3944
R9022 gnd.n5408 gnd.n5040 19.3944
R9023 gnd.n5408 gnd.n5023 19.3944
R9024 gnd.n5429 gnd.n5023 19.3944
R9025 gnd.n5429 gnd.n5428 19.3944
R9026 gnd.n5428 gnd.n5002 19.3944
R9027 gnd.n5459 gnd.n5002 19.3944
R9028 gnd.n5459 gnd.n4947 19.3944
R9029 gnd.n5509 gnd.n4947 19.3944
R9030 gnd.n5509 gnd.n5508 19.3944
R9031 gnd.n5508 gnd.n5507 19.3944
R9032 gnd.n5507 gnd.n4951 19.3944
R9033 gnd.n4969 gnd.n4951 19.3944
R9034 gnd.n5495 gnd.n4969 19.3944
R9035 gnd.n5495 gnd.n5494 19.3944
R9036 gnd.n5494 gnd.n5493 19.3944
R9037 gnd.n5493 gnd.n4973 19.3944
R9038 gnd.n4973 gnd.n4884 19.3944
R9039 gnd.n5550 gnd.n4884 19.3944
R9040 gnd.n5550 gnd.n4877 19.3944
R9041 gnd.n5561 gnd.n4877 19.3944
R9042 gnd.n5561 gnd.n4873 19.3944
R9043 gnd.n5574 gnd.n4873 19.3944
R9044 gnd.n5574 gnd.n5573 19.3944
R9045 gnd.n5573 gnd.n4852 19.3944
R9046 gnd.n5598 gnd.n4852 19.3944
R9047 gnd.n5598 gnd.n5597 19.3944
R9048 gnd.n5597 gnd.n935 19.3944
R9049 gnd.n6102 gnd.n935 19.3944
R9050 gnd.n6102 gnd.n6101 19.3944
R9051 gnd.n6101 gnd.n6100 19.3944
R9052 gnd.n6100 gnd.n939 19.3944
R9053 gnd.n958 gnd.n939 19.3944
R9054 gnd.n6088 gnd.n958 19.3944
R9055 gnd.n6088 gnd.n6087 19.3944
R9056 gnd.n6087 gnd.n6086 19.3944
R9057 gnd.n6086 gnd.n962 19.3944
R9058 gnd.n983 gnd.n962 19.3944
R9059 gnd.n6074 gnd.n983 19.3944
R9060 gnd.n6074 gnd.n6073 19.3944
R9061 gnd.n6073 gnd.n6072 19.3944
R9062 gnd.n6072 gnd.n987 19.3944
R9063 gnd.n1009 gnd.n987 19.3944
R9064 gnd.n6060 gnd.n1009 19.3944
R9065 gnd.n6060 gnd.n6059 19.3944
R9066 gnd.n6059 gnd.n6058 19.3944
R9067 gnd.n4146 gnd.n1597 19.3944
R9068 gnd.n4146 gnd.n1592 19.3944
R9069 gnd.n4178 gnd.n1592 19.3944
R9070 gnd.n4178 gnd.n1589 19.3944
R9071 gnd.n4183 gnd.n1589 19.3944
R9072 gnd.n4183 gnd.n1590 19.3944
R9073 gnd.n1590 gnd.n1553 19.3944
R9074 gnd.n4209 gnd.n1553 19.3944
R9075 gnd.n4209 gnd.n1550 19.3944
R9076 gnd.n4220 gnd.n1550 19.3944
R9077 gnd.n4220 gnd.n1551 19.3944
R9078 gnd.n4216 gnd.n1551 19.3944
R9079 gnd.n4216 gnd.n4215 19.3944
R9080 gnd.n4215 gnd.n1505 19.3944
R9081 gnd.n4324 gnd.n1505 19.3944
R9082 gnd.n4324 gnd.n1506 19.3944
R9083 gnd.n4320 gnd.n1506 19.3944
R9084 gnd.n4320 gnd.n4319 19.3944
R9085 gnd.n4319 gnd.n4318 19.3944
R9086 gnd.n4318 gnd.n4316 19.3944
R9087 gnd.n4316 gnd.n52 19.3944
R9088 gnd.n7358 gnd.n52 19.3944
R9089 gnd.n7358 gnd.n7357 19.3944
R9090 gnd.n7357 gnd.n7356 19.3944
R9091 gnd.n7356 gnd.n57 19.3944
R9092 gnd.n7352 gnd.n57 19.3944
R9093 gnd.n7352 gnd.n7351 19.3944
R9094 gnd.n7351 gnd.n7350 19.3944
R9095 gnd.n7350 gnd.n62 19.3944
R9096 gnd.n7346 gnd.n62 19.3944
R9097 gnd.n7346 gnd.n7345 19.3944
R9098 gnd.n7345 gnd.n7344 19.3944
R9099 gnd.n7344 gnd.n67 19.3944
R9100 gnd.n7340 gnd.n67 19.3944
R9101 gnd.n7340 gnd.n7339 19.3944
R9102 gnd.n7339 gnd.n7338 19.3944
R9103 gnd.n7338 gnd.n72 19.3944
R9104 gnd.n7334 gnd.n72 19.3944
R9105 gnd.n7334 gnd.n7333 19.3944
R9106 gnd.n7333 gnd.n7332 19.3944
R9107 gnd.n7332 gnd.n77 19.3944
R9108 gnd.n7328 gnd.n77 19.3944
R9109 gnd.n7241 gnd.n7240 19.3944
R9110 gnd.n7240 gnd.n7239 19.3944
R9111 gnd.n7239 gnd.n7182 19.3944
R9112 gnd.n7235 gnd.n7182 19.3944
R9113 gnd.n7235 gnd.n7234 19.3944
R9114 gnd.n7234 gnd.n7233 19.3944
R9115 gnd.n7233 gnd.n7190 19.3944
R9116 gnd.n7229 gnd.n7190 19.3944
R9117 gnd.n7229 gnd.n7228 19.3944
R9118 gnd.n7228 gnd.n7227 19.3944
R9119 gnd.n7227 gnd.n7198 19.3944
R9120 gnd.n7223 gnd.n7198 19.3944
R9121 gnd.n7223 gnd.n7222 19.3944
R9122 gnd.n7222 gnd.n7221 19.3944
R9123 gnd.n7221 gnd.n7206 19.3944
R9124 gnd.n7217 gnd.n7206 19.3944
R9125 gnd.n1648 gnd.n1642 19.3944
R9126 gnd.n1654 gnd.n1642 19.3944
R9127 gnd.n1654 gnd.n1635 19.3944
R9128 gnd.n1667 gnd.n1635 19.3944
R9129 gnd.n1667 gnd.n1633 19.3944
R9130 gnd.n1673 gnd.n1633 19.3944
R9131 gnd.n1673 gnd.n1626 19.3944
R9132 gnd.n1686 gnd.n1626 19.3944
R9133 gnd.n1686 gnd.n1624 19.3944
R9134 gnd.n1692 gnd.n1624 19.3944
R9135 gnd.n1692 gnd.n1617 19.3944
R9136 gnd.n1705 gnd.n1617 19.3944
R9137 gnd.n1705 gnd.n1615 19.3944
R9138 gnd.n1711 gnd.n1615 19.3944
R9139 gnd.n1711 gnd.n1608 19.3944
R9140 gnd.n1724 gnd.n1608 19.3944
R9141 gnd.n1645 gnd.n1477 19.3944
R9142 gnd.n4353 gnd.n1477 19.3944
R9143 gnd.n4353 gnd.n1478 19.3944
R9144 gnd.n4349 gnd.n1478 19.3944
R9145 gnd.n4349 gnd.n4348 19.3944
R9146 gnd.n4348 gnd.n4347 19.3944
R9147 gnd.n4347 gnd.n1484 19.3944
R9148 gnd.n4343 gnd.n1484 19.3944
R9149 gnd.n4343 gnd.n4342 19.3944
R9150 gnd.n4342 gnd.n4341 19.3944
R9151 gnd.n4341 gnd.n1489 19.3944
R9152 gnd.n4337 gnd.n1489 19.3944
R9153 gnd.n4337 gnd.n4336 19.3944
R9154 gnd.n4336 gnd.n4335 19.3944
R9155 gnd.n4335 gnd.n1494 19.3944
R9156 gnd.n4331 gnd.n1494 19.3944
R9157 gnd.n4331 gnd.n239 19.3944
R9158 gnd.n7111 gnd.n239 19.3944
R9159 gnd.n7111 gnd.n240 19.3944
R9160 gnd.n7107 gnd.n240 19.3944
R9161 gnd.n7107 gnd.n7106 19.3944
R9162 gnd.n7106 gnd.n7105 19.3944
R9163 gnd.n7105 gnd.n246 19.3944
R9164 gnd.n7101 gnd.n246 19.3944
R9165 gnd.n7101 gnd.n7100 19.3944
R9166 gnd.n7100 gnd.n218 19.3944
R9167 gnd.n7124 gnd.n218 19.3944
R9168 gnd.n7124 gnd.n216 19.3944
R9169 gnd.n7128 gnd.n216 19.3944
R9170 gnd.n7128 gnd.n201 19.3944
R9171 gnd.n7140 gnd.n201 19.3944
R9172 gnd.n7140 gnd.n199 19.3944
R9173 gnd.n7144 gnd.n199 19.3944
R9174 gnd.n7144 gnd.n186 19.3944
R9175 gnd.n7156 gnd.n186 19.3944
R9176 gnd.n7156 gnd.n184 19.3944
R9177 gnd.n7160 gnd.n184 19.3944
R9178 gnd.n7160 gnd.n167 19.3944
R9179 gnd.n7174 gnd.n167 19.3944
R9180 gnd.n7174 gnd.n164 19.3944
R9181 gnd.n7245 gnd.n164 19.3944
R9182 gnd.n7245 gnd.n165 19.3944
R9183 gnd.n3017 gnd.n1332 19.3944
R9184 gnd.n3017 gnd.n3016 19.3944
R9185 gnd.n3120 gnd.n3016 19.3944
R9186 gnd.n3120 gnd.n3119 19.3944
R9187 gnd.n3119 gnd.n3024 19.3944
R9188 gnd.n3112 gnd.n3024 19.3944
R9189 gnd.n3112 gnd.n3111 19.3944
R9190 gnd.n3111 gnd.n3035 19.3944
R9191 gnd.n3104 gnd.n3035 19.3944
R9192 gnd.n3104 gnd.n3103 19.3944
R9193 gnd.n3103 gnd.n3046 19.3944
R9194 gnd.n3096 gnd.n3046 19.3944
R9195 gnd.n3096 gnd.n3095 19.3944
R9196 gnd.n3095 gnd.n3058 19.3944
R9197 gnd.n3088 gnd.n3058 19.3944
R9198 gnd.n3088 gnd.n3087 19.3944
R9199 gnd.n6797 gnd.n449 19.3944
R9200 gnd.n6801 gnd.n449 19.3944
R9201 gnd.n6801 gnd.n445 19.3944
R9202 gnd.n6807 gnd.n445 19.3944
R9203 gnd.n6807 gnd.n443 19.3944
R9204 gnd.n6811 gnd.n443 19.3944
R9205 gnd.n6811 gnd.n439 19.3944
R9206 gnd.n6817 gnd.n439 19.3944
R9207 gnd.n6817 gnd.n437 19.3944
R9208 gnd.n6821 gnd.n437 19.3944
R9209 gnd.n6821 gnd.n433 19.3944
R9210 gnd.n6827 gnd.n433 19.3944
R9211 gnd.n6827 gnd.n431 19.3944
R9212 gnd.n6831 gnd.n431 19.3944
R9213 gnd.n6831 gnd.n427 19.3944
R9214 gnd.n6837 gnd.n427 19.3944
R9215 gnd.n6837 gnd.n425 19.3944
R9216 gnd.n6841 gnd.n425 19.3944
R9217 gnd.n6841 gnd.n421 19.3944
R9218 gnd.n6847 gnd.n421 19.3944
R9219 gnd.n6847 gnd.n419 19.3944
R9220 gnd.n6851 gnd.n419 19.3944
R9221 gnd.n6851 gnd.n415 19.3944
R9222 gnd.n6857 gnd.n415 19.3944
R9223 gnd.n6857 gnd.n413 19.3944
R9224 gnd.n6861 gnd.n413 19.3944
R9225 gnd.n6861 gnd.n409 19.3944
R9226 gnd.n6867 gnd.n409 19.3944
R9227 gnd.n6867 gnd.n407 19.3944
R9228 gnd.n6871 gnd.n407 19.3944
R9229 gnd.n6871 gnd.n403 19.3944
R9230 gnd.n6877 gnd.n403 19.3944
R9231 gnd.n6877 gnd.n401 19.3944
R9232 gnd.n6881 gnd.n401 19.3944
R9233 gnd.n6881 gnd.n397 19.3944
R9234 gnd.n6887 gnd.n397 19.3944
R9235 gnd.n6887 gnd.n395 19.3944
R9236 gnd.n6891 gnd.n395 19.3944
R9237 gnd.n6891 gnd.n391 19.3944
R9238 gnd.n6897 gnd.n391 19.3944
R9239 gnd.n6897 gnd.n389 19.3944
R9240 gnd.n6901 gnd.n389 19.3944
R9241 gnd.n6901 gnd.n385 19.3944
R9242 gnd.n6907 gnd.n385 19.3944
R9243 gnd.n6907 gnd.n383 19.3944
R9244 gnd.n6911 gnd.n383 19.3944
R9245 gnd.n6911 gnd.n379 19.3944
R9246 gnd.n6917 gnd.n379 19.3944
R9247 gnd.n6917 gnd.n377 19.3944
R9248 gnd.n6921 gnd.n377 19.3944
R9249 gnd.n6921 gnd.n373 19.3944
R9250 gnd.n6927 gnd.n373 19.3944
R9251 gnd.n6927 gnd.n371 19.3944
R9252 gnd.n6931 gnd.n371 19.3944
R9253 gnd.n6931 gnd.n367 19.3944
R9254 gnd.n6937 gnd.n367 19.3944
R9255 gnd.n6937 gnd.n365 19.3944
R9256 gnd.n6941 gnd.n365 19.3944
R9257 gnd.n6941 gnd.n361 19.3944
R9258 gnd.n6947 gnd.n361 19.3944
R9259 gnd.n6947 gnd.n359 19.3944
R9260 gnd.n6951 gnd.n359 19.3944
R9261 gnd.n6951 gnd.n355 19.3944
R9262 gnd.n6957 gnd.n355 19.3944
R9263 gnd.n6957 gnd.n353 19.3944
R9264 gnd.n6961 gnd.n353 19.3944
R9265 gnd.n6961 gnd.n349 19.3944
R9266 gnd.n6967 gnd.n349 19.3944
R9267 gnd.n6967 gnd.n347 19.3944
R9268 gnd.n6971 gnd.n347 19.3944
R9269 gnd.n6971 gnd.n343 19.3944
R9270 gnd.n6977 gnd.n343 19.3944
R9271 gnd.n6977 gnd.n341 19.3944
R9272 gnd.n6981 gnd.n341 19.3944
R9273 gnd.n6981 gnd.n337 19.3944
R9274 gnd.n6987 gnd.n337 19.3944
R9275 gnd.n6987 gnd.n335 19.3944
R9276 gnd.n6991 gnd.n335 19.3944
R9277 gnd.n6991 gnd.n331 19.3944
R9278 gnd.n6997 gnd.n331 19.3944
R9279 gnd.n6997 gnd.n329 19.3944
R9280 gnd.n7001 gnd.n329 19.3944
R9281 gnd.n7001 gnd.n325 19.3944
R9282 gnd.n7007 gnd.n325 19.3944
R9283 gnd.n6276 gnd.n760 19.3944
R9284 gnd.n6280 gnd.n760 19.3944
R9285 gnd.n6280 gnd.n756 19.3944
R9286 gnd.n6286 gnd.n756 19.3944
R9287 gnd.n6286 gnd.n754 19.3944
R9288 gnd.n6290 gnd.n754 19.3944
R9289 gnd.n6290 gnd.n750 19.3944
R9290 gnd.n6296 gnd.n750 19.3944
R9291 gnd.n6296 gnd.n748 19.3944
R9292 gnd.n6300 gnd.n748 19.3944
R9293 gnd.n6300 gnd.n744 19.3944
R9294 gnd.n6306 gnd.n744 19.3944
R9295 gnd.n6306 gnd.n742 19.3944
R9296 gnd.n6310 gnd.n742 19.3944
R9297 gnd.n6310 gnd.n738 19.3944
R9298 gnd.n6316 gnd.n738 19.3944
R9299 gnd.n6316 gnd.n736 19.3944
R9300 gnd.n6320 gnd.n736 19.3944
R9301 gnd.n6320 gnd.n732 19.3944
R9302 gnd.n6326 gnd.n732 19.3944
R9303 gnd.n6326 gnd.n730 19.3944
R9304 gnd.n6330 gnd.n730 19.3944
R9305 gnd.n6330 gnd.n726 19.3944
R9306 gnd.n6336 gnd.n726 19.3944
R9307 gnd.n6336 gnd.n724 19.3944
R9308 gnd.n6340 gnd.n724 19.3944
R9309 gnd.n6340 gnd.n720 19.3944
R9310 gnd.n6346 gnd.n720 19.3944
R9311 gnd.n6346 gnd.n718 19.3944
R9312 gnd.n6350 gnd.n718 19.3944
R9313 gnd.n6350 gnd.n714 19.3944
R9314 gnd.n6356 gnd.n714 19.3944
R9315 gnd.n6356 gnd.n712 19.3944
R9316 gnd.n6360 gnd.n712 19.3944
R9317 gnd.n6360 gnd.n708 19.3944
R9318 gnd.n6366 gnd.n708 19.3944
R9319 gnd.n6366 gnd.n706 19.3944
R9320 gnd.n6370 gnd.n706 19.3944
R9321 gnd.n6370 gnd.n702 19.3944
R9322 gnd.n6376 gnd.n702 19.3944
R9323 gnd.n6376 gnd.n700 19.3944
R9324 gnd.n6380 gnd.n700 19.3944
R9325 gnd.n6380 gnd.n696 19.3944
R9326 gnd.n6386 gnd.n696 19.3944
R9327 gnd.n6386 gnd.n694 19.3944
R9328 gnd.n6390 gnd.n694 19.3944
R9329 gnd.n6390 gnd.n690 19.3944
R9330 gnd.n6396 gnd.n690 19.3944
R9331 gnd.n6396 gnd.n688 19.3944
R9332 gnd.n6400 gnd.n688 19.3944
R9333 gnd.n6400 gnd.n684 19.3944
R9334 gnd.n6406 gnd.n684 19.3944
R9335 gnd.n6406 gnd.n682 19.3944
R9336 gnd.n6410 gnd.n682 19.3944
R9337 gnd.n6410 gnd.n678 19.3944
R9338 gnd.n6416 gnd.n678 19.3944
R9339 gnd.n6416 gnd.n676 19.3944
R9340 gnd.n6420 gnd.n676 19.3944
R9341 gnd.n6420 gnd.n672 19.3944
R9342 gnd.n6426 gnd.n672 19.3944
R9343 gnd.n6426 gnd.n670 19.3944
R9344 gnd.n6430 gnd.n670 19.3944
R9345 gnd.n6430 gnd.n666 19.3944
R9346 gnd.n6436 gnd.n666 19.3944
R9347 gnd.n6436 gnd.n664 19.3944
R9348 gnd.n6440 gnd.n664 19.3944
R9349 gnd.n6440 gnd.n660 19.3944
R9350 gnd.n6446 gnd.n660 19.3944
R9351 gnd.n6446 gnd.n658 19.3944
R9352 gnd.n6450 gnd.n658 19.3944
R9353 gnd.n6450 gnd.n654 19.3944
R9354 gnd.n6456 gnd.n654 19.3944
R9355 gnd.n6456 gnd.n652 19.3944
R9356 gnd.n6460 gnd.n652 19.3944
R9357 gnd.n6460 gnd.n648 19.3944
R9358 gnd.n6466 gnd.n648 19.3944
R9359 gnd.n6466 gnd.n646 19.3944
R9360 gnd.n6470 gnd.n646 19.3944
R9361 gnd.n6470 gnd.n642 19.3944
R9362 gnd.n6476 gnd.n642 19.3944
R9363 gnd.n6476 gnd.n640 19.3944
R9364 gnd.n6480 gnd.n640 19.3944
R9365 gnd.n6480 gnd.n636 19.3944
R9366 gnd.n6486 gnd.n636 19.3944
R9367 gnd.n6486 gnd.n634 19.3944
R9368 gnd.n6490 gnd.n634 19.3944
R9369 gnd.n6490 gnd.n630 19.3944
R9370 gnd.n6496 gnd.n630 19.3944
R9371 gnd.n6496 gnd.n628 19.3944
R9372 gnd.n6500 gnd.n628 19.3944
R9373 gnd.n6500 gnd.n624 19.3944
R9374 gnd.n6506 gnd.n624 19.3944
R9375 gnd.n6506 gnd.n622 19.3944
R9376 gnd.n6510 gnd.n622 19.3944
R9377 gnd.n6510 gnd.n618 19.3944
R9378 gnd.n6516 gnd.n618 19.3944
R9379 gnd.n6516 gnd.n616 19.3944
R9380 gnd.n6520 gnd.n616 19.3944
R9381 gnd.n6520 gnd.n612 19.3944
R9382 gnd.n6526 gnd.n612 19.3944
R9383 gnd.n6526 gnd.n610 19.3944
R9384 gnd.n6530 gnd.n610 19.3944
R9385 gnd.n6530 gnd.n606 19.3944
R9386 gnd.n6536 gnd.n606 19.3944
R9387 gnd.n6536 gnd.n604 19.3944
R9388 gnd.n6540 gnd.n604 19.3944
R9389 gnd.n6540 gnd.n600 19.3944
R9390 gnd.n6546 gnd.n600 19.3944
R9391 gnd.n6546 gnd.n598 19.3944
R9392 gnd.n6550 gnd.n598 19.3944
R9393 gnd.n6550 gnd.n594 19.3944
R9394 gnd.n6556 gnd.n594 19.3944
R9395 gnd.n6556 gnd.n592 19.3944
R9396 gnd.n6560 gnd.n592 19.3944
R9397 gnd.n6560 gnd.n588 19.3944
R9398 gnd.n6566 gnd.n588 19.3944
R9399 gnd.n6566 gnd.n586 19.3944
R9400 gnd.n6570 gnd.n586 19.3944
R9401 gnd.n6570 gnd.n582 19.3944
R9402 gnd.n6576 gnd.n582 19.3944
R9403 gnd.n6576 gnd.n580 19.3944
R9404 gnd.n6580 gnd.n580 19.3944
R9405 gnd.n6580 gnd.n576 19.3944
R9406 gnd.n6586 gnd.n576 19.3944
R9407 gnd.n6586 gnd.n574 19.3944
R9408 gnd.n6590 gnd.n574 19.3944
R9409 gnd.n6590 gnd.n570 19.3944
R9410 gnd.n6596 gnd.n570 19.3944
R9411 gnd.n6596 gnd.n568 19.3944
R9412 gnd.n6600 gnd.n568 19.3944
R9413 gnd.n6600 gnd.n564 19.3944
R9414 gnd.n6606 gnd.n564 19.3944
R9415 gnd.n6606 gnd.n562 19.3944
R9416 gnd.n6610 gnd.n562 19.3944
R9417 gnd.n6610 gnd.n558 19.3944
R9418 gnd.n6616 gnd.n558 19.3944
R9419 gnd.n6616 gnd.n556 19.3944
R9420 gnd.n6620 gnd.n556 19.3944
R9421 gnd.n6620 gnd.n552 19.3944
R9422 gnd.n6626 gnd.n552 19.3944
R9423 gnd.n6626 gnd.n550 19.3944
R9424 gnd.n6630 gnd.n550 19.3944
R9425 gnd.n6630 gnd.n546 19.3944
R9426 gnd.n6636 gnd.n546 19.3944
R9427 gnd.n6636 gnd.n544 19.3944
R9428 gnd.n6640 gnd.n544 19.3944
R9429 gnd.n6640 gnd.n540 19.3944
R9430 gnd.n6646 gnd.n540 19.3944
R9431 gnd.n6646 gnd.n538 19.3944
R9432 gnd.n6650 gnd.n538 19.3944
R9433 gnd.n6650 gnd.n534 19.3944
R9434 gnd.n6656 gnd.n534 19.3944
R9435 gnd.n6656 gnd.n532 19.3944
R9436 gnd.n6660 gnd.n532 19.3944
R9437 gnd.n6660 gnd.n528 19.3944
R9438 gnd.n6666 gnd.n528 19.3944
R9439 gnd.n6666 gnd.n526 19.3944
R9440 gnd.n6670 gnd.n526 19.3944
R9441 gnd.n6670 gnd.n522 19.3944
R9442 gnd.n6676 gnd.n522 19.3944
R9443 gnd.n6676 gnd.n520 19.3944
R9444 gnd.n6680 gnd.n520 19.3944
R9445 gnd.n6680 gnd.n516 19.3944
R9446 gnd.n6686 gnd.n516 19.3944
R9447 gnd.n6686 gnd.n514 19.3944
R9448 gnd.n6690 gnd.n514 19.3944
R9449 gnd.n6690 gnd.n510 19.3944
R9450 gnd.n6696 gnd.n510 19.3944
R9451 gnd.n6696 gnd.n508 19.3944
R9452 gnd.n6700 gnd.n508 19.3944
R9453 gnd.n6700 gnd.n504 19.3944
R9454 gnd.n6706 gnd.n504 19.3944
R9455 gnd.n6706 gnd.n502 19.3944
R9456 gnd.n6710 gnd.n502 19.3944
R9457 gnd.n6710 gnd.n498 19.3944
R9458 gnd.n6716 gnd.n498 19.3944
R9459 gnd.n6716 gnd.n496 19.3944
R9460 gnd.n6720 gnd.n496 19.3944
R9461 gnd.n6720 gnd.n492 19.3944
R9462 gnd.n6726 gnd.n492 19.3944
R9463 gnd.n6726 gnd.n490 19.3944
R9464 gnd.n6730 gnd.n490 19.3944
R9465 gnd.n6730 gnd.n486 19.3944
R9466 gnd.n6736 gnd.n486 19.3944
R9467 gnd.n6736 gnd.n484 19.3944
R9468 gnd.n6740 gnd.n484 19.3944
R9469 gnd.n6740 gnd.n480 19.3944
R9470 gnd.n6746 gnd.n480 19.3944
R9471 gnd.n6746 gnd.n478 19.3944
R9472 gnd.n6750 gnd.n478 19.3944
R9473 gnd.n6750 gnd.n474 19.3944
R9474 gnd.n6756 gnd.n474 19.3944
R9475 gnd.n6756 gnd.n472 19.3944
R9476 gnd.n6760 gnd.n472 19.3944
R9477 gnd.n6760 gnd.n468 19.3944
R9478 gnd.n6766 gnd.n468 19.3944
R9479 gnd.n6766 gnd.n466 19.3944
R9480 gnd.n6770 gnd.n466 19.3944
R9481 gnd.n6770 gnd.n462 19.3944
R9482 gnd.n6776 gnd.n462 19.3944
R9483 gnd.n6776 gnd.n460 19.3944
R9484 gnd.n6780 gnd.n460 19.3944
R9485 gnd.n6780 gnd.n456 19.3944
R9486 gnd.n6786 gnd.n456 19.3944
R9487 gnd.n6786 gnd.n454 19.3944
R9488 gnd.n6791 gnd.n454 19.3944
R9489 gnd.n6791 gnd.n6790 19.3944
R9490 gnd.n1843 gnd.n1840 19.3944
R9491 gnd.n1843 gnd.n1838 19.3944
R9492 gnd.n1847 gnd.n1838 19.3944
R9493 gnd.n1847 gnd.n1836 19.3944
R9494 gnd.n1853 gnd.n1836 19.3944
R9495 gnd.n1853 gnd.n1834 19.3944
R9496 gnd.n1857 gnd.n1834 19.3944
R9497 gnd.n1857 gnd.n1832 19.3944
R9498 gnd.n1863 gnd.n1832 19.3944
R9499 gnd.n1863 gnd.n1830 19.3944
R9500 gnd.n1868 gnd.n1830 19.3944
R9501 gnd.n1868 gnd.n1828 19.3944
R9502 gnd.n1828 gnd.n1825 19.3944
R9503 gnd.n1875 gnd.n1825 19.3944
R9504 gnd.n1875 gnd.n1822 19.3944
R9505 gnd.n1956 gnd.n1882 19.3944
R9506 gnd.n1950 gnd.n1882 19.3944
R9507 gnd.n1950 gnd.n1949 19.3944
R9508 gnd.n1949 gnd.n1948 19.3944
R9509 gnd.n1948 gnd.n1888 19.3944
R9510 gnd.n1942 gnd.n1888 19.3944
R9511 gnd.n1942 gnd.n1941 19.3944
R9512 gnd.n1941 gnd.n1940 19.3944
R9513 gnd.n1940 gnd.n1894 19.3944
R9514 gnd.n1934 gnd.n1894 19.3944
R9515 gnd.n1934 gnd.n1933 19.3944
R9516 gnd.n1933 gnd.n1932 19.3944
R9517 gnd.n1932 gnd.n1900 19.3944
R9518 gnd.n1926 gnd.n1900 19.3944
R9519 gnd.n1926 gnd.n1925 19.3944
R9520 gnd.n1925 gnd.n1924 19.3944
R9521 gnd.n1924 gnd.n1906 19.3944
R9522 gnd.n1918 gnd.n1906 19.3944
R9523 gnd.n4150 gnd.n1596 19.3944
R9524 gnd.n4150 gnd.n1594 19.3944
R9525 gnd.n4173 gnd.n1594 19.3944
R9526 gnd.n4173 gnd.n4172 19.3944
R9527 gnd.n4172 gnd.n4171 19.3944
R9528 gnd.n4171 gnd.n4170 19.3944
R9529 gnd.n4170 gnd.n4169 19.3944
R9530 gnd.n4169 gnd.n4167 19.3944
R9531 gnd.n4167 gnd.n4166 19.3944
R9532 gnd.n4166 gnd.n4163 19.3944
R9533 gnd.n4163 gnd.n4162 19.3944
R9534 gnd.n4162 gnd.n1527 19.3944
R9535 gnd.n4262 gnd.n1527 19.3944
R9536 gnd.n4262 gnd.n1525 19.3944
R9537 gnd.n4266 gnd.n1525 19.3944
R9538 gnd.n4267 gnd.n4266 19.3944
R9539 gnd.n4270 gnd.n4267 19.3944
R9540 gnd.n4270 gnd.n1523 19.3944
R9541 gnd.n4296 gnd.n1523 19.3944
R9542 gnd.n4296 gnd.n4295 19.3944
R9543 gnd.n4295 gnd.n4294 19.3944
R9544 gnd.n4294 gnd.n4293 19.3944
R9545 gnd.n4293 gnd.n4287 19.3944
R9546 gnd.n4287 gnd.n4286 19.3944
R9547 gnd.n4286 gnd.n4285 19.3944
R9548 gnd.n4285 gnd.n4284 19.3944
R9549 gnd.n4284 gnd.n263 19.3944
R9550 gnd.n7082 gnd.n263 19.3944
R9551 gnd.n7082 gnd.n7081 19.3944
R9552 gnd.n7081 gnd.n7080 19.3944
R9553 gnd.n7080 gnd.n7077 19.3944
R9554 gnd.n7077 gnd.n7076 19.3944
R9555 gnd.n7076 gnd.n269 19.3944
R9556 gnd.n7050 gnd.n269 19.3944
R9557 gnd.n7050 gnd.n7046 19.3944
R9558 gnd.n7063 gnd.n7046 19.3944
R9559 gnd.n7063 gnd.n7062 19.3944
R9560 gnd.n7062 gnd.n7061 19.3944
R9561 gnd.n7061 gnd.n7058 19.3944
R9562 gnd.n7058 gnd.n160 19.3944
R9563 gnd.n7249 gnd.n160 19.3944
R9564 gnd.n7250 gnd.n7249 19.3944
R9565 gnd.n7288 gnd.n121 19.3944
R9566 gnd.n7283 gnd.n121 19.3944
R9567 gnd.n7283 gnd.n7282 19.3944
R9568 gnd.n7282 gnd.n7281 19.3944
R9569 gnd.n7281 gnd.n128 19.3944
R9570 gnd.n7276 gnd.n128 19.3944
R9571 gnd.n7276 gnd.n7275 19.3944
R9572 gnd.n7275 gnd.n7274 19.3944
R9573 gnd.n7274 gnd.n135 19.3944
R9574 gnd.n7269 gnd.n135 19.3944
R9575 gnd.n7269 gnd.n7268 19.3944
R9576 gnd.n7268 gnd.n7267 19.3944
R9577 gnd.n7267 gnd.n142 19.3944
R9578 gnd.n7262 gnd.n142 19.3944
R9579 gnd.n7262 gnd.n7261 19.3944
R9580 gnd.n7261 gnd.n7260 19.3944
R9581 gnd.n7260 gnd.n149 19.3944
R9582 gnd.n7255 gnd.n149 19.3944
R9583 gnd.n7321 gnd.n7320 19.3944
R9584 gnd.n7320 gnd.n7319 19.3944
R9585 gnd.n7319 gnd.n92 19.3944
R9586 gnd.n7314 gnd.n92 19.3944
R9587 gnd.n7314 gnd.n7313 19.3944
R9588 gnd.n7313 gnd.n7312 19.3944
R9589 gnd.n7312 gnd.n100 19.3944
R9590 gnd.n7307 gnd.n100 19.3944
R9591 gnd.n7307 gnd.n7306 19.3944
R9592 gnd.n7306 gnd.n7305 19.3944
R9593 gnd.n7305 gnd.n107 19.3944
R9594 gnd.n7300 gnd.n107 19.3944
R9595 gnd.n7300 gnd.n7299 19.3944
R9596 gnd.n7299 gnd.n7298 19.3944
R9597 gnd.n7298 gnd.n114 19.3944
R9598 gnd.n7293 gnd.n114 19.3944
R9599 gnd.n7293 gnd.n7292 19.3944
R9600 gnd.n4359 gnd.n4358 19.3944
R9601 gnd.n4358 gnd.n4357 19.3944
R9602 gnd.n4357 gnd.n1469 19.3944
R9603 gnd.n1584 gnd.n1469 19.3944
R9604 gnd.n1584 gnd.n1562 19.3944
R9605 gnd.n4199 gnd.n1562 19.3944
R9606 gnd.n4199 gnd.n1560 19.3944
R9607 gnd.n4205 gnd.n1560 19.3944
R9608 gnd.n4205 gnd.n4204 19.3944
R9609 gnd.n4204 gnd.n1537 19.3944
R9610 gnd.n4252 gnd.n1537 19.3944
R9611 gnd.n4252 gnd.n1535 19.3944
R9612 gnd.n4258 gnd.n1535 19.3944
R9613 gnd.n4258 gnd.n4257 19.3944
R9614 gnd.n4257 gnd.n1501 19.3944
R9615 gnd.n1501 gnd.n230 19.3944
R9616 gnd.n7116 gnd.n7115 19.3944
R9617 gnd.n4312 gnd.n4311 19.3944
R9618 gnd.n1516 gnd.n1515 19.3944
R9619 gnd.n254 gnd.n253 19.3944
R9620 gnd.n7096 gnd.n223 19.3944
R9621 gnd.n7120 gnd.n223 19.3944
R9622 gnd.n7120 gnd.n209 19.3944
R9623 gnd.n7132 gnd.n209 19.3944
R9624 gnd.n7132 gnd.n207 19.3944
R9625 gnd.n7136 gnd.n207 19.3944
R9626 gnd.n7136 gnd.n193 19.3944
R9627 gnd.n7148 gnd.n193 19.3944
R9628 gnd.n7148 gnd.n191 19.3944
R9629 gnd.n7152 gnd.n191 19.3944
R9630 gnd.n7152 gnd.n177 19.3944
R9631 gnd.n7164 gnd.n177 19.3944
R9632 gnd.n7164 gnd.n175 19.3944
R9633 gnd.n7170 gnd.n175 19.3944
R9634 gnd.n7170 gnd.n7169 19.3944
R9635 gnd.n7169 gnd.n87 19.3944
R9636 gnd.n7324 gnd.n87 19.3944
R9637 gnd.n4737 gnd.n4736 19.3944
R9638 gnd.n4736 gnd.n4735 19.3944
R9639 gnd.n4735 gnd.n1023 19.3944
R9640 gnd.n4729 gnd.n1023 19.3944
R9641 gnd.n4729 gnd.n4728 19.3944
R9642 gnd.n4728 gnd.n4727 19.3944
R9643 gnd.n4727 gnd.n1031 19.3944
R9644 gnd.n4721 gnd.n1031 19.3944
R9645 gnd.n4721 gnd.n4720 19.3944
R9646 gnd.n4720 gnd.n4719 19.3944
R9647 gnd.n4719 gnd.n1039 19.3944
R9648 gnd.n2761 gnd.n1039 19.3944
R9649 gnd.n2761 gnd.n2758 19.3944
R9650 gnd.n2765 gnd.n2758 19.3944
R9651 gnd.n2765 gnd.n2756 19.3944
R9652 gnd.n2769 gnd.n2756 19.3944
R9653 gnd.n2769 gnd.n2660 19.3944
R9654 gnd.n2773 gnd.n2660 19.3944
R9655 gnd.n2773 gnd.n2658 19.3944
R9656 gnd.n2797 gnd.n2658 19.3944
R9657 gnd.n2797 gnd.n2796 19.3944
R9658 gnd.n2796 gnd.n2795 19.3944
R9659 gnd.n2795 gnd.n2779 19.3944
R9660 gnd.n2791 gnd.n2779 19.3944
R9661 gnd.n2791 gnd.n2790 19.3944
R9662 gnd.n2790 gnd.n2789 19.3944
R9663 gnd.n2789 gnd.n2786 19.3944
R9664 gnd.n2786 gnd.n2607 19.3944
R9665 gnd.n2897 gnd.n2607 19.3944
R9666 gnd.n2897 gnd.n2608 19.3944
R9667 gnd.n2621 gnd.n2620 19.3944
R9668 gnd.n2884 gnd.n2883 19.3944
R9669 gnd.n2880 gnd.n2879 19.3944
R9670 gnd.n2627 gnd.n2626 19.3944
R9671 gnd.n2623 gnd.n2600 19.3944
R9672 gnd.n2904 gnd.n2600 19.3944
R9673 gnd.n2904 gnd.n2903 19.3944
R9674 gnd.n2903 gnd.n2575 19.3944
R9675 gnd.n2963 gnd.n2575 19.3944
R9676 gnd.n2963 gnd.n2573 19.3944
R9677 gnd.n2967 gnd.n2573 19.3944
R9678 gnd.n2967 gnd.n2571 19.3944
R9679 gnd.n2971 gnd.n2571 19.3944
R9680 gnd.n2971 gnd.n2569 19.3944
R9681 gnd.n2975 gnd.n2569 19.3944
R9682 gnd.n2975 gnd.n2567 19.3944
R9683 gnd.n2979 gnd.n2567 19.3944
R9684 gnd.n2979 gnd.n2565 19.3944
R9685 gnd.n2983 gnd.n2565 19.3944
R9686 gnd.n2983 gnd.n2563 19.3944
R9687 gnd.n2987 gnd.n2563 19.3944
R9688 gnd.n2987 gnd.n2561 19.3944
R9689 gnd.n2991 gnd.n2561 19.3944
R9690 gnd.n2991 gnd.n2557 19.3944
R9691 gnd.n3130 gnd.n2557 19.3944
R9692 gnd.n3130 gnd.n2555 19.3944
R9693 gnd.n3134 gnd.n2555 19.3944
R9694 gnd.n3134 gnd.n2551 19.3944
R9695 gnd.n3144 gnd.n2551 19.3944
R9696 gnd.n3144 gnd.n2549 19.3944
R9697 gnd.n3148 gnd.n2549 19.3944
R9698 gnd.n3148 gnd.n2543 19.3944
R9699 gnd.n3158 gnd.n2543 19.3944
R9700 gnd.n3158 gnd.n2541 19.3944
R9701 gnd.n3162 gnd.n2541 19.3944
R9702 gnd.n3162 gnd.n2535 19.3944
R9703 gnd.n3172 gnd.n2535 19.3944
R9704 gnd.n3172 gnd.n2533 19.3944
R9705 gnd.n3176 gnd.n2533 19.3944
R9706 gnd.n3176 gnd.n2258 19.3944
R9707 gnd.n3361 gnd.n2258 19.3944
R9708 gnd.n3361 gnd.n2256 19.3944
R9709 gnd.n3365 gnd.n2256 19.3944
R9710 gnd.n3365 gnd.n2240 19.3944
R9711 gnd.n3452 gnd.n2240 19.3944
R9712 gnd.n3452 gnd.n2238 19.3944
R9713 gnd.n3456 gnd.n2238 19.3944
R9714 gnd.n3456 gnd.n2219 19.3944
R9715 gnd.n3483 gnd.n2219 19.3944
R9716 gnd.n3483 gnd.n2217 19.3944
R9717 gnd.n3487 gnd.n2217 19.3944
R9718 gnd.n3487 gnd.n2197 19.3944
R9719 gnd.n3511 gnd.n2197 19.3944
R9720 gnd.n3511 gnd.n2195 19.3944
R9721 gnd.n3517 gnd.n2195 19.3944
R9722 gnd.n3517 gnd.n3516 19.3944
R9723 gnd.n3516 gnd.n2168 19.3944
R9724 gnd.n3548 gnd.n2168 19.3944
R9725 gnd.n3548 gnd.n2166 19.3944
R9726 gnd.n3552 gnd.n2166 19.3944
R9727 gnd.n3552 gnd.n2145 19.3944
R9728 gnd.n3576 gnd.n2145 19.3944
R9729 gnd.n3576 gnd.n2143 19.3944
R9730 gnd.n3582 gnd.n2143 19.3944
R9731 gnd.n3582 gnd.n3581 19.3944
R9732 gnd.n3581 gnd.n2116 19.3944
R9733 gnd.n3627 gnd.n2116 19.3944
R9734 gnd.n3627 gnd.n2114 19.3944
R9735 gnd.n3631 gnd.n2114 19.3944
R9736 gnd.n3631 gnd.n2095 19.3944
R9737 gnd.n3657 gnd.n2095 19.3944
R9738 gnd.n3657 gnd.n2093 19.3944
R9739 gnd.n3663 gnd.n2093 19.3944
R9740 gnd.n3663 gnd.n3662 19.3944
R9741 gnd.n3662 gnd.n2065 19.3944
R9742 gnd.n3707 gnd.n2065 19.3944
R9743 gnd.n3707 gnd.n2063 19.3944
R9744 gnd.n3711 gnd.n2063 19.3944
R9745 gnd.n3711 gnd.n2042 19.3944
R9746 gnd.n3747 gnd.n2042 19.3944
R9747 gnd.n3747 gnd.n2040 19.3944
R9748 gnd.n3751 gnd.n2040 19.3944
R9749 gnd.n3751 gnd.n2019 19.3944
R9750 gnd.n3786 gnd.n2019 19.3944
R9751 gnd.n3786 gnd.n2017 19.3944
R9752 gnd.n3790 gnd.n2017 19.3944
R9753 gnd.n3790 gnd.n1997 19.3944
R9754 gnd.n3827 gnd.n1997 19.3944
R9755 gnd.n3827 gnd.n1995 19.3944
R9756 gnd.n3831 gnd.n1995 19.3944
R9757 gnd.n3831 gnd.n1975 19.3944
R9758 gnd.n3872 gnd.n1975 19.3944
R9759 gnd.n3872 gnd.n1973 19.3944
R9760 gnd.n3882 gnd.n1973 19.3944
R9761 gnd.n3882 gnd.n3881 19.3944
R9762 gnd.n3881 gnd.n3880 19.3944
R9763 gnd.n3880 gnd.n1779 19.3944
R9764 gnd.n4063 gnd.n1779 19.3944
R9765 gnd.n4063 gnd.n1777 19.3944
R9766 gnd.n4067 gnd.n1777 19.3944
R9767 gnd.n4067 gnd.n1767 19.3944
R9768 gnd.n4084 gnd.n1767 19.3944
R9769 gnd.n4084 gnd.n1765 19.3944
R9770 gnd.n4088 gnd.n1765 19.3944
R9771 gnd.n4088 gnd.n1755 19.3944
R9772 gnd.n4107 gnd.n1755 19.3944
R9773 gnd.n4107 gnd.n1753 19.3944
R9774 gnd.n4112 gnd.n1753 19.3944
R9775 gnd.n4112 gnd.n1444 19.3944
R9776 gnd.n4374 gnd.n1444 19.3944
R9777 gnd.n4374 gnd.n4373 19.3944
R9778 gnd.n4373 gnd.n4372 19.3944
R9779 gnd.n4372 gnd.n1448 19.3944
R9780 gnd.n4366 gnd.n1448 19.3944
R9781 gnd.n4366 gnd.n4365 19.3944
R9782 gnd.n4365 gnd.n4364 19.3944
R9783 gnd.n4364 gnd.n1457 19.3944
R9784 gnd.n1575 gnd.n1457 19.3944
R9785 gnd.n1579 gnd.n1575 19.3944
R9786 gnd.n1579 gnd.n1573 19.3944
R9787 gnd.n4188 gnd.n1573 19.3944
R9788 gnd.n4188 gnd.n1571 19.3944
R9789 gnd.n4194 gnd.n1571 19.3944
R9790 gnd.n4194 gnd.n4193 19.3944
R9791 gnd.n4193 gnd.n1546 19.3944
R9792 gnd.n4225 gnd.n1546 19.3944
R9793 gnd.n4225 gnd.n1544 19.3944
R9794 gnd.n4246 gnd.n1544 19.3944
R9795 gnd.n4246 gnd.n4245 19.3944
R9796 gnd.n4245 gnd.n4244 19.3944
R9797 gnd.n4244 gnd.n4231 19.3944
R9798 gnd.n4240 gnd.n4231 19.3944
R9799 gnd.n4240 gnd.n4239 19.3944
R9800 gnd.n4237 gnd.n4235 19.3944
R9801 gnd.n4302 gnd.n4301 19.3944
R9802 gnd.n4306 gnd.n4305 19.3944
R9803 gnd.n7091 gnd.n259 19.3944
R9804 gnd.n7089 gnd.n7088 19.3944
R9805 gnd.n7088 gnd.n261 19.3944
R9806 gnd.n276 gnd.n261 19.3944
R9807 gnd.n277 gnd.n276 19.3944
R9808 gnd.n280 gnd.n277 19.3944
R9809 gnd.n280 gnd.n272 19.3944
R9810 gnd.n7071 gnd.n272 19.3944
R9811 gnd.n7071 gnd.n7070 19.3944
R9812 gnd.n7070 gnd.n7069 19.3944
R9813 gnd.n7069 gnd.n286 19.3944
R9814 gnd.n7044 gnd.n286 19.3944
R9815 gnd.n7044 gnd.n7043 19.3944
R9816 gnd.n7043 gnd.n7042 19.3944
R9817 gnd.n7042 gnd.n292 19.3944
R9818 gnd.n7038 gnd.n292 19.3944
R9819 gnd.n7038 gnd.n7037 19.3944
R9820 gnd.n7037 gnd.n7036 19.3944
R9821 gnd.n7036 gnd.n298 19.3944
R9822 gnd.n300 gnd.n298 19.3944
R9823 gnd.n303 gnd.n300 19.3944
R9824 gnd.n7027 gnd.n303 19.3944
R9825 gnd.n7027 gnd.n7026 19.3944
R9826 gnd.n7026 gnd.n7025 19.3944
R9827 gnd.n7025 gnd.n310 19.3944
R9828 gnd.n7019 gnd.n310 19.3944
R9829 gnd.n7019 gnd.n7018 19.3944
R9830 gnd.n7018 gnd.n7017 19.3944
R9831 gnd.n7017 gnd.n318 19.3944
R9832 gnd.n7011 gnd.n318 19.3944
R9833 gnd.n7011 gnd.n7010 19.3944
R9834 gnd.n4712 gnd.n4711 19.3944
R9835 gnd.n4711 gnd.n4710 19.3944
R9836 gnd.n4710 gnd.n4709 19.3944
R9837 gnd.n4709 gnd.n4707 19.3944
R9838 gnd.n4707 gnd.n4704 19.3944
R9839 gnd.n4704 gnd.n4703 19.3944
R9840 gnd.n4703 gnd.n4700 19.3944
R9841 gnd.n4700 gnd.n4699 19.3944
R9842 gnd.n4699 gnd.n4696 19.3944
R9843 gnd.n4696 gnd.n4695 19.3944
R9844 gnd.n4695 gnd.n4692 19.3944
R9845 gnd.n4692 gnd.n4691 19.3944
R9846 gnd.n4691 gnd.n4688 19.3944
R9847 gnd.n4688 gnd.n4687 19.3944
R9848 gnd.n4687 gnd.n4684 19.3944
R9849 gnd.n4684 gnd.n4683 19.3944
R9850 gnd.n4683 gnd.n4680 19.3944
R9851 gnd.n4678 gnd.n4675 19.3944
R9852 gnd.n4675 gnd.n4674 19.3944
R9853 gnd.n4674 gnd.n4671 19.3944
R9854 gnd.n4671 gnd.n4670 19.3944
R9855 gnd.n4670 gnd.n4667 19.3944
R9856 gnd.n4667 gnd.n4666 19.3944
R9857 gnd.n4666 gnd.n4663 19.3944
R9858 gnd.n4663 gnd.n4662 19.3944
R9859 gnd.n4662 gnd.n4659 19.3944
R9860 gnd.n4659 gnd.n4658 19.3944
R9861 gnd.n4658 gnd.n4655 19.3944
R9862 gnd.n4655 gnd.n4654 19.3944
R9863 gnd.n4654 gnd.n4651 19.3944
R9864 gnd.n4651 gnd.n4650 19.3944
R9865 gnd.n4650 gnd.n4647 19.3944
R9866 gnd.n4647 gnd.n4646 19.3944
R9867 gnd.n4646 gnd.n4643 19.3944
R9868 gnd.n4643 gnd.n4642 19.3944
R9869 gnd.n4633 gnd.n4632 19.3944
R9870 gnd.n4632 gnd.n1125 19.3944
R9871 gnd.n4628 gnd.n1125 19.3944
R9872 gnd.n4628 gnd.n1127 19.3944
R9873 gnd.n4618 gnd.n1127 19.3944
R9874 gnd.n4618 gnd.n4617 19.3944
R9875 gnd.n4617 gnd.n4616 19.3944
R9876 gnd.n4616 gnd.n1150 19.3944
R9877 gnd.n4606 gnd.n1150 19.3944
R9878 gnd.n4606 gnd.n4605 19.3944
R9879 gnd.n4605 gnd.n4604 19.3944
R9880 gnd.n4604 gnd.n1170 19.3944
R9881 gnd.n4594 gnd.n1170 19.3944
R9882 gnd.n4594 gnd.n4593 19.3944
R9883 gnd.n4593 gnd.n4592 19.3944
R9884 gnd.n4592 gnd.n1192 19.3944
R9885 gnd.n1210 gnd.n1192 19.3944
R9886 gnd.n4580 gnd.n1210 19.3944
R9887 gnd.n4580 gnd.n4579 19.3944
R9888 gnd.n4579 gnd.n4578 19.3944
R9889 gnd.n4578 gnd.n1216 19.3944
R9890 gnd.n4567 gnd.n1216 19.3944
R9891 gnd.n4567 gnd.n4566 19.3944
R9892 gnd.n4566 gnd.n4565 19.3944
R9893 gnd.n4565 gnd.n1232 19.3944
R9894 gnd.n4554 gnd.n1232 19.3944
R9895 gnd.n4554 gnd.n4553 19.3944
R9896 gnd.n4553 gnd.n4552 19.3944
R9897 gnd.n4552 gnd.n1251 19.3944
R9898 gnd.n4542 gnd.n1251 19.3944
R9899 gnd.n4542 gnd.n4541 19.3944
R9900 gnd.n4541 gnd.n4540 19.3944
R9901 gnd.n4540 gnd.n1271 19.3944
R9902 gnd.n4530 gnd.n1271 19.3944
R9903 gnd.n4530 gnd.n4529 19.3944
R9904 gnd.n4529 gnd.n4528 19.3944
R9905 gnd.n4528 gnd.n1293 19.3944
R9906 gnd.n4518 gnd.n1293 19.3944
R9907 gnd.n4518 gnd.n4517 19.3944
R9908 gnd.n4517 gnd.n4516 19.3944
R9909 gnd.n4516 gnd.n1314 19.3944
R9910 gnd.n4506 gnd.n1314 19.3944
R9911 gnd.n2687 gnd.n2686 19.3944
R9912 gnd.n2690 gnd.n2687 19.3944
R9913 gnd.n2690 gnd.n2683 19.3944
R9914 gnd.n2696 gnd.n2683 19.3944
R9915 gnd.n2697 gnd.n2696 19.3944
R9916 gnd.n2700 gnd.n2697 19.3944
R9917 gnd.n2700 gnd.n2681 19.3944
R9918 gnd.n2706 gnd.n2681 19.3944
R9919 gnd.n2707 gnd.n2706 19.3944
R9920 gnd.n2710 gnd.n2707 19.3944
R9921 gnd.n2710 gnd.n2679 19.3944
R9922 gnd.n2716 gnd.n2679 19.3944
R9923 gnd.n2717 gnd.n2716 19.3944
R9924 gnd.n2720 gnd.n2717 19.3944
R9925 gnd.n2720 gnd.n2675 19.3944
R9926 gnd.n2724 gnd.n2675 19.3944
R9927 gnd.n2728 gnd.n2670 19.3944
R9928 gnd.n2751 gnd.n2670 19.3944
R9929 gnd.n2751 gnd.n2750 19.3944
R9930 gnd.n2750 gnd.n2749 19.3944
R9931 gnd.n2749 gnd.n2737 19.3944
R9932 gnd.n2737 gnd.n2736 19.3944
R9933 gnd.n2736 gnd.n2651 19.3944
R9934 gnd.n2810 gnd.n2651 19.3944
R9935 gnd.n2810 gnd.n2649 19.3944
R9936 gnd.n2814 gnd.n2649 19.3944
R9937 gnd.n2814 gnd.n2644 19.3944
R9938 gnd.n2827 gnd.n2644 19.3944
R9939 gnd.n2827 gnd.n2642 19.3944
R9940 gnd.n2834 gnd.n2642 19.3944
R9941 gnd.n2834 gnd.n2833 19.3944
R9942 gnd.n2833 gnd.n2614 19.3944
R9943 gnd.n2891 gnd.n2614 19.3944
R9944 gnd.n2891 gnd.n2890 19.3944
R9945 gnd.n2890 gnd.n2889 19.3944
R9946 gnd.n2889 gnd.n2618 19.3944
R9947 gnd.n2852 gnd.n2618 19.3944
R9948 gnd.n2852 gnd.n2630 19.3944
R9949 gnd.n2874 gnd.n2630 19.3944
R9950 gnd.n2874 gnd.n2631 19.3944
R9951 gnd.n2870 gnd.n2631 19.3944
R9952 gnd.n2870 gnd.n2596 19.3944
R9953 gnd.n2909 gnd.n2596 19.3944
R9954 gnd.n2909 gnd.n2594 19.3944
R9955 gnd.n2913 gnd.n2594 19.3944
R9956 gnd.n2913 gnd.n2578 19.3944
R9957 gnd.n2958 gnd.n2578 19.3944
R9958 gnd.n2958 gnd.n2579 19.3944
R9959 gnd.n2954 gnd.n2579 19.3944
R9960 gnd.n2954 gnd.n2953 19.3944
R9961 gnd.n2953 gnd.n2952 19.3944
R9962 gnd.n2952 gnd.n2584 19.3944
R9963 gnd.n2948 gnd.n2584 19.3944
R9964 gnd.n2948 gnd.n2947 19.3944
R9965 gnd.n2947 gnd.n2946 19.3944
R9966 gnd.n2946 gnd.n2494 19.3944
R9967 gnd.n3237 gnd.n2494 19.3944
R9968 gnd.n3237 gnd.n2495 19.3944
R9969 gnd.n2740 gnd.n1118 19.3944
R9970 gnd.n2741 gnd.n2740 19.3944
R9971 gnd.n2741 gnd.n2738 19.3944
R9972 gnd.n2745 gnd.n2738 19.3944
R9973 gnd.n2745 gnd.n2654 19.3944
R9974 gnd.n2802 gnd.n2654 19.3944
R9975 gnd.n2802 gnd.n2652 19.3944
R9976 gnd.n2806 gnd.n2652 19.3944
R9977 gnd.n2806 gnd.n2647 19.3944
R9978 gnd.n2818 gnd.n2647 19.3944
R9979 gnd.n2818 gnd.n2645 19.3944
R9980 gnd.n2823 gnd.n2645 19.3944
R9981 gnd.n2823 gnd.n2641 19.3944
R9982 gnd.n2839 gnd.n2641 19.3944
R9983 gnd.n2840 gnd.n2839 19.3944
R9984 gnd.n2840 gnd.n2639 19.3944
R9985 gnd.n2844 gnd.n2639 19.3944
R9986 gnd.n2845 gnd.n2844 19.3944
R9987 gnd.n2846 gnd.n2845 19.3944
R9988 gnd.n2846 gnd.n2635 19.3944
R9989 gnd.n2856 gnd.n2635 19.3944
R9990 gnd.n2857 gnd.n2856 19.3944
R9991 gnd.n2858 gnd.n2857 19.3944
R9992 gnd.n2858 gnd.n2633 19.3944
R9993 gnd.n2866 gnd.n2633 19.3944
R9994 gnd.n2866 gnd.n2865 19.3944
R9995 gnd.n2865 gnd.n2864 19.3944
R9996 gnd.n2864 gnd.n2593 19.3944
R9997 gnd.n2917 gnd.n2593 19.3944
R9998 gnd.n2917 gnd.n2591 19.3944
R9999 gnd.n2921 gnd.n2591 19.3944
R10000 gnd.n2922 gnd.n2921 19.3944
R10001 gnd.n2925 gnd.n2922 19.3944
R10002 gnd.n2925 gnd.n2589 19.3944
R10003 gnd.n2932 gnd.n2589 19.3944
R10004 gnd.n2933 gnd.n2932 19.3944
R10005 gnd.n2936 gnd.n2933 19.3944
R10006 gnd.n2936 gnd.n2587 19.3944
R10007 gnd.n2941 gnd.n2587 19.3944
R10008 gnd.n2941 gnd.n2493 19.3944
R10009 gnd.n3241 gnd.n2493 19.3944
R10010 gnd.n3242 gnd.n3241 19.3944
R10011 gnd.n3280 gnd.n2396 19.3944
R10012 gnd.n3280 gnd.n2403 19.3944
R10013 gnd.n2460 gnd.n2403 19.3944
R10014 gnd.n3273 gnd.n2460 19.3944
R10015 gnd.n3273 gnd.n3272 19.3944
R10016 gnd.n3272 gnd.n3271 19.3944
R10017 gnd.n3271 gnd.n2466 19.3944
R10018 gnd.n3266 gnd.n2466 19.3944
R10019 gnd.n3266 gnd.n3265 19.3944
R10020 gnd.n3265 gnd.n3264 19.3944
R10021 gnd.n3264 gnd.n2473 19.3944
R10022 gnd.n3259 gnd.n2473 19.3944
R10023 gnd.n3259 gnd.n3258 19.3944
R10024 gnd.n3258 gnd.n3257 19.3944
R10025 gnd.n3257 gnd.n2480 19.3944
R10026 gnd.n3252 gnd.n2480 19.3944
R10027 gnd.n3252 gnd.n3251 19.3944
R10028 gnd.n3251 gnd.n3250 19.3944
R10029 gnd.n2416 gnd.n2415 19.3944
R10030 gnd.n2456 gnd.n2415 19.3944
R10031 gnd.n2456 gnd.n2455 19.3944
R10032 gnd.n2455 gnd.n2454 19.3944
R10033 gnd.n2454 gnd.n2451 19.3944
R10034 gnd.n2451 gnd.n2450 19.3944
R10035 gnd.n2450 gnd.n2447 19.3944
R10036 gnd.n2447 gnd.n2446 19.3944
R10037 gnd.n2446 gnd.n2443 19.3944
R10038 gnd.n2443 gnd.n2442 19.3944
R10039 gnd.n2442 gnd.n2439 19.3944
R10040 gnd.n2439 gnd.n2438 19.3944
R10041 gnd.n2438 gnd.n2435 19.3944
R10042 gnd.n2435 gnd.n2434 19.3944
R10043 gnd.n2434 gnd.n2397 19.3944
R10044 gnd.n2665 gnd.n2661 19.3944
R10045 gnd.n2665 gnd.n1136 19.3944
R10046 gnd.n4624 gnd.n1136 19.3944
R10047 gnd.n4624 gnd.n4623 19.3944
R10048 gnd.n4623 gnd.n4622 19.3944
R10049 gnd.n4622 gnd.n1140 19.3944
R10050 gnd.n4612 gnd.n1140 19.3944
R10051 gnd.n4612 gnd.n4611 19.3944
R10052 gnd.n4611 gnd.n4610 19.3944
R10053 gnd.n4610 gnd.n1160 19.3944
R10054 gnd.n4600 gnd.n1160 19.3944
R10055 gnd.n4600 gnd.n4599 19.3944
R10056 gnd.n4599 gnd.n4598 19.3944
R10057 gnd.n4598 gnd.n1181 19.3944
R10058 gnd.n4588 gnd.n1181 19.3944
R10059 gnd.n4588 gnd.n4587 19.3944
R10060 gnd.n4585 gnd.n4584 19.3944
R10061 gnd.n4574 gnd.n1222 19.3944
R10062 gnd.n4572 gnd.n4571 19.3944
R10063 gnd.n4561 gnd.n1239 19.3944
R10064 gnd.n4559 gnd.n4558 19.3944
R10065 gnd.n4558 gnd.n1240 19.3944
R10066 gnd.n4548 gnd.n1240 19.3944
R10067 gnd.n4548 gnd.n4547 19.3944
R10068 gnd.n4547 gnd.n4546 19.3944
R10069 gnd.n4546 gnd.n1261 19.3944
R10070 gnd.n4536 gnd.n1261 19.3944
R10071 gnd.n4536 gnd.n4535 19.3944
R10072 gnd.n4535 gnd.n4534 19.3944
R10073 gnd.n4534 gnd.n1282 19.3944
R10074 gnd.n4524 gnd.n1282 19.3944
R10075 gnd.n4524 gnd.n4523 19.3944
R10076 gnd.n4523 gnd.n4522 19.3944
R10077 gnd.n4522 gnd.n1303 19.3944
R10078 gnd.n4512 gnd.n1303 19.3944
R10079 gnd.n4512 gnd.n4511 19.3944
R10080 gnd.n4511 gnd.n4510 19.3944
R10081 gnd.n6270 gnd.n765 19.3944
R10082 gnd.n6270 gnd.n6269 19.3944
R10083 gnd.n6269 gnd.n6268 19.3944
R10084 gnd.n6268 gnd.n769 19.3944
R10085 gnd.n6262 gnd.n769 19.3944
R10086 gnd.n6262 gnd.n6261 19.3944
R10087 gnd.n6261 gnd.n6260 19.3944
R10088 gnd.n6260 gnd.n777 19.3944
R10089 gnd.n6254 gnd.n777 19.3944
R10090 gnd.n6254 gnd.n6253 19.3944
R10091 gnd.n6253 gnd.n6252 19.3944
R10092 gnd.n6252 gnd.n785 19.3944
R10093 gnd.n6246 gnd.n785 19.3944
R10094 gnd.n6246 gnd.n6245 19.3944
R10095 gnd.n6245 gnd.n6244 19.3944
R10096 gnd.n6244 gnd.n793 19.3944
R10097 gnd.n6238 gnd.n793 19.3944
R10098 gnd.n6238 gnd.n6237 19.3944
R10099 gnd.n6237 gnd.n6236 19.3944
R10100 gnd.n6236 gnd.n801 19.3944
R10101 gnd.n6230 gnd.n801 19.3944
R10102 gnd.n6230 gnd.n6229 19.3944
R10103 gnd.n6229 gnd.n6228 19.3944
R10104 gnd.n6228 gnd.n809 19.3944
R10105 gnd.n6222 gnd.n809 19.3944
R10106 gnd.n6222 gnd.n6221 19.3944
R10107 gnd.n6221 gnd.n6220 19.3944
R10108 gnd.n6220 gnd.n817 19.3944
R10109 gnd.n6214 gnd.n817 19.3944
R10110 gnd.n6214 gnd.n6213 19.3944
R10111 gnd.n6213 gnd.n6212 19.3944
R10112 gnd.n6212 gnd.n825 19.3944
R10113 gnd.n6206 gnd.n825 19.3944
R10114 gnd.n6206 gnd.n6205 19.3944
R10115 gnd.n6205 gnd.n6204 19.3944
R10116 gnd.n6204 gnd.n833 19.3944
R10117 gnd.n6198 gnd.n833 19.3944
R10118 gnd.n6198 gnd.n6197 19.3944
R10119 gnd.n6197 gnd.n6196 19.3944
R10120 gnd.n6196 gnd.n841 19.3944
R10121 gnd.n6190 gnd.n841 19.3944
R10122 gnd.n6190 gnd.n6189 19.3944
R10123 gnd.n6189 gnd.n6188 19.3944
R10124 gnd.n6188 gnd.n849 19.3944
R10125 gnd.n6182 gnd.n849 19.3944
R10126 gnd.n6182 gnd.n6181 19.3944
R10127 gnd.n6181 gnd.n6180 19.3944
R10128 gnd.n6180 gnd.n857 19.3944
R10129 gnd.n6174 gnd.n857 19.3944
R10130 gnd.n6174 gnd.n6173 19.3944
R10131 gnd.n6173 gnd.n6172 19.3944
R10132 gnd.n6172 gnd.n865 19.3944
R10133 gnd.n6166 gnd.n865 19.3944
R10134 gnd.n6166 gnd.n6165 19.3944
R10135 gnd.n6165 gnd.n6164 19.3944
R10136 gnd.n6164 gnd.n873 19.3944
R10137 gnd.n6158 gnd.n873 19.3944
R10138 gnd.n6158 gnd.n6157 19.3944
R10139 gnd.n6157 gnd.n6156 19.3944
R10140 gnd.n6156 gnd.n881 19.3944
R10141 gnd.n6150 gnd.n881 19.3944
R10142 gnd.n6150 gnd.n6149 19.3944
R10143 gnd.n6149 gnd.n6148 19.3944
R10144 gnd.n6148 gnd.n889 19.3944
R10145 gnd.n6142 gnd.n889 19.3944
R10146 gnd.n6142 gnd.n6141 19.3944
R10147 gnd.n6141 gnd.n6140 19.3944
R10148 gnd.n6140 gnd.n897 19.3944
R10149 gnd.n6134 gnd.n897 19.3944
R10150 gnd.n6134 gnd.n6133 19.3944
R10151 gnd.n6133 gnd.n6132 19.3944
R10152 gnd.n6132 gnd.n905 19.3944
R10153 gnd.n6126 gnd.n905 19.3944
R10154 gnd.n6126 gnd.n6125 19.3944
R10155 gnd.n6125 gnd.n6124 19.3944
R10156 gnd.n6124 gnd.n913 19.3944
R10157 gnd.n6118 gnd.n913 19.3944
R10158 gnd.n6118 gnd.n6117 19.3944
R10159 gnd.n6117 gnd.n6116 19.3944
R10160 gnd.n6116 gnd.n921 19.3944
R10161 gnd.n6110 gnd.n921 19.3944
R10162 gnd.n6110 gnd.n6109 19.3944
R10163 gnd.n6109 gnd.n6108 19.3944
R10164 gnd.n6108 gnd.n929 19.3944
R10165 gnd.n4501 gnd.n4500 19.3944
R10166 gnd.n4500 gnd.n4499 19.3944
R10167 gnd.n4499 gnd.n1338 19.3944
R10168 gnd.n4495 gnd.n1338 19.3944
R10169 gnd.n4495 gnd.n4494 19.3944
R10170 gnd.n4494 gnd.n4493 19.3944
R10171 gnd.n4493 gnd.n1343 19.3944
R10172 gnd.n4489 gnd.n1343 19.3944
R10173 gnd.n4489 gnd.n4488 19.3944
R10174 gnd.n4488 gnd.n4487 19.3944
R10175 gnd.n4487 gnd.n1348 19.3944
R10176 gnd.n4483 gnd.n1348 19.3944
R10177 gnd.n4483 gnd.n4482 19.3944
R10178 gnd.n4482 gnd.n4481 19.3944
R10179 gnd.n4481 gnd.n1353 19.3944
R10180 gnd.n4477 gnd.n1353 19.3944
R10181 gnd.n4477 gnd.n4476 19.3944
R10182 gnd.n4476 gnd.n4475 19.3944
R10183 gnd.n4475 gnd.n1358 19.3944
R10184 gnd.n4471 gnd.n1358 19.3944
R10185 gnd.n4471 gnd.n4470 19.3944
R10186 gnd.n4470 gnd.n4469 19.3944
R10187 gnd.n4469 gnd.n1363 19.3944
R10188 gnd.n4465 gnd.n1363 19.3944
R10189 gnd.n4465 gnd.n4464 19.3944
R10190 gnd.n4464 gnd.n4463 19.3944
R10191 gnd.n4463 gnd.n1368 19.3944
R10192 gnd.n4459 gnd.n1368 19.3944
R10193 gnd.n4459 gnd.n4458 19.3944
R10194 gnd.n4458 gnd.n4457 19.3944
R10195 gnd.n4457 gnd.n1373 19.3944
R10196 gnd.n4453 gnd.n1373 19.3944
R10197 gnd.n4453 gnd.n4452 19.3944
R10198 gnd.n4452 gnd.n4451 19.3944
R10199 gnd.n4451 gnd.n1378 19.3944
R10200 gnd.n4447 gnd.n1378 19.3944
R10201 gnd.n4447 gnd.n4446 19.3944
R10202 gnd.n4446 gnd.n4445 19.3944
R10203 gnd.n4445 gnd.n1383 19.3944
R10204 gnd.n4441 gnd.n1383 19.3944
R10205 gnd.n4441 gnd.n4440 19.3944
R10206 gnd.n4440 gnd.n4439 19.3944
R10207 gnd.n4439 gnd.n1388 19.3944
R10208 gnd.n4435 gnd.n1388 19.3944
R10209 gnd.n4435 gnd.n4434 19.3944
R10210 gnd.n4434 gnd.n4433 19.3944
R10211 gnd.n4433 gnd.n1393 19.3944
R10212 gnd.n4429 gnd.n1393 19.3944
R10213 gnd.n4429 gnd.n4428 19.3944
R10214 gnd.n4428 gnd.n4427 19.3944
R10215 gnd.n4427 gnd.n1398 19.3944
R10216 gnd.n4423 gnd.n1398 19.3944
R10217 gnd.n4423 gnd.n4422 19.3944
R10218 gnd.n4422 gnd.n4421 19.3944
R10219 gnd.n4421 gnd.n1403 19.3944
R10220 gnd.n4417 gnd.n1403 19.3944
R10221 gnd.n4417 gnd.n4416 19.3944
R10222 gnd.n4416 gnd.n4415 19.3944
R10223 gnd.n4415 gnd.n1408 19.3944
R10224 gnd.n4411 gnd.n1408 19.3944
R10225 gnd.n4411 gnd.n4410 19.3944
R10226 gnd.n4410 gnd.n4409 19.3944
R10227 gnd.n4409 gnd.n1413 19.3944
R10228 gnd.n4405 gnd.n1413 19.3944
R10229 gnd.n4405 gnd.n4404 19.3944
R10230 gnd.n4404 gnd.n4403 19.3944
R10231 gnd.n4403 gnd.n1418 19.3944
R10232 gnd.n4399 gnd.n1418 19.3944
R10233 gnd.n4399 gnd.n4398 19.3944
R10234 gnd.n4398 gnd.n4397 19.3944
R10235 gnd.n4397 gnd.n1423 19.3944
R10236 gnd.n4393 gnd.n1423 19.3944
R10237 gnd.n4393 gnd.n4392 19.3944
R10238 gnd.n4392 gnd.n4391 19.3944
R10239 gnd.n4391 gnd.n1428 19.3944
R10240 gnd.n4387 gnd.n1428 19.3944
R10241 gnd.n4387 gnd.n4386 19.3944
R10242 gnd.n4386 gnd.n4385 19.3944
R10243 gnd.n4385 gnd.n1433 19.3944
R10244 gnd.n4381 gnd.n1433 19.3944
R10245 gnd.n4381 gnd.n4380 19.3944
R10246 gnd.n4380 gnd.n4379 19.3944
R10247 gnd.n4130 gnd.n1748 19.3944
R10248 gnd.n4126 gnd.n1748 19.3944
R10249 gnd.n4126 gnd.n4125 19.3944
R10250 gnd.n1658 gnd.n1640 19.3944
R10251 gnd.n1658 gnd.n1638 19.3944
R10252 gnd.n1664 gnd.n1638 19.3944
R10253 gnd.n1664 gnd.n1631 19.3944
R10254 gnd.n1677 gnd.n1631 19.3944
R10255 gnd.n1677 gnd.n1629 19.3944
R10256 gnd.n1683 gnd.n1629 19.3944
R10257 gnd.n1683 gnd.n1622 19.3944
R10258 gnd.n1696 gnd.n1622 19.3944
R10259 gnd.n1696 gnd.n1620 19.3944
R10260 gnd.n1702 gnd.n1620 19.3944
R10261 gnd.n1702 gnd.n1613 19.3944
R10262 gnd.n1715 gnd.n1613 19.3944
R10263 gnd.n1715 gnd.n1611 19.3944
R10264 gnd.n1721 gnd.n1611 19.3944
R10265 gnd.n1721 gnd.n1602 19.3944
R10266 gnd.n1732 gnd.n1602 19.3944
R10267 gnd.n1732 gnd.n1600 19.3944
R10268 gnd.n4141 gnd.n1600 19.3944
R10269 gnd.n4141 gnd.n4140 19.3944
R10270 gnd.n4140 gnd.n4139 19.3944
R10271 gnd.n4139 gnd.n1740 19.3944
R10272 gnd.n4135 gnd.n1740 19.3944
R10273 gnd.n4135 gnd.n4134 19.3944
R10274 gnd.n5505 gnd.t17 18.8012
R10275 gnd.n5490 gnd.t0 18.8012
R10276 gnd.n5349 gnd.n5348 18.4825
R10277 gnd.n1957 gnd.n1822 18.4247
R10278 gnd.n3284 gnd.n2397 18.4247
R10279 gnd.n7217 gnd.n7216 18.2308
R10280 gnd.n1724 gnd.n1606 18.2308
R10281 gnd.n3087 gnd.n3071 18.2308
R10282 gnd.n2725 gnd.n2724 18.2308
R10283 gnd.t9 gnd.n5029 18.1639
R10284 gnd.n6105 gnd.n6104 18.1639
R10285 gnd.n5057 gnd.t16 17.5266
R10286 gnd.n5456 gnd.t13 16.8893
R10287 gnd.n3239 gnd.t64 16.8893
R10288 gnd.n4148 gnd.t46 16.8893
R10289 gnd.n5284 gnd.t123 16.2519
R10290 gnd.n4984 gnd.t11 16.2519
R10291 gnd.n3128 gnd.n3127 15.9333
R10292 gnd.n3127 gnd.n2553 15.9333
R10293 gnd.n3137 gnd.n3136 15.9333
R10294 gnd.n3138 gnd.n3137 15.9333
R10295 gnd.n3139 gnd.n3138 15.9333
R10296 gnd.n3142 gnd.n3139 15.9333
R10297 gnd.n3141 gnd.n3140 15.9333
R10298 gnd.n3140 gnd.n2547 15.9333
R10299 gnd.n3150 gnd.n2547 15.9333
R10300 gnd.n3151 gnd.n3150 15.9333
R10301 gnd.n3152 gnd.n3151 15.9333
R10302 gnd.n3153 gnd.n3152 15.9333
R10303 gnd.n3156 gnd.n3153 15.9333
R10304 gnd.n3156 gnd.n3155 15.9333
R10305 gnd.n3154 gnd.n2539 15.9333
R10306 gnd.n3164 gnd.n2539 15.9333
R10307 gnd.n3165 gnd.n3164 15.9333
R10308 gnd.n3166 gnd.n3165 15.9333
R10309 gnd.n3167 gnd.n3166 15.9333
R10310 gnd.n3170 gnd.n3167 15.9333
R10311 gnd.n3170 gnd.n3169 15.9333
R10312 gnd.n3169 gnd.n3168 15.9333
R10313 gnd.n3180 gnd.n3178 15.9333
R10314 gnd.n3178 gnd.n2289 15.9333
R10315 gnd.n3183 gnd.n2322 15.9333
R10316 gnd.n3359 gnd.n3358 15.9333
R10317 gnd.n3367 gnd.n2254 15.9333
R10318 gnd.n3450 gnd.n2242 15.9333
R10319 gnd.n3460 gnd.n3458 15.9333
R10320 gnd.n3491 gnd.n3489 15.9333
R10321 gnd.n3411 gnd.n2191 15.9333
R10322 gnd.n3546 gnd.n3545 15.9333
R10323 gnd.n3555 gnd.n3554 15.9333
R10324 gnd.n3554 gnd.n2153 15.9333
R10325 gnd.n3382 gnd.n2124 15.9333
R10326 gnd.n3374 gnd.n2120 15.9333
R10327 gnd.n3633 gnd.n2112 15.9333
R10328 gnd.n3655 gnd.n3654 15.9333
R10329 gnd.n3686 gnd.n2068 15.9333
R10330 gnd.n3686 gnd.n3685 15.9333
R10331 gnd.n3715 gnd.n2051 15.9333
R10332 gnd.n3755 gnd.n2028 15.9333
R10333 gnd.n3794 gnd.n3792 15.9333
R10334 gnd.n3835 gnd.n3833 15.9333
R10335 gnd.n3870 gnd.n3869 15.9333
R10336 gnd.n4050 gnd.n4049 15.9333
R10337 gnd.n4061 gnd.n4060 15.9333
R10338 gnd.n4058 gnd.n1775 15.9333
R10339 gnd.n4069 gnd.n1775 15.9333
R10340 gnd.n4071 gnd.n4069 15.9333
R10341 gnd.n4071 gnd.n4070 15.9333
R10342 gnd.n4070 gnd.n1769 15.9333
R10343 gnd.n4082 gnd.n1769 15.9333
R10344 gnd.n4082 gnd.n4081 15.9333
R10345 gnd.n4081 gnd.n4079 15.9333
R10346 gnd.n4090 gnd.n1763 15.9333
R10347 gnd.n4092 gnd.n4090 15.9333
R10348 gnd.n4092 gnd.n4091 15.9333
R10349 gnd.n4091 gnd.n1757 15.9333
R10350 gnd.n4105 gnd.n1757 15.9333
R10351 gnd.n4105 gnd.n4104 15.9333
R10352 gnd.n4104 gnd.n4102 15.9333
R10353 gnd.n4102 gnd.n4101 15.9333
R10354 gnd.n4115 gnd.n4114 15.9333
R10355 gnd.n4115 gnd.n1439 15.9333
R10356 gnd.n4377 gnd.n1439 15.9333
R10357 gnd.n4377 gnd.n4376 15.9333
R10358 gnd.n1450 gnd.n1441 15.9333
R10359 gnd.n4370 gnd.n1450 15.9333
R10360 gnd.n5901 gnd.n5899 15.6674
R10361 gnd.n5869 gnd.n5867 15.6674
R10362 gnd.n5837 gnd.n5835 15.6674
R10363 gnd.n5806 gnd.n5804 15.6674
R10364 gnd.n5774 gnd.n5772 15.6674
R10365 gnd.n5742 gnd.n5740 15.6674
R10366 gnd.n5710 gnd.n5708 15.6674
R10367 gnd.n5679 gnd.n5677 15.6674
R10368 gnd.n5275 gnd.t123 15.6146
R10369 gnd.t36 gnd.n6062 15.6146
R10370 gnd.n5966 gnd.t90 15.6146
R10371 gnd.t97 gnd.n3141 15.6146
R10372 gnd.n4101 gnd.t74 15.6146
R10373 gnd.n3421 gnd.n2214 15.296
R10374 gnd.n3509 gnd.n2199 15.296
R10375 gnd.n3625 gnd.n3624 15.296
R10376 gnd.n2111 gnd.n2102 15.296
R10377 gnd.n3784 gnd.n3783 15.296
R10378 gnd.n3795 gnd.n2007 15.296
R10379 gnd.n3892 gnd.n3891 15.0827
R10380 gnd.n2275 gnd.n2270 15.0481
R10381 gnd.n3902 gnd.n3901 15.0481
R10382 gnd.n6097 gnd.t20 14.9773
R10383 gnd.t116 gnd.n2753 14.9773
R10384 gnd.n3168 gnd.t270 14.9773
R10385 gnd.t171 gnd.n4058 14.9773
R10386 gnd.n173 gnd.t32 14.9773
R10387 gnd.n3449 gnd.n2244 14.6587
R10388 gnd.n3468 gnd.t2 14.6587
R10389 gnd.n3535 gnd.n2170 14.6587
R10390 gnd.n3573 gnd.n2149 14.6587
R10391 gnd.n3695 gnd.n2074 14.6587
R10392 gnd.n3735 gnd.n3734 14.6587
R10393 gnd.t5 gnd.n3824 14.6587
R10394 gnd.n3861 gnd.n1977 14.6587
R10395 gnd.n4050 gnd.n1786 14.6587
R10396 gnd.n4061 gnd.t113 14.6587
R10397 gnd.n6083 gnd.t23 14.34
R10398 gnd.t14 gnd.n980 14.34
R10399 gnd.n3470 gnd.n3469 14.0214
R10400 gnd.n3520 gnd.n3519 14.0214
R10401 gnd.n3383 gnd.n2135 14.0214
R10402 gnd.n3653 gnd.n2088 14.0214
R10403 gnd.n3756 gnd.n3753 14.0214
R10404 gnd.n3823 gnd.n2002 14.0214
R10405 gnd.n5431 gnd.t145 13.7027
R10406 gnd.n3574 gnd.t159 13.7027
R10407 gnd.n3694 gnd.t161 13.7027
R10408 gnd.n5141 gnd.n5140 13.5763
R10409 gnd.n6022 gnd.n4773 13.5763
R10410 gnd.n1918 gnd.n1910 13.5763
R10411 gnd.n7255 gnd.n7254 13.5763
R10412 gnd.n4642 gnd.n1115 13.5763
R10413 gnd.n3250 gnd.n2489 13.5763
R10414 gnd.n5349 gnd.n5087 13.384
R10415 gnd.n3527 gnd.n3526 13.384
R10416 gnd.n3593 gnd.n2133 13.384
R10417 gnd.n3667 gnd.n3666 13.384
R10418 gnd.n3726 gnd.n3725 13.384
R10419 gnd.n3805 gnd.n1993 13.384
R10420 gnd.n2286 gnd.n2267 13.1884
R10421 gnd.n2281 gnd.n2280 13.1884
R10422 gnd.n2280 gnd.n2279 13.1884
R10423 gnd.n3895 gnd.n3890 13.1884
R10424 gnd.n3896 gnd.n3895 13.1884
R10425 gnd.n2282 gnd.n2269 13.146
R10426 gnd.n2278 gnd.n2269 13.146
R10427 gnd.n3894 gnd.n3893 13.146
R10428 gnd.n3894 gnd.n3889 13.146
R10429 gnd.t140 gnd.n2249 13.0654
R10430 gnd.n3848 gnd.t137 13.0654
R10431 gnd.n5902 gnd.n5898 12.8005
R10432 gnd.n5870 gnd.n5866 12.8005
R10433 gnd.n5838 gnd.n5834 12.8005
R10434 gnd.n5807 gnd.n5803 12.8005
R10435 gnd.n5775 gnd.n5771 12.8005
R10436 gnd.n5743 gnd.n5739 12.8005
R10437 gnd.n5711 gnd.n5707 12.8005
R10438 gnd.n5680 gnd.n5676 12.8005
R10439 gnd.n3431 gnd.n2234 12.7467
R10440 gnd.n3586 gnd.n2139 12.7467
R10441 gnd.n3674 gnd.n2084 12.7467
R10442 gnd.n3348 gnd.n2322 12.4281
R10443 gnd.n4049 gnd.n4048 12.4281
R10444 gnd.n5140 gnd.n5135 12.4126
R10445 gnd.n6027 gnd.n4773 12.4126
R10446 gnd.n1914 gnd.n1910 12.4126
R10447 gnd.n7254 gnd.n156 12.4126
R10448 gnd.n4638 gnd.n1115 12.4126
R10449 gnd.n3245 gnd.n2489 12.4126
R10450 gnd.n3352 gnd.n3351 12.1761
R10451 gnd.n3975 gnd.n3974 12.1761
R10452 gnd.n3480 gnd.n2222 12.1094
R10453 gnd.t156 gnd.n2201 12.1094
R10454 gnd.t173 gnd.n3774 12.1094
R10455 gnd.n3813 gnd.n1999 12.1094
R10456 gnd.t40 gnd.n1965 12.1094
R10457 gnd.n5906 gnd.n5905 12.0247
R10458 gnd.n5874 gnd.n5873 12.0247
R10459 gnd.n5842 gnd.n5841 12.0247
R10460 gnd.n5811 gnd.n5810 12.0247
R10461 gnd.n5779 gnd.n5778 12.0247
R10462 gnd.n5747 gnd.n5746 12.0247
R10463 gnd.n5715 gnd.n5714 12.0247
R10464 gnd.n5684 gnd.n5683 12.0247
R10465 gnd.n4526 gnd.t176 11.7908
R10466 gnd.n4197 gnd.t228 11.7908
R10467 gnd.n2993 gnd.n2459 11.4721
R10468 gnd.t43 gnd.n2260 11.4721
R10469 gnd.n3357 gnd.n2263 11.4721
R10470 gnd.n3979 gnd.n1964 11.4721
R10471 gnd.n4368 gnd.n1451 11.4721
R10472 gnd.n5909 gnd.n5896 11.249
R10473 gnd.n5877 gnd.n5864 11.249
R10474 gnd.n5845 gnd.n5832 11.249
R10475 gnd.n5814 gnd.n5801 11.249
R10476 gnd.n5782 gnd.n5769 11.249
R10477 gnd.n5750 gnd.n5737 11.249
R10478 gnd.n5718 gnd.n5705 11.249
R10479 gnd.n5687 gnd.n5674 11.249
R10480 gnd.n5419 gnd.t145 11.1535
R10481 gnd.t197 gnd.n1175 11.1535
R10482 gnd.n4550 gnd.t174 11.1535
R10483 gnd.n3155 gnd.t272 11.1535
R10484 gnd.n3404 gnd.t151 11.1535
R10485 gnd.t280 gnd.n3744 11.1535
R10486 gnd.t147 gnd.n1763 11.1535
R10487 gnd.n1532 gnd.t180 11.1535
R10488 gnd.t192 gnd.n203 11.1535
R10489 gnd.n4635 gnd.n1121 10.8348
R10490 gnd.n2754 gnd.n2667 10.8348
R10491 gnd.n2753 gnd.n1130 10.8348
R10492 gnd.n4626 gnd.n1133 10.8348
R10493 gnd.n2747 gnd.n1142 10.8348
R10494 gnd.n4620 gnd.n1145 10.8348
R10495 gnd.n2800 gnd.n2799 10.8348
R10496 gnd.n4614 gnd.n1154 10.8348
R10497 gnd.n2808 gnd.n1162 10.8348
R10498 gnd.n2816 gnd.n1172 10.8348
R10499 gnd.n4602 gnd.n1175 10.8348
R10500 gnd.n2825 gnd.n1183 10.8348
R10501 gnd.n4596 gnd.n1186 10.8348
R10502 gnd.n2837 gnd.n2836 10.8348
R10503 gnd.n4590 gnd.n1196 10.8348
R10504 gnd.n2894 gnd.n2611 10.8348
R10505 gnd.n4582 gnd.n1207 10.8348
R10506 gnd.n2887 gnd.n2886 10.8348
R10507 gnd.n4576 gnd.n1220 10.8348
R10508 gnd.n2854 gnd.n1225 10.8348
R10509 gnd.n2876 gnd.n1234 10.8348
R10510 gnd.n4563 gnd.n1237 10.8348
R10511 gnd.n2868 gnd.n1242 10.8348
R10512 gnd.n4556 gnd.n1245 10.8348
R10513 gnd.n2907 gnd.n2906 10.8348
R10514 gnd.n4550 gnd.n1255 10.8348
R10515 gnd.n2915 gnd.n1263 10.8348
R10516 gnd.n2960 gnd.n1273 10.8348
R10517 gnd.n4538 gnd.n1276 10.8348
R10518 gnd.n2923 gnd.n1284 10.8348
R10519 gnd.n4532 gnd.n1287 10.8348
R10520 gnd.n2930 gnd.n2929 10.8348
R10521 gnd.n4526 gnd.n1297 10.8348
R10522 gnd.n2934 gnd.n1305 10.8348
R10523 gnd.n4520 gnd.n1308 10.8348
R10524 gnd.n2943 gnd.n1316 10.8348
R10525 gnd.n4514 gnd.n1319 10.8348
R10526 gnd.n3239 gnd.n1326 10.8348
R10527 gnd.n4508 gnd.n1329 10.8348
R10528 gnd.n3502 gnd.n2205 10.8348
R10529 gnd.t155 gnd.n2186 10.8348
R10530 gnd.n3375 gnd.n2109 10.8348
R10531 gnd.n3634 gnd.n2109 10.8348
R10532 gnd.n2058 gnd.t3 10.8348
R10533 gnd.n3766 gnd.n3765 10.8348
R10534 gnd.n4362 gnd.n4361 10.8348
R10535 gnd.n4148 gnd.n1462 10.8348
R10536 gnd.n4355 gnd.n1471 10.8348
R10537 gnd.n4176 gnd.n1474 10.8348
R10538 gnd.n4175 gnd.n1586 10.8348
R10539 gnd.n4186 gnd.n4185 10.8348
R10540 gnd.n4197 gnd.n1564 10.8348
R10541 gnd.n4196 gnd.n1568 10.8348
R10542 gnd.n4207 gnd.n1555 10.8348
R10543 gnd.n4164 gnd.n1557 10.8348
R10544 gnd.n4223 gnd.n4222 10.8348
R10545 gnd.n4250 gnd.n1539 10.8348
R10546 gnd.n4260 gnd.n1530 10.8348
R10547 gnd.n1533 gnd.n1532 10.8348
R10548 gnd.n4326 gnd.n1502 10.8348
R10549 gnd.n4329 gnd.n1496 10.8348
R10550 gnd.n4268 gnd.n1499 10.8348
R10551 gnd.n7113 gnd.n233 10.8348
R10552 gnd.n4298 gnd.n236 10.8348
R10553 gnd.n4309 gnd.n1513 10.8348
R10554 gnd.n4308 gnd.n1518 10.8348
R10555 gnd.n4290 gnd.n4288 10.8348
R10556 gnd.n7094 gnd.n255 10.8348
R10557 gnd.n4282 gnd.n251 10.8348
R10558 gnd.n7122 gnd.n220 10.8348
R10559 gnd.n7085 gnd.n7084 10.8348
R10560 gnd.n7130 gnd.n211 10.8348
R10561 gnd.n7078 gnd.n214 10.8348
R10562 gnd.n7138 gnd.n203 10.8348
R10563 gnd.n7074 gnd.n205 10.8348
R10564 gnd.n7048 gnd.n197 10.8348
R10565 gnd.n7154 gnd.n188 10.8348
R10566 gnd.n7066 gnd.n7065 10.8348
R10567 gnd.n7162 gnd.n179 10.8348
R10568 gnd.n7059 gnd.n182 10.8348
R10569 gnd.n7172 gnd.n169 10.8348
R10570 gnd.n173 gnd.n171 10.8348
R10571 gnd.n7247 gnd.n162 10.8348
R10572 gnd.n7326 gnd.n81 10.8348
R10573 gnd.n4045 gnd.n4044 10.6151
R10574 gnd.n4044 gnd.n4041 10.6151
R10575 gnd.n4039 gnd.n4036 10.6151
R10576 gnd.n4036 gnd.n4035 10.6151
R10577 gnd.n4035 gnd.n4032 10.6151
R10578 gnd.n4032 gnd.n4031 10.6151
R10579 gnd.n4031 gnd.n4028 10.6151
R10580 gnd.n4028 gnd.n4027 10.6151
R10581 gnd.n4027 gnd.n4024 10.6151
R10582 gnd.n4024 gnd.n4023 10.6151
R10583 gnd.n4023 gnd.n4020 10.6151
R10584 gnd.n4020 gnd.n4019 10.6151
R10585 gnd.n4019 gnd.n4016 10.6151
R10586 gnd.n4016 gnd.n4015 10.6151
R10587 gnd.n4015 gnd.n4012 10.6151
R10588 gnd.n4012 gnd.n4011 10.6151
R10589 gnd.n4011 gnd.n4008 10.6151
R10590 gnd.n4008 gnd.n4007 10.6151
R10591 gnd.n4007 gnd.n4004 10.6151
R10592 gnd.n4004 gnd.n4003 10.6151
R10593 gnd.n4003 gnd.n4000 10.6151
R10594 gnd.n4000 gnd.n3999 10.6151
R10595 gnd.n3999 gnd.n3996 10.6151
R10596 gnd.n3996 gnd.n3995 10.6151
R10597 gnd.n3995 gnd.n3992 10.6151
R10598 gnd.n3992 gnd.n3991 10.6151
R10599 gnd.n3991 gnd.n3988 10.6151
R10600 gnd.n3988 gnd.n3987 10.6151
R10601 gnd.n3987 gnd.n3984 10.6151
R10602 gnd.n3984 gnd.n3983 10.6151
R10603 gnd.n2330 gnd.n2329 10.6151
R10604 gnd.n2329 gnd.n2251 10.6151
R10605 gnd.n3369 gnd.n2251 10.6151
R10606 gnd.n3370 gnd.n3369 10.6151
R10607 gnd.n3436 gnd.n3370 10.6151
R10608 gnd.n3436 gnd.n3435 10.6151
R10609 gnd.n3435 gnd.n3434 10.6151
R10610 gnd.n3434 gnd.n3371 10.6151
R10611 gnd.n3428 gnd.n3371 10.6151
R10612 gnd.n3428 gnd.n3427 10.6151
R10613 gnd.n3427 gnd.n3426 10.6151
R10614 gnd.n3426 gnd.n3425 10.6151
R10615 gnd.n3425 gnd.n3424 10.6151
R10616 gnd.n3424 gnd.n3372 10.6151
R10617 gnd.n3418 gnd.n3372 10.6151
R10618 gnd.n3418 gnd.n3417 10.6151
R10619 gnd.n3417 gnd.n3416 10.6151
R10620 gnd.n3416 gnd.n3414 10.6151
R10621 gnd.n3414 gnd.n3413 10.6151
R10622 gnd.n3413 gnd.n3410 10.6151
R10623 gnd.n3410 gnd.n3409 10.6151
R10624 gnd.n3409 gnd.n3407 10.6151
R10625 gnd.n3407 gnd.n3406 10.6151
R10626 gnd.n3406 gnd.n3402 10.6151
R10627 gnd.n3402 gnd.n3401 10.6151
R10628 gnd.n3401 gnd.n3399 10.6151
R10629 gnd.n3399 gnd.n3398 10.6151
R10630 gnd.n3398 gnd.n3396 10.6151
R10631 gnd.n3396 gnd.n3395 10.6151
R10632 gnd.n3395 gnd.n3394 10.6151
R10633 gnd.n3394 gnd.n3393 10.6151
R10634 gnd.n3393 gnd.n3392 10.6151
R10635 gnd.n3392 gnd.n3389 10.6151
R10636 gnd.n3389 gnd.n3388 10.6151
R10637 gnd.n3388 gnd.n3386 10.6151
R10638 gnd.n3386 gnd.n3385 10.6151
R10639 gnd.n3385 gnd.n3381 10.6151
R10640 gnd.n3381 gnd.n3380 10.6151
R10641 gnd.n3380 gnd.n3378 10.6151
R10642 gnd.n3378 gnd.n3377 10.6151
R10643 gnd.n3377 gnd.n3373 10.6151
R10644 gnd.n3373 gnd.n2100 10.6151
R10645 gnd.n3643 gnd.n2100 10.6151
R10646 gnd.n3644 gnd.n3643 10.6151
R10647 gnd.n3651 gnd.n3644 10.6151
R10648 gnd.n3651 gnd.n3650 10.6151
R10649 gnd.n3650 gnd.n3649 10.6151
R10650 gnd.n3649 gnd.n3648 10.6151
R10651 gnd.n3648 gnd.n3647 10.6151
R10652 gnd.n3647 gnd.n2077 10.6151
R10653 gnd.n3690 gnd.n2077 10.6151
R10654 gnd.n3690 gnd.n3689 10.6151
R10655 gnd.n3689 gnd.n3688 10.6151
R10656 gnd.n3688 gnd.n2059 10.6151
R10657 gnd.n3718 gnd.n2059 10.6151
R10658 gnd.n3719 gnd.n3718 10.6151
R10659 gnd.n3721 gnd.n3719 10.6151
R10660 gnd.n3722 gnd.n3721 10.6151
R10661 gnd.n3723 gnd.n3722 10.6151
R10662 gnd.n3723 gnd.n2036 10.6151
R10663 gnd.n3758 gnd.n2036 10.6151
R10664 gnd.n3759 gnd.n3758 10.6151
R10665 gnd.n3761 gnd.n3759 10.6151
R10666 gnd.n3762 gnd.n3761 10.6151
R10667 gnd.n3763 gnd.n3762 10.6151
R10668 gnd.n3763 gnd.n2013 10.6151
R10669 gnd.n3797 gnd.n2013 10.6151
R10670 gnd.n3798 gnd.n3797 10.6151
R10671 gnd.n3800 gnd.n3798 10.6151
R10672 gnd.n3801 gnd.n3800 10.6151
R10673 gnd.n3802 gnd.n3801 10.6151
R10674 gnd.n3802 gnd.n1991 10.6151
R10675 gnd.n3838 gnd.n1991 10.6151
R10676 gnd.n3839 gnd.n3838 10.6151
R10677 gnd.n3841 gnd.n3839 10.6151
R10678 gnd.n3842 gnd.n3841 10.6151
R10679 gnd.n3845 gnd.n3842 10.6151
R10680 gnd.n3845 gnd.n3844 10.6151
R10681 gnd.n3844 gnd.n3843 10.6151
R10682 gnd.n3843 gnd.n1963 10.6151
R10683 gnd.n1963 gnd.n1961 10.6151
R10684 gnd.n2395 gnd.n2394 10.6151
R10685 gnd.n2394 gnd.n2391 10.6151
R10686 gnd.n2389 gnd.n2386 10.6151
R10687 gnd.n2386 gnd.n2385 10.6151
R10688 gnd.n2385 gnd.n2382 10.6151
R10689 gnd.n2382 gnd.n2381 10.6151
R10690 gnd.n2381 gnd.n2378 10.6151
R10691 gnd.n2378 gnd.n2377 10.6151
R10692 gnd.n2377 gnd.n2374 10.6151
R10693 gnd.n2374 gnd.n2373 10.6151
R10694 gnd.n2373 gnd.n2370 10.6151
R10695 gnd.n2370 gnd.n2369 10.6151
R10696 gnd.n2369 gnd.n2366 10.6151
R10697 gnd.n2366 gnd.n2365 10.6151
R10698 gnd.n2365 gnd.n2362 10.6151
R10699 gnd.n2362 gnd.n2361 10.6151
R10700 gnd.n2361 gnd.n2358 10.6151
R10701 gnd.n2358 gnd.n2357 10.6151
R10702 gnd.n2357 gnd.n2354 10.6151
R10703 gnd.n2354 gnd.n2353 10.6151
R10704 gnd.n2353 gnd.n2350 10.6151
R10705 gnd.n2350 gnd.n2349 10.6151
R10706 gnd.n2349 gnd.n2346 10.6151
R10707 gnd.n2346 gnd.n2345 10.6151
R10708 gnd.n2345 gnd.n2342 10.6151
R10709 gnd.n2342 gnd.n2341 10.6151
R10710 gnd.n2341 gnd.n2338 10.6151
R10711 gnd.n2338 gnd.n2337 10.6151
R10712 gnd.n2337 gnd.n2334 10.6151
R10713 gnd.n2334 gnd.n2333 10.6151
R10714 gnd.n3351 gnd.n2287 10.6151
R10715 gnd.n3346 gnd.n2287 10.6151
R10716 gnd.n3346 gnd.n3345 10.6151
R10717 gnd.n3345 gnd.n3344 10.6151
R10718 gnd.n3344 gnd.n3341 10.6151
R10719 gnd.n3341 gnd.n3340 10.6151
R10720 gnd.n3340 gnd.n3337 10.6151
R10721 gnd.n3337 gnd.n3336 10.6151
R10722 gnd.n3336 gnd.n3333 10.6151
R10723 gnd.n3333 gnd.n3332 10.6151
R10724 gnd.n3332 gnd.n3329 10.6151
R10725 gnd.n3329 gnd.n3328 10.6151
R10726 gnd.n3328 gnd.n3325 10.6151
R10727 gnd.n3325 gnd.n3324 10.6151
R10728 gnd.n3324 gnd.n3321 10.6151
R10729 gnd.n3321 gnd.n3320 10.6151
R10730 gnd.n3320 gnd.n3317 10.6151
R10731 gnd.n3317 gnd.n3316 10.6151
R10732 gnd.n3316 gnd.n3313 10.6151
R10733 gnd.n3313 gnd.n3312 10.6151
R10734 gnd.n3312 gnd.n3309 10.6151
R10735 gnd.n3309 gnd.n3308 10.6151
R10736 gnd.n3308 gnd.n3305 10.6151
R10737 gnd.n3305 gnd.n3304 10.6151
R10738 gnd.n3304 gnd.n3301 10.6151
R10739 gnd.n3301 gnd.n3300 10.6151
R10740 gnd.n3300 gnd.n3297 10.6151
R10741 gnd.n3297 gnd.n3296 10.6151
R10742 gnd.n3293 gnd.n3292 10.6151
R10743 gnd.n3292 gnd.n3289 10.6151
R10744 gnd.n3974 gnd.n3972 10.6151
R10745 gnd.n3972 gnd.n3969 10.6151
R10746 gnd.n3969 gnd.n3968 10.6151
R10747 gnd.n3968 gnd.n3965 10.6151
R10748 gnd.n3965 gnd.n3964 10.6151
R10749 gnd.n3964 gnd.n3961 10.6151
R10750 gnd.n3961 gnd.n3960 10.6151
R10751 gnd.n3960 gnd.n3957 10.6151
R10752 gnd.n3957 gnd.n3956 10.6151
R10753 gnd.n3956 gnd.n3953 10.6151
R10754 gnd.n3953 gnd.n3952 10.6151
R10755 gnd.n3952 gnd.n3949 10.6151
R10756 gnd.n3949 gnd.n3948 10.6151
R10757 gnd.n3948 gnd.n3945 10.6151
R10758 gnd.n3945 gnd.n3944 10.6151
R10759 gnd.n3944 gnd.n3941 10.6151
R10760 gnd.n3941 gnd.n3940 10.6151
R10761 gnd.n3940 gnd.n3937 10.6151
R10762 gnd.n3937 gnd.n3936 10.6151
R10763 gnd.n3936 gnd.n3933 10.6151
R10764 gnd.n3933 gnd.n3932 10.6151
R10765 gnd.n3932 gnd.n3929 10.6151
R10766 gnd.n3929 gnd.n3928 10.6151
R10767 gnd.n3928 gnd.n3925 10.6151
R10768 gnd.n3925 gnd.n3924 10.6151
R10769 gnd.n3924 gnd.n3921 10.6151
R10770 gnd.n3921 gnd.n3920 10.6151
R10771 gnd.n3920 gnd.n3917 10.6151
R10772 gnd.n3915 gnd.n3912 10.6151
R10773 gnd.n3912 gnd.n3911 10.6151
R10774 gnd.n3355 gnd.n3353 10.6151
R10775 gnd.n3355 gnd.n3354 10.6151
R10776 gnd.n3354 gnd.n2247 10.6151
R10777 gnd.n3442 gnd.n2247 10.6151
R10778 gnd.n3443 gnd.n3442 10.6151
R10779 gnd.n3447 gnd.n3443 10.6151
R10780 gnd.n3447 gnd.n3446 10.6151
R10781 gnd.n3446 gnd.n3445 10.6151
R10782 gnd.n3445 gnd.n2225 10.6151
R10783 gnd.n3473 gnd.n2225 10.6151
R10784 gnd.n3474 gnd.n3473 10.6151
R10785 gnd.n3478 gnd.n3474 10.6151
R10786 gnd.n3478 gnd.n3477 10.6151
R10787 gnd.n3477 gnd.n3476 10.6151
R10788 gnd.n3476 gnd.n2203 10.6151
R10789 gnd.n3504 gnd.n2203 10.6151
R10790 gnd.n3505 gnd.n3504 10.6151
R10791 gnd.n3506 gnd.n3505 10.6151
R10792 gnd.n3506 gnd.n2188 10.6151
R10793 gnd.n3522 gnd.n2188 10.6151
R10794 gnd.n3523 gnd.n3522 10.6151
R10795 gnd.n3524 gnd.n3523 10.6151
R10796 gnd.n3524 gnd.n2175 10.6151
R10797 gnd.n3538 gnd.n2175 10.6151
R10798 gnd.n3539 gnd.n3538 10.6151
R10799 gnd.n3541 gnd.n3539 10.6151
R10800 gnd.n3541 gnd.n3540 10.6151
R10801 gnd.n3540 gnd.n2151 10.6151
R10802 gnd.n3569 gnd.n2151 10.6151
R10803 gnd.n3570 gnd.n3569 10.6151
R10804 gnd.n3571 gnd.n3570 10.6151
R10805 gnd.n3571 gnd.n2137 10.6151
R10806 gnd.n3588 gnd.n2137 10.6151
R10807 gnd.n3589 gnd.n3588 10.6151
R10808 gnd.n3590 gnd.n3589 10.6151
R10809 gnd.n3590 gnd.n2122 10.6151
R10810 gnd.n3620 gnd.n2122 10.6151
R10811 gnd.n3621 gnd.n3620 10.6151
R10812 gnd.n3622 gnd.n3621 10.6151
R10813 gnd.n3622 gnd.n2107 10.6151
R10814 gnd.n3636 gnd.n2107 10.6151
R10815 gnd.n3637 gnd.n3636 10.6151
R10816 gnd.n3639 gnd.n3637 10.6151
R10817 gnd.n3639 gnd.n3638 10.6151
R10818 gnd.n3638 gnd.n2086 10.6151
R10819 gnd.n3670 gnd.n2086 10.6151
R10820 gnd.n3671 gnd.n3670 10.6151
R10821 gnd.n3672 gnd.n3671 10.6151
R10822 gnd.n3672 gnd.n2071 10.6151
R10823 gnd.n3697 gnd.n2071 10.6151
R10824 gnd.n3698 gnd.n3697 10.6151
R10825 gnd.n3702 gnd.n3698 10.6151
R10826 gnd.n3702 gnd.n3701 10.6151
R10827 gnd.n3701 gnd.n3700 10.6151
R10828 gnd.n3700 gnd.n2049 10.6151
R10829 gnd.n3737 gnd.n2049 10.6151
R10830 gnd.n3738 gnd.n3737 10.6151
R10831 gnd.n3742 gnd.n3738 10.6151
R10832 gnd.n3742 gnd.n3741 10.6151
R10833 gnd.n3741 gnd.n3740 10.6151
R10834 gnd.n3740 gnd.n2026 10.6151
R10835 gnd.n3776 gnd.n2026 10.6151
R10836 gnd.n3777 gnd.n3776 10.6151
R10837 gnd.n3781 gnd.n3777 10.6151
R10838 gnd.n3781 gnd.n3780 10.6151
R10839 gnd.n3780 gnd.n3779 10.6151
R10840 gnd.n3779 gnd.n2005 10.6151
R10841 gnd.n3816 gnd.n2005 10.6151
R10842 gnd.n3817 gnd.n3816 10.6151
R10843 gnd.n3821 gnd.n3817 10.6151
R10844 gnd.n3821 gnd.n3820 10.6151
R10845 gnd.n3820 gnd.n3819 10.6151
R10846 gnd.n3819 gnd.n1981 10.6151
R10847 gnd.n3864 gnd.n1981 10.6151
R10848 gnd.n3865 gnd.n3864 10.6151
R10849 gnd.n3866 gnd.n3865 10.6151
R10850 gnd.n3866 gnd.n1968 10.6151
R10851 gnd.n3886 gnd.n1968 10.6151
R10852 gnd.n3887 gnd.n3886 10.6151
R10853 gnd.n3977 gnd.n3887 10.6151
R10854 gnd.n3977 gnd.n3976 10.6151
R10855 gnd.n5338 gnd.t163 10.5161
R10856 gnd.n5948 gnd.t23 10.5161
R10857 gnd.n5955 gnd.t14 10.5161
R10858 gnd.t211 gnd.n1204 10.5161
R10859 gnd.n2886 gnd.t186 10.5161
R10860 gnd.n4576 gnd.t186 10.5161
R10861 gnd.n4569 gnd.t182 10.5161
R10862 gnd.n3501 gnd.t143 10.5161
R10863 gnd.n2035 gnd.t276 10.5161
R10864 gnd.n4314 gnd.t204 10.5161
R10865 gnd.t195 gnd.n1518 10.5161
R10866 gnd.n4288 gnd.t195 10.5161
R10867 gnd.n7093 gnd.t230 10.5161
R10868 gnd.n5910 gnd.n5894 10.4732
R10869 gnd.n5878 gnd.n5862 10.4732
R10870 gnd.n5846 gnd.n5830 10.4732
R10871 gnd.n5815 gnd.n5799 10.4732
R10872 gnd.n5783 gnd.n5767 10.4732
R10873 gnd.n5751 gnd.n5735 10.4732
R10874 gnd.n5719 gnd.n5703 10.4732
R10875 gnd.n5688 gnd.n5672 10.4732
R10876 gnd.n4715 gnd.n1069 10.1975
R10877 gnd.n3439 gnd.t28 10.1975
R10878 gnd.n2172 gnd.n2163 10.1975
R10879 gnd.n3567 gnd.n3566 10.1975
R10880 gnd.n3705 gnd.n3704 10.1975
R10881 gnd.n3713 gnd.n2061 10.1975
R10882 gnd.n1990 gnd.t57 10.1975
R10883 gnd.n3847 gnd.n1990 10.1975
R10884 gnd.n3850 gnd.n1964 10.1975
R10885 gnd.n7033 gnd.n94 10.1975
R10886 gnd.n5623 gnd.t20 9.87883
R10887 gnd.n2648 gnd.t184 9.87883
R10888 gnd.n2825 gnd.t197 9.87883
R10889 gnd.n2906 gnd.t174 9.87883
R10890 gnd.n4544 gnd.t188 9.87883
R10891 gnd.t282 gnd.n3617 9.87883
R10892 gnd.n2104 gnd.t278 9.87883
R10893 gnd.n4213 gnd.t240 9.87883
R10894 gnd.t180 gnd.n1502 9.87883
R10895 gnd.n7078 gnd.t192 9.87883
R10896 gnd.n7073 gnd.t237 9.87883
R10897 gnd.n5914 gnd.n5913 9.69747
R10898 gnd.n5882 gnd.n5881 9.69747
R10899 gnd.n5850 gnd.n5849 9.69747
R10900 gnd.n5819 gnd.n5818 9.69747
R10901 gnd.n5787 gnd.n5786 9.69747
R10902 gnd.n5755 gnd.n5754 9.69747
R10903 gnd.n5723 gnd.n5722 9.69747
R10904 gnd.n5692 gnd.n5691 9.69747
R10905 gnd.n7361 gnd.n50 9.6512
R10906 gnd.n3422 gnd.n2222 9.56018
R10907 gnd.n3508 gnd.n2201 9.56018
R10908 gnd.n3617 gnd.n2118 9.56018
R10909 gnd.n3641 gnd.n2104 9.56018
R10910 gnd.n3774 gnd.n2021 9.56018
R10911 gnd.n3814 gnd.n3813 9.56018
R10912 gnd.n3836 gnd.t78 9.56018
R10913 gnd.n4504 gnd.n1332 9.45599
R10914 gnd.n1648 gnd.n1647 9.45599
R10915 gnd.n5920 gnd.n5919 9.45567
R10916 gnd.n5888 gnd.n5887 9.45567
R10917 gnd.n5856 gnd.n5855 9.45567
R10918 gnd.n5825 gnd.n5824 9.45567
R10919 gnd.n5793 gnd.n5792 9.45567
R10920 gnd.n5761 gnd.n5760 9.45567
R10921 gnd.n5729 gnd.n5728 9.45567
R10922 gnd.n5698 gnd.n5697 9.45567
R10923 gnd.n4936 gnd.n4935 9.39724
R10924 gnd.n5919 gnd.n5918 9.3005
R10925 gnd.n5892 gnd.n5891 9.3005
R10926 gnd.n5913 gnd.n5912 9.3005
R10927 gnd.n5911 gnd.n5910 9.3005
R10928 gnd.n5896 gnd.n5895 9.3005
R10929 gnd.n5905 gnd.n5904 9.3005
R10930 gnd.n5903 gnd.n5902 9.3005
R10931 gnd.n5887 gnd.n5886 9.3005
R10932 gnd.n5860 gnd.n5859 9.3005
R10933 gnd.n5881 gnd.n5880 9.3005
R10934 gnd.n5879 gnd.n5878 9.3005
R10935 gnd.n5864 gnd.n5863 9.3005
R10936 gnd.n5873 gnd.n5872 9.3005
R10937 gnd.n5871 gnd.n5870 9.3005
R10938 gnd.n5855 gnd.n5854 9.3005
R10939 gnd.n5828 gnd.n5827 9.3005
R10940 gnd.n5849 gnd.n5848 9.3005
R10941 gnd.n5847 gnd.n5846 9.3005
R10942 gnd.n5832 gnd.n5831 9.3005
R10943 gnd.n5841 gnd.n5840 9.3005
R10944 gnd.n5839 gnd.n5838 9.3005
R10945 gnd.n5824 gnd.n5823 9.3005
R10946 gnd.n5797 gnd.n5796 9.3005
R10947 gnd.n5818 gnd.n5817 9.3005
R10948 gnd.n5816 gnd.n5815 9.3005
R10949 gnd.n5801 gnd.n5800 9.3005
R10950 gnd.n5810 gnd.n5809 9.3005
R10951 gnd.n5808 gnd.n5807 9.3005
R10952 gnd.n5792 gnd.n5791 9.3005
R10953 gnd.n5765 gnd.n5764 9.3005
R10954 gnd.n5786 gnd.n5785 9.3005
R10955 gnd.n5784 gnd.n5783 9.3005
R10956 gnd.n5769 gnd.n5768 9.3005
R10957 gnd.n5778 gnd.n5777 9.3005
R10958 gnd.n5776 gnd.n5775 9.3005
R10959 gnd.n5760 gnd.n5759 9.3005
R10960 gnd.n5733 gnd.n5732 9.3005
R10961 gnd.n5754 gnd.n5753 9.3005
R10962 gnd.n5752 gnd.n5751 9.3005
R10963 gnd.n5737 gnd.n5736 9.3005
R10964 gnd.n5746 gnd.n5745 9.3005
R10965 gnd.n5744 gnd.n5743 9.3005
R10966 gnd.n5728 gnd.n5727 9.3005
R10967 gnd.n5701 gnd.n5700 9.3005
R10968 gnd.n5722 gnd.n5721 9.3005
R10969 gnd.n5720 gnd.n5719 9.3005
R10970 gnd.n5705 gnd.n5704 9.3005
R10971 gnd.n5714 gnd.n5713 9.3005
R10972 gnd.n5712 gnd.n5711 9.3005
R10973 gnd.n5697 gnd.n5696 9.3005
R10974 gnd.n5670 gnd.n5669 9.3005
R10975 gnd.n5691 gnd.n5690 9.3005
R10976 gnd.n5689 gnd.n5688 9.3005
R10977 gnd.n5674 gnd.n5673 9.3005
R10978 gnd.n5683 gnd.n5682 9.3005
R10979 gnd.n5681 gnd.n5680 9.3005
R10980 gnd.n6049 gnd.n4747 9.3005
R10981 gnd.n6048 gnd.n4749 9.3005
R10982 gnd.n4753 gnd.n4750 9.3005
R10983 gnd.n6043 gnd.n4754 9.3005
R10984 gnd.n6042 gnd.n4755 9.3005
R10985 gnd.n6041 gnd.n4756 9.3005
R10986 gnd.n4760 gnd.n4757 9.3005
R10987 gnd.n6036 gnd.n4761 9.3005
R10988 gnd.n6035 gnd.n4762 9.3005
R10989 gnd.n6034 gnd.n4763 9.3005
R10990 gnd.n4767 gnd.n4764 9.3005
R10991 gnd.n6029 gnd.n4768 9.3005
R10992 gnd.n6028 gnd.n4769 9.3005
R10993 gnd.n6027 gnd.n4770 9.3005
R10994 gnd.n4775 gnd.n4773 9.3005
R10995 gnd.n6022 gnd.n6021 9.3005
R10996 gnd.n6051 gnd.n6050 9.3005
R10997 gnd.n5357 gnd.n5356 9.3005
R10998 gnd.n5061 gnd.n5060 9.3005
R10999 gnd.n5384 gnd.n5383 9.3005
R11000 gnd.n5385 gnd.n5059 9.3005
R11001 gnd.n5389 gnd.n5386 9.3005
R11002 gnd.n5388 gnd.n5387 9.3005
R11003 gnd.n5033 gnd.n5032 9.3005
R11004 gnd.n5414 gnd.n5413 9.3005
R11005 gnd.n5415 gnd.n5031 9.3005
R11006 gnd.n5417 gnd.n5416 9.3005
R11007 gnd.n5011 gnd.n5010 9.3005
R11008 gnd.n5445 gnd.n5444 9.3005
R11009 gnd.n5446 gnd.n5009 9.3005
R11010 gnd.n5454 gnd.n5447 9.3005
R11011 gnd.n5453 gnd.n5448 9.3005
R11012 gnd.n5452 gnd.n5450 9.3005
R11013 gnd.n5449 gnd.n4958 9.3005
R11014 gnd.n5502 gnd.n4959 9.3005
R11015 gnd.n5501 gnd.n4960 9.3005
R11016 gnd.n5500 gnd.n4961 9.3005
R11017 gnd.n4980 gnd.n4962 9.3005
R11018 gnd.n4982 gnd.n4981 9.3005
R11019 gnd.n4892 gnd.n4891 9.3005
R11020 gnd.n5540 gnd.n5539 9.3005
R11021 gnd.n5541 gnd.n4890 9.3005
R11022 gnd.n5545 gnd.n5542 9.3005
R11023 gnd.n5544 gnd.n5543 9.3005
R11024 gnd.n4865 gnd.n4864 9.3005
R11025 gnd.n5580 gnd.n5579 9.3005
R11026 gnd.n5581 gnd.n4863 9.3005
R11027 gnd.n5585 gnd.n5582 9.3005
R11028 gnd.n5584 gnd.n5583 9.3005
R11029 gnd.n4839 gnd.n4838 9.3005
R11030 gnd.n5636 gnd.n5635 9.3005
R11031 gnd.n5637 gnd.n4837 9.3005
R11032 gnd.n5640 gnd.n5639 9.3005
R11033 gnd.n5638 gnd.n946 9.3005
R11034 gnd.n6095 gnd.n947 9.3005
R11035 gnd.n6094 gnd.n948 9.3005
R11036 gnd.n6093 gnd.n949 9.3005
R11037 gnd.n970 gnd.n950 9.3005
R11038 gnd.n971 gnd.n969 9.3005
R11039 gnd.n6081 gnd.n972 9.3005
R11040 gnd.n6080 gnd.n973 9.3005
R11041 gnd.n6079 gnd.n974 9.3005
R11042 gnd.n996 gnd.n975 9.3005
R11043 gnd.n997 gnd.n995 9.3005
R11044 gnd.n6067 gnd.n998 9.3005
R11045 gnd.n6066 gnd.n999 9.3005
R11046 gnd.n6065 gnd.n1000 9.3005
R11047 gnd.n4745 gnd.n1001 9.3005
R11048 gnd.n4746 gnd.n4744 9.3005
R11049 gnd.n6053 gnd.n6052 9.3005
R11050 gnd.n5358 gnd.n5355 9.3005
R11051 gnd.n5140 gnd.n5099 9.3005
R11052 gnd.n5135 gnd.n5134 9.3005
R11053 gnd.n5133 gnd.n5100 9.3005
R11054 gnd.n5132 gnd.n5131 9.3005
R11055 gnd.n5128 gnd.n5101 9.3005
R11056 gnd.n5125 gnd.n5124 9.3005
R11057 gnd.n5123 gnd.n5102 9.3005
R11058 gnd.n5122 gnd.n5121 9.3005
R11059 gnd.n5118 gnd.n5103 9.3005
R11060 gnd.n5115 gnd.n5114 9.3005
R11061 gnd.n5113 gnd.n5104 9.3005
R11062 gnd.n5112 gnd.n5111 9.3005
R11063 gnd.n5108 gnd.n5106 9.3005
R11064 gnd.n5105 gnd.n5085 9.3005
R11065 gnd.n5352 gnd.n5084 9.3005
R11066 gnd.n5354 gnd.n5353 9.3005
R11067 gnd.n5142 gnd.n5141 9.3005
R11068 gnd.n5365 gnd.n5071 9.3005
R11069 gnd.n5372 gnd.n5072 9.3005
R11070 gnd.n5374 gnd.n5373 9.3005
R11071 gnd.n5375 gnd.n5052 9.3005
R11072 gnd.n5394 gnd.n5393 9.3005
R11073 gnd.n5396 gnd.n5044 9.3005
R11074 gnd.n5403 gnd.n5046 9.3005
R11075 gnd.n5404 gnd.n5041 9.3005
R11076 gnd.n5406 gnd.n5405 9.3005
R11077 gnd.n5042 gnd.n5027 9.3005
R11078 gnd.n5422 gnd.n5025 9.3005
R11079 gnd.n5426 gnd.n5425 9.3005
R11080 gnd.n5424 gnd.n5001 9.3005
R11081 gnd.n5461 gnd.n5000 9.3005
R11082 gnd.n5464 gnd.n5463 9.3005
R11083 gnd.n4997 gnd.n4996 9.3005
R11084 gnd.n5470 gnd.n4998 9.3005
R11085 gnd.n5472 gnd.n5471 9.3005
R11086 gnd.n5474 gnd.n4995 9.3005
R11087 gnd.n5477 gnd.n5476 9.3005
R11088 gnd.n5480 gnd.n5478 9.3005
R11089 gnd.n5482 gnd.n5481 9.3005
R11090 gnd.n5488 gnd.n5483 9.3005
R11091 gnd.n5487 gnd.n5486 9.3005
R11092 gnd.n4883 gnd.n4882 9.3005
R11093 gnd.n5554 gnd.n5553 9.3005
R11094 gnd.n5555 gnd.n4876 9.3005
R11095 gnd.n5563 gnd.n4875 9.3005
R11096 gnd.n5566 gnd.n5565 9.3005
R11097 gnd.n5568 gnd.n5567 9.3005
R11098 gnd.n5571 gnd.n4858 9.3005
R11099 gnd.n5569 gnd.n4856 9.3005
R11100 gnd.n5591 gnd.n4854 9.3005
R11101 gnd.n5595 gnd.n5594 9.3005
R11102 gnd.n5593 gnd.n5592 9.3005
R11103 gnd.n4832 gnd.n4831 9.3005
R11104 gnd.n5645 gnd.n4833 9.3005
R11105 gnd.n5647 gnd.n5646 9.3005
R11106 gnd.n5649 gnd.n4830 9.3005
R11107 gnd.n5652 gnd.n5651 9.3005
R11108 gnd.n5654 gnd.n5653 9.3005
R11109 gnd.n5658 gnd.n5655 9.3005
R11110 gnd.n5660 gnd.n5659 9.3005
R11111 gnd.n5945 gnd.n5662 9.3005
R11112 gnd.n5944 gnd.n5664 9.3005
R11113 gnd.n5943 gnd.n5665 9.3005
R11114 gnd.n5940 gnd.n5666 9.3005
R11115 gnd.n5939 gnd.n5667 9.3005
R11116 gnd.n5938 gnd.n5925 9.3005
R11117 gnd.n5935 gnd.n5927 9.3005
R11118 gnd.n5934 gnd.n5928 9.3005
R11119 gnd.n5931 gnd.n5929 9.3005
R11120 gnd.n5930 gnd.n4776 9.3005
R11121 gnd.n5363 gnd.n5362 9.3005
R11122 gnd.n6017 gnd.n4777 9.3005
R11123 gnd.n6016 gnd.n4779 9.3005
R11124 gnd.n4783 gnd.n4780 9.3005
R11125 gnd.n6011 gnd.n4784 9.3005
R11126 gnd.n6010 gnd.n4785 9.3005
R11127 gnd.n6009 gnd.n4786 9.3005
R11128 gnd.n4790 gnd.n4787 9.3005
R11129 gnd.n6004 gnd.n4791 9.3005
R11130 gnd.n6003 gnd.n4792 9.3005
R11131 gnd.n6002 gnd.n4793 9.3005
R11132 gnd.n4797 gnd.n4794 9.3005
R11133 gnd.n5997 gnd.n4798 9.3005
R11134 gnd.n5996 gnd.n4799 9.3005
R11135 gnd.n5995 gnd.n4800 9.3005
R11136 gnd.n4804 gnd.n4801 9.3005
R11137 gnd.n5990 gnd.n4805 9.3005
R11138 gnd.n5989 gnd.n4806 9.3005
R11139 gnd.n5988 gnd.n4807 9.3005
R11140 gnd.n4811 gnd.n4808 9.3005
R11141 gnd.n5983 gnd.n4812 9.3005
R11142 gnd.n5982 gnd.n4813 9.3005
R11143 gnd.n5981 gnd.n4814 9.3005
R11144 gnd.n4821 gnd.n4819 9.3005
R11145 gnd.n5976 gnd.n4822 9.3005
R11146 gnd.n5975 gnd.n4823 9.3005
R11147 gnd.n5974 gnd.n5971 9.3005
R11148 gnd.n6019 gnd.n6018 9.3005
R11149 gnd.n5532 gnd.n5516 9.3005
R11150 gnd.n5531 gnd.n5517 9.3005
R11151 gnd.n5530 gnd.n5518 9.3005
R11152 gnd.n5528 gnd.n5519 9.3005
R11153 gnd.n5527 gnd.n5520 9.3005
R11154 gnd.n5525 gnd.n5521 9.3005
R11155 gnd.n5524 gnd.n5522 9.3005
R11156 gnd.n4846 gnd.n4845 9.3005
R11157 gnd.n5603 gnd.n5602 9.3005
R11158 gnd.n5604 gnd.n4844 9.3005
R11159 gnd.n5630 gnd.n5605 9.3005
R11160 gnd.n5629 gnd.n5606 9.3005
R11161 gnd.n5628 gnd.n5607 9.3005
R11162 gnd.n5626 gnd.n5608 9.3005
R11163 gnd.n5625 gnd.n5609 9.3005
R11164 gnd.n5619 gnd.n5610 9.3005
R11165 gnd.n5618 gnd.n5611 9.3005
R11166 gnd.n5617 gnd.n5612 9.3005
R11167 gnd.n5614 gnd.n5613 9.3005
R11168 gnd.n4829 gnd.n4828 9.3005
R11169 gnd.n5952 gnd.n5951 9.3005
R11170 gnd.n5953 gnd.n4827 9.3005
R11171 gnd.n5957 gnd.n5954 9.3005
R11172 gnd.n5958 gnd.n4826 9.3005
R11173 gnd.n5962 gnd.n5961 9.3005
R11174 gnd.n5963 gnd.n4825 9.3005
R11175 gnd.n5965 gnd.n5964 9.3005
R11176 gnd.n5968 gnd.n4824 9.3005
R11177 gnd.n5970 gnd.n5969 9.3005
R11178 gnd.n5273 gnd.n5272 9.3005
R11179 gnd.n5163 gnd.n5162 9.3005
R11180 gnd.n5287 gnd.n5286 9.3005
R11181 gnd.n5288 gnd.n5161 9.3005
R11182 gnd.n5290 gnd.n5289 9.3005
R11183 gnd.n5151 gnd.n5150 9.3005
R11184 gnd.n5303 gnd.n5302 9.3005
R11185 gnd.n5304 gnd.n5149 9.3005
R11186 gnd.n5336 gnd.n5305 9.3005
R11187 gnd.n5335 gnd.n5306 9.3005
R11188 gnd.n5334 gnd.n5307 9.3005
R11189 gnd.n5333 gnd.n5308 9.3005
R11190 gnd.n5330 gnd.n5309 9.3005
R11191 gnd.n5329 gnd.n5310 9.3005
R11192 gnd.n5328 gnd.n5311 9.3005
R11193 gnd.n5326 gnd.n5312 9.3005
R11194 gnd.n5325 gnd.n5313 9.3005
R11195 gnd.n5322 gnd.n5314 9.3005
R11196 gnd.n5321 gnd.n5315 9.3005
R11197 gnd.n5320 gnd.n5316 9.3005
R11198 gnd.n5318 gnd.n5317 9.3005
R11199 gnd.n5017 gnd.n5016 9.3005
R11200 gnd.n5434 gnd.n5433 9.3005
R11201 gnd.n5435 gnd.n5015 9.3005
R11202 gnd.n5439 gnd.n5436 9.3005
R11203 gnd.n5438 gnd.n5437 9.3005
R11204 gnd.n4939 gnd.n4938 9.3005
R11205 gnd.n5514 gnd.n5513 9.3005
R11206 gnd.n5271 gnd.n5172 9.3005
R11207 gnd.n5174 gnd.n5173 9.3005
R11208 gnd.n5218 gnd.n5216 9.3005
R11209 gnd.n5219 gnd.n5215 9.3005
R11210 gnd.n5222 gnd.n5211 9.3005
R11211 gnd.n5223 gnd.n5210 9.3005
R11212 gnd.n5226 gnd.n5209 9.3005
R11213 gnd.n5227 gnd.n5208 9.3005
R11214 gnd.n5230 gnd.n5207 9.3005
R11215 gnd.n5231 gnd.n5206 9.3005
R11216 gnd.n5234 gnd.n5205 9.3005
R11217 gnd.n5235 gnd.n5204 9.3005
R11218 gnd.n5238 gnd.n5203 9.3005
R11219 gnd.n5239 gnd.n5202 9.3005
R11220 gnd.n5242 gnd.n5201 9.3005
R11221 gnd.n5243 gnd.n5200 9.3005
R11222 gnd.n5246 gnd.n5199 9.3005
R11223 gnd.n5247 gnd.n5198 9.3005
R11224 gnd.n5250 gnd.n5197 9.3005
R11225 gnd.n5251 gnd.n5196 9.3005
R11226 gnd.n5254 gnd.n5195 9.3005
R11227 gnd.n5255 gnd.n5194 9.3005
R11228 gnd.n5258 gnd.n5193 9.3005
R11229 gnd.n5260 gnd.n5192 9.3005
R11230 gnd.n5261 gnd.n5191 9.3005
R11231 gnd.n5262 gnd.n5190 9.3005
R11232 gnd.n5263 gnd.n5189 9.3005
R11233 gnd.n5270 gnd.n5269 9.3005
R11234 gnd.n5279 gnd.n5278 9.3005
R11235 gnd.n5280 gnd.n5166 9.3005
R11236 gnd.n5282 gnd.n5281 9.3005
R11237 gnd.n5157 gnd.n5156 9.3005
R11238 gnd.n5295 gnd.n5294 9.3005
R11239 gnd.n5296 gnd.n5155 9.3005
R11240 gnd.n5298 gnd.n5297 9.3005
R11241 gnd.n5144 gnd.n5143 9.3005
R11242 gnd.n5341 gnd.n5340 9.3005
R11243 gnd.n5342 gnd.n5098 9.3005
R11244 gnd.n5346 gnd.n5344 9.3005
R11245 gnd.n5345 gnd.n5077 9.3005
R11246 gnd.n5364 gnd.n5076 9.3005
R11247 gnd.n5367 gnd.n5366 9.3005
R11248 gnd.n5070 gnd.n5069 9.3005
R11249 gnd.n5378 gnd.n5376 9.3005
R11250 gnd.n5377 gnd.n5051 9.3005
R11251 gnd.n5395 gnd.n5050 9.3005
R11252 gnd.n5398 gnd.n5397 9.3005
R11253 gnd.n5045 gnd.n5040 9.3005
R11254 gnd.n5408 gnd.n5407 9.3005
R11255 gnd.n5043 gnd.n5023 9.3005
R11256 gnd.n5429 gnd.n5024 9.3005
R11257 gnd.n5428 gnd.n5427 9.3005
R11258 gnd.n5026 gnd.n5002 9.3005
R11259 gnd.n5460 gnd.n5459 9.3005
R11260 gnd.n5462 gnd.n4947 9.3005
R11261 gnd.n5509 gnd.n4948 9.3005
R11262 gnd.n5508 gnd.n4949 9.3005
R11263 gnd.n5507 gnd.n4950 9.3005
R11264 gnd.n5473 gnd.n4951 9.3005
R11265 gnd.n5475 gnd.n4969 9.3005
R11266 gnd.n5495 gnd.n4970 9.3005
R11267 gnd.n5494 gnd.n4971 9.3005
R11268 gnd.n5493 gnd.n4972 9.3005
R11269 gnd.n5484 gnd.n4973 9.3005
R11270 gnd.n5485 gnd.n4884 9.3005
R11271 gnd.n5551 gnd.n5550 9.3005
R11272 gnd.n5552 gnd.n4877 9.3005
R11273 gnd.n5562 gnd.n5561 9.3005
R11274 gnd.n5564 gnd.n4873 9.3005
R11275 gnd.n5574 gnd.n4874 9.3005
R11276 gnd.n5573 gnd.n5572 9.3005
R11277 gnd.n5570 gnd.n4852 9.3005
R11278 gnd.n5598 gnd.n4853 9.3005
R11279 gnd.n5597 gnd.n5596 9.3005
R11280 gnd.n4855 gnd.n935 9.3005
R11281 gnd.n6102 gnd.n936 9.3005
R11282 gnd.n6101 gnd.n937 9.3005
R11283 gnd.n6100 gnd.n938 9.3005
R11284 gnd.n5648 gnd.n939 9.3005
R11285 gnd.n5650 gnd.n958 9.3005
R11286 gnd.n6088 gnd.n959 9.3005
R11287 gnd.n6087 gnd.n960 9.3005
R11288 gnd.n6086 gnd.n961 9.3005
R11289 gnd.n5661 gnd.n962 9.3005
R11290 gnd.n5663 gnd.n983 9.3005
R11291 gnd.n6074 gnd.n984 9.3005
R11292 gnd.n6073 gnd.n985 9.3005
R11293 gnd.n6072 gnd.n986 9.3005
R11294 gnd.n5924 gnd.n987 9.3005
R11295 gnd.n5926 gnd.n1009 9.3005
R11296 gnd.n6060 gnd.n1010 9.3005
R11297 gnd.n6059 gnd.n1011 9.3005
R11298 gnd.n6058 gnd.n1012 9.3005
R11299 gnd.n5168 gnd.n5167 9.3005
R11300 gnd.n6277 gnd.n6276 9.3005
R11301 gnd.n6278 gnd.n760 9.3005
R11302 gnd.n6280 gnd.n6279 9.3005
R11303 gnd.n756 gnd.n755 9.3005
R11304 gnd.n6287 gnd.n6286 9.3005
R11305 gnd.n6288 gnd.n754 9.3005
R11306 gnd.n6290 gnd.n6289 9.3005
R11307 gnd.n750 gnd.n749 9.3005
R11308 gnd.n6297 gnd.n6296 9.3005
R11309 gnd.n6298 gnd.n748 9.3005
R11310 gnd.n6300 gnd.n6299 9.3005
R11311 gnd.n744 gnd.n743 9.3005
R11312 gnd.n6307 gnd.n6306 9.3005
R11313 gnd.n6308 gnd.n742 9.3005
R11314 gnd.n6310 gnd.n6309 9.3005
R11315 gnd.n738 gnd.n737 9.3005
R11316 gnd.n6317 gnd.n6316 9.3005
R11317 gnd.n6318 gnd.n736 9.3005
R11318 gnd.n6320 gnd.n6319 9.3005
R11319 gnd.n732 gnd.n731 9.3005
R11320 gnd.n6327 gnd.n6326 9.3005
R11321 gnd.n6328 gnd.n730 9.3005
R11322 gnd.n6330 gnd.n6329 9.3005
R11323 gnd.n726 gnd.n725 9.3005
R11324 gnd.n6337 gnd.n6336 9.3005
R11325 gnd.n6338 gnd.n724 9.3005
R11326 gnd.n6340 gnd.n6339 9.3005
R11327 gnd.n720 gnd.n719 9.3005
R11328 gnd.n6347 gnd.n6346 9.3005
R11329 gnd.n6348 gnd.n718 9.3005
R11330 gnd.n6350 gnd.n6349 9.3005
R11331 gnd.n714 gnd.n713 9.3005
R11332 gnd.n6357 gnd.n6356 9.3005
R11333 gnd.n6358 gnd.n712 9.3005
R11334 gnd.n6360 gnd.n6359 9.3005
R11335 gnd.n708 gnd.n707 9.3005
R11336 gnd.n6367 gnd.n6366 9.3005
R11337 gnd.n6368 gnd.n706 9.3005
R11338 gnd.n6370 gnd.n6369 9.3005
R11339 gnd.n702 gnd.n701 9.3005
R11340 gnd.n6377 gnd.n6376 9.3005
R11341 gnd.n6378 gnd.n700 9.3005
R11342 gnd.n6380 gnd.n6379 9.3005
R11343 gnd.n696 gnd.n695 9.3005
R11344 gnd.n6387 gnd.n6386 9.3005
R11345 gnd.n6388 gnd.n694 9.3005
R11346 gnd.n6390 gnd.n6389 9.3005
R11347 gnd.n690 gnd.n689 9.3005
R11348 gnd.n6397 gnd.n6396 9.3005
R11349 gnd.n6398 gnd.n688 9.3005
R11350 gnd.n6400 gnd.n6399 9.3005
R11351 gnd.n684 gnd.n683 9.3005
R11352 gnd.n6407 gnd.n6406 9.3005
R11353 gnd.n6408 gnd.n682 9.3005
R11354 gnd.n6410 gnd.n6409 9.3005
R11355 gnd.n678 gnd.n677 9.3005
R11356 gnd.n6417 gnd.n6416 9.3005
R11357 gnd.n6418 gnd.n676 9.3005
R11358 gnd.n6420 gnd.n6419 9.3005
R11359 gnd.n672 gnd.n671 9.3005
R11360 gnd.n6427 gnd.n6426 9.3005
R11361 gnd.n6428 gnd.n670 9.3005
R11362 gnd.n6430 gnd.n6429 9.3005
R11363 gnd.n666 gnd.n665 9.3005
R11364 gnd.n6437 gnd.n6436 9.3005
R11365 gnd.n6438 gnd.n664 9.3005
R11366 gnd.n6440 gnd.n6439 9.3005
R11367 gnd.n660 gnd.n659 9.3005
R11368 gnd.n6447 gnd.n6446 9.3005
R11369 gnd.n6448 gnd.n658 9.3005
R11370 gnd.n6450 gnd.n6449 9.3005
R11371 gnd.n654 gnd.n653 9.3005
R11372 gnd.n6457 gnd.n6456 9.3005
R11373 gnd.n6458 gnd.n652 9.3005
R11374 gnd.n6460 gnd.n6459 9.3005
R11375 gnd.n648 gnd.n647 9.3005
R11376 gnd.n6467 gnd.n6466 9.3005
R11377 gnd.n6468 gnd.n646 9.3005
R11378 gnd.n6470 gnd.n6469 9.3005
R11379 gnd.n642 gnd.n641 9.3005
R11380 gnd.n6477 gnd.n6476 9.3005
R11381 gnd.n6478 gnd.n640 9.3005
R11382 gnd.n6480 gnd.n6479 9.3005
R11383 gnd.n636 gnd.n635 9.3005
R11384 gnd.n6487 gnd.n6486 9.3005
R11385 gnd.n6488 gnd.n634 9.3005
R11386 gnd.n6490 gnd.n6489 9.3005
R11387 gnd.n630 gnd.n629 9.3005
R11388 gnd.n6497 gnd.n6496 9.3005
R11389 gnd.n6498 gnd.n628 9.3005
R11390 gnd.n6500 gnd.n6499 9.3005
R11391 gnd.n624 gnd.n623 9.3005
R11392 gnd.n6507 gnd.n6506 9.3005
R11393 gnd.n6508 gnd.n622 9.3005
R11394 gnd.n6510 gnd.n6509 9.3005
R11395 gnd.n618 gnd.n617 9.3005
R11396 gnd.n6517 gnd.n6516 9.3005
R11397 gnd.n6518 gnd.n616 9.3005
R11398 gnd.n6520 gnd.n6519 9.3005
R11399 gnd.n612 gnd.n611 9.3005
R11400 gnd.n6527 gnd.n6526 9.3005
R11401 gnd.n6528 gnd.n610 9.3005
R11402 gnd.n6530 gnd.n6529 9.3005
R11403 gnd.n606 gnd.n605 9.3005
R11404 gnd.n6537 gnd.n6536 9.3005
R11405 gnd.n6538 gnd.n604 9.3005
R11406 gnd.n6540 gnd.n6539 9.3005
R11407 gnd.n600 gnd.n599 9.3005
R11408 gnd.n6547 gnd.n6546 9.3005
R11409 gnd.n6548 gnd.n598 9.3005
R11410 gnd.n6550 gnd.n6549 9.3005
R11411 gnd.n594 gnd.n593 9.3005
R11412 gnd.n6557 gnd.n6556 9.3005
R11413 gnd.n6558 gnd.n592 9.3005
R11414 gnd.n6560 gnd.n6559 9.3005
R11415 gnd.n588 gnd.n587 9.3005
R11416 gnd.n6567 gnd.n6566 9.3005
R11417 gnd.n6568 gnd.n586 9.3005
R11418 gnd.n6570 gnd.n6569 9.3005
R11419 gnd.n582 gnd.n581 9.3005
R11420 gnd.n6577 gnd.n6576 9.3005
R11421 gnd.n6578 gnd.n580 9.3005
R11422 gnd.n6580 gnd.n6579 9.3005
R11423 gnd.n576 gnd.n575 9.3005
R11424 gnd.n6587 gnd.n6586 9.3005
R11425 gnd.n6588 gnd.n574 9.3005
R11426 gnd.n6590 gnd.n6589 9.3005
R11427 gnd.n570 gnd.n569 9.3005
R11428 gnd.n6597 gnd.n6596 9.3005
R11429 gnd.n6598 gnd.n568 9.3005
R11430 gnd.n6600 gnd.n6599 9.3005
R11431 gnd.n564 gnd.n563 9.3005
R11432 gnd.n6607 gnd.n6606 9.3005
R11433 gnd.n6608 gnd.n562 9.3005
R11434 gnd.n6610 gnd.n6609 9.3005
R11435 gnd.n558 gnd.n557 9.3005
R11436 gnd.n6617 gnd.n6616 9.3005
R11437 gnd.n6618 gnd.n556 9.3005
R11438 gnd.n6620 gnd.n6619 9.3005
R11439 gnd.n552 gnd.n551 9.3005
R11440 gnd.n6627 gnd.n6626 9.3005
R11441 gnd.n6628 gnd.n550 9.3005
R11442 gnd.n6630 gnd.n6629 9.3005
R11443 gnd.n546 gnd.n545 9.3005
R11444 gnd.n6637 gnd.n6636 9.3005
R11445 gnd.n6638 gnd.n544 9.3005
R11446 gnd.n6640 gnd.n6639 9.3005
R11447 gnd.n540 gnd.n539 9.3005
R11448 gnd.n6647 gnd.n6646 9.3005
R11449 gnd.n6648 gnd.n538 9.3005
R11450 gnd.n6650 gnd.n6649 9.3005
R11451 gnd.n534 gnd.n533 9.3005
R11452 gnd.n6657 gnd.n6656 9.3005
R11453 gnd.n6658 gnd.n532 9.3005
R11454 gnd.n6660 gnd.n6659 9.3005
R11455 gnd.n528 gnd.n527 9.3005
R11456 gnd.n6667 gnd.n6666 9.3005
R11457 gnd.n6668 gnd.n526 9.3005
R11458 gnd.n6670 gnd.n6669 9.3005
R11459 gnd.n522 gnd.n521 9.3005
R11460 gnd.n6677 gnd.n6676 9.3005
R11461 gnd.n6678 gnd.n520 9.3005
R11462 gnd.n6680 gnd.n6679 9.3005
R11463 gnd.n516 gnd.n515 9.3005
R11464 gnd.n6687 gnd.n6686 9.3005
R11465 gnd.n6688 gnd.n514 9.3005
R11466 gnd.n6690 gnd.n6689 9.3005
R11467 gnd.n510 gnd.n509 9.3005
R11468 gnd.n6697 gnd.n6696 9.3005
R11469 gnd.n6698 gnd.n508 9.3005
R11470 gnd.n6700 gnd.n6699 9.3005
R11471 gnd.n504 gnd.n503 9.3005
R11472 gnd.n6707 gnd.n6706 9.3005
R11473 gnd.n6708 gnd.n502 9.3005
R11474 gnd.n6710 gnd.n6709 9.3005
R11475 gnd.n498 gnd.n497 9.3005
R11476 gnd.n6717 gnd.n6716 9.3005
R11477 gnd.n6718 gnd.n496 9.3005
R11478 gnd.n6720 gnd.n6719 9.3005
R11479 gnd.n492 gnd.n491 9.3005
R11480 gnd.n6727 gnd.n6726 9.3005
R11481 gnd.n6728 gnd.n490 9.3005
R11482 gnd.n6730 gnd.n6729 9.3005
R11483 gnd.n486 gnd.n485 9.3005
R11484 gnd.n6737 gnd.n6736 9.3005
R11485 gnd.n6738 gnd.n484 9.3005
R11486 gnd.n6740 gnd.n6739 9.3005
R11487 gnd.n480 gnd.n479 9.3005
R11488 gnd.n6747 gnd.n6746 9.3005
R11489 gnd.n6748 gnd.n478 9.3005
R11490 gnd.n6750 gnd.n6749 9.3005
R11491 gnd.n474 gnd.n473 9.3005
R11492 gnd.n6757 gnd.n6756 9.3005
R11493 gnd.n6758 gnd.n472 9.3005
R11494 gnd.n6760 gnd.n6759 9.3005
R11495 gnd.n468 gnd.n467 9.3005
R11496 gnd.n6767 gnd.n6766 9.3005
R11497 gnd.n6768 gnd.n466 9.3005
R11498 gnd.n6770 gnd.n6769 9.3005
R11499 gnd.n462 gnd.n461 9.3005
R11500 gnd.n6777 gnd.n6776 9.3005
R11501 gnd.n6778 gnd.n460 9.3005
R11502 gnd.n6780 gnd.n6779 9.3005
R11503 gnd.n456 gnd.n455 9.3005
R11504 gnd.n6787 gnd.n6786 9.3005
R11505 gnd.n6788 gnd.n454 9.3005
R11506 gnd.n6791 gnd.n6789 9.3005
R11507 gnd.n6790 gnd.n450 9.3005
R11508 gnd.n6799 gnd.n449 9.3005
R11509 gnd.n6801 gnd.n6800 9.3005
R11510 gnd.n445 gnd.n444 9.3005
R11511 gnd.n6808 gnd.n6807 9.3005
R11512 gnd.n6809 gnd.n443 9.3005
R11513 gnd.n6811 gnd.n6810 9.3005
R11514 gnd.n439 gnd.n438 9.3005
R11515 gnd.n6818 gnd.n6817 9.3005
R11516 gnd.n6819 gnd.n437 9.3005
R11517 gnd.n6821 gnd.n6820 9.3005
R11518 gnd.n433 gnd.n432 9.3005
R11519 gnd.n6828 gnd.n6827 9.3005
R11520 gnd.n6829 gnd.n431 9.3005
R11521 gnd.n6831 gnd.n6830 9.3005
R11522 gnd.n427 gnd.n426 9.3005
R11523 gnd.n6838 gnd.n6837 9.3005
R11524 gnd.n6839 gnd.n425 9.3005
R11525 gnd.n6841 gnd.n6840 9.3005
R11526 gnd.n421 gnd.n420 9.3005
R11527 gnd.n6848 gnd.n6847 9.3005
R11528 gnd.n6849 gnd.n419 9.3005
R11529 gnd.n6851 gnd.n6850 9.3005
R11530 gnd.n415 gnd.n414 9.3005
R11531 gnd.n6858 gnd.n6857 9.3005
R11532 gnd.n6859 gnd.n413 9.3005
R11533 gnd.n6861 gnd.n6860 9.3005
R11534 gnd.n409 gnd.n408 9.3005
R11535 gnd.n6868 gnd.n6867 9.3005
R11536 gnd.n6869 gnd.n407 9.3005
R11537 gnd.n6871 gnd.n6870 9.3005
R11538 gnd.n403 gnd.n402 9.3005
R11539 gnd.n6878 gnd.n6877 9.3005
R11540 gnd.n6879 gnd.n401 9.3005
R11541 gnd.n6881 gnd.n6880 9.3005
R11542 gnd.n397 gnd.n396 9.3005
R11543 gnd.n6888 gnd.n6887 9.3005
R11544 gnd.n6889 gnd.n395 9.3005
R11545 gnd.n6891 gnd.n6890 9.3005
R11546 gnd.n391 gnd.n390 9.3005
R11547 gnd.n6898 gnd.n6897 9.3005
R11548 gnd.n6899 gnd.n389 9.3005
R11549 gnd.n6901 gnd.n6900 9.3005
R11550 gnd.n385 gnd.n384 9.3005
R11551 gnd.n6908 gnd.n6907 9.3005
R11552 gnd.n6909 gnd.n383 9.3005
R11553 gnd.n6911 gnd.n6910 9.3005
R11554 gnd.n379 gnd.n378 9.3005
R11555 gnd.n6918 gnd.n6917 9.3005
R11556 gnd.n6919 gnd.n377 9.3005
R11557 gnd.n6921 gnd.n6920 9.3005
R11558 gnd.n373 gnd.n372 9.3005
R11559 gnd.n6928 gnd.n6927 9.3005
R11560 gnd.n6929 gnd.n371 9.3005
R11561 gnd.n6931 gnd.n6930 9.3005
R11562 gnd.n367 gnd.n366 9.3005
R11563 gnd.n6938 gnd.n6937 9.3005
R11564 gnd.n6939 gnd.n365 9.3005
R11565 gnd.n6941 gnd.n6940 9.3005
R11566 gnd.n361 gnd.n360 9.3005
R11567 gnd.n6948 gnd.n6947 9.3005
R11568 gnd.n6949 gnd.n359 9.3005
R11569 gnd.n6951 gnd.n6950 9.3005
R11570 gnd.n355 gnd.n354 9.3005
R11571 gnd.n6958 gnd.n6957 9.3005
R11572 gnd.n6959 gnd.n353 9.3005
R11573 gnd.n6961 gnd.n6960 9.3005
R11574 gnd.n349 gnd.n348 9.3005
R11575 gnd.n6968 gnd.n6967 9.3005
R11576 gnd.n6969 gnd.n347 9.3005
R11577 gnd.n6971 gnd.n6970 9.3005
R11578 gnd.n343 gnd.n342 9.3005
R11579 gnd.n6978 gnd.n6977 9.3005
R11580 gnd.n6979 gnd.n341 9.3005
R11581 gnd.n6981 gnd.n6980 9.3005
R11582 gnd.n337 gnd.n336 9.3005
R11583 gnd.n6988 gnd.n6987 9.3005
R11584 gnd.n6989 gnd.n335 9.3005
R11585 gnd.n6991 gnd.n6990 9.3005
R11586 gnd.n331 gnd.n330 9.3005
R11587 gnd.n6998 gnd.n6997 9.3005
R11588 gnd.n6999 gnd.n329 9.3005
R11589 gnd.n7001 gnd.n7000 9.3005
R11590 gnd.n325 gnd.n324 9.3005
R11591 gnd.n7008 gnd.n7007 9.3005
R11592 gnd.n6798 gnd.n6797 9.3005
R11593 gnd.n7320 gnd.n89 9.3005
R11594 gnd.n7319 gnd.n91 9.3005
R11595 gnd.n96 gnd.n92 9.3005
R11596 gnd.n7314 gnd.n97 9.3005
R11597 gnd.n7313 gnd.n98 9.3005
R11598 gnd.n7312 gnd.n99 9.3005
R11599 gnd.n103 gnd.n100 9.3005
R11600 gnd.n7307 gnd.n104 9.3005
R11601 gnd.n7306 gnd.n105 9.3005
R11602 gnd.n7305 gnd.n106 9.3005
R11603 gnd.n110 gnd.n107 9.3005
R11604 gnd.n7300 gnd.n111 9.3005
R11605 gnd.n7299 gnd.n112 9.3005
R11606 gnd.n7298 gnd.n113 9.3005
R11607 gnd.n117 gnd.n114 9.3005
R11608 gnd.n7293 gnd.n118 9.3005
R11609 gnd.n7292 gnd.n119 9.3005
R11610 gnd.n7288 gnd.n120 9.3005
R11611 gnd.n124 gnd.n121 9.3005
R11612 gnd.n7283 gnd.n125 9.3005
R11613 gnd.n7282 gnd.n126 9.3005
R11614 gnd.n7281 gnd.n127 9.3005
R11615 gnd.n131 gnd.n128 9.3005
R11616 gnd.n7276 gnd.n132 9.3005
R11617 gnd.n7275 gnd.n133 9.3005
R11618 gnd.n7274 gnd.n134 9.3005
R11619 gnd.n138 gnd.n135 9.3005
R11620 gnd.n7269 gnd.n139 9.3005
R11621 gnd.n7268 gnd.n140 9.3005
R11622 gnd.n7267 gnd.n141 9.3005
R11623 gnd.n145 gnd.n142 9.3005
R11624 gnd.n7262 gnd.n146 9.3005
R11625 gnd.n7261 gnd.n147 9.3005
R11626 gnd.n7260 gnd.n148 9.3005
R11627 gnd.n152 gnd.n149 9.3005
R11628 gnd.n7255 gnd.n153 9.3005
R11629 gnd.n7254 gnd.n7253 9.3005
R11630 gnd.n7252 gnd.n156 9.3005
R11631 gnd.n7322 gnd.n7321 9.3005
R11632 gnd.n4151 gnd.n4150 9.3005
R11633 gnd.n4152 gnd.n1594 9.3005
R11634 gnd.n4173 gnd.n4153 9.3005
R11635 gnd.n4172 gnd.n4154 9.3005
R11636 gnd.n4171 gnd.n4155 9.3005
R11637 gnd.n4170 gnd.n4156 9.3005
R11638 gnd.n4169 gnd.n4157 9.3005
R11639 gnd.n4167 gnd.n4158 9.3005
R11640 gnd.n4166 gnd.n4159 9.3005
R11641 gnd.n4163 gnd.n4160 9.3005
R11642 gnd.n4162 gnd.n4161 9.3005
R11643 gnd.n1527 gnd.n1526 9.3005
R11644 gnd.n4263 gnd.n4262 9.3005
R11645 gnd.n4264 gnd.n1525 9.3005
R11646 gnd.n4266 gnd.n4265 9.3005
R11647 gnd.n4267 gnd.n1524 9.3005
R11648 gnd.n4271 gnd.n4270 9.3005
R11649 gnd.n4272 gnd.n1523 9.3005
R11650 gnd.n4296 gnd.n4273 9.3005
R11651 gnd.n4295 gnd.n4274 9.3005
R11652 gnd.n4294 gnd.n4275 9.3005
R11653 gnd.n4293 gnd.n4276 9.3005
R11654 gnd.n4287 gnd.n4277 9.3005
R11655 gnd.n4286 gnd.n4278 9.3005
R11656 gnd.n4285 gnd.n4279 9.3005
R11657 gnd.n4284 gnd.n4281 9.3005
R11658 gnd.n4280 gnd.n263 9.3005
R11659 gnd.n7082 gnd.n264 9.3005
R11660 gnd.n7081 gnd.n265 9.3005
R11661 gnd.n7080 gnd.n266 9.3005
R11662 gnd.n7077 gnd.n267 9.3005
R11663 gnd.n7076 gnd.n268 9.3005
R11664 gnd.n7047 gnd.n269 9.3005
R11665 gnd.n7051 gnd.n7050 9.3005
R11666 gnd.n7052 gnd.n7046 9.3005
R11667 gnd.n7063 gnd.n7053 9.3005
R11668 gnd.n7062 gnd.n7054 9.3005
R11669 gnd.n7061 gnd.n7055 9.3005
R11670 gnd.n7058 gnd.n7057 9.3005
R11671 gnd.n7056 gnd.n160 9.3005
R11672 gnd.n7249 gnd.n159 9.3005
R11673 gnd.n7251 gnd.n7250 9.3005
R11674 gnd.n1596 gnd.n1595 9.3005
R11675 gnd.n1918 gnd.n1917 9.3005
R11676 gnd.n1911 gnd.n1906 9.3005
R11677 gnd.n1924 gnd.n1905 9.3005
R11678 gnd.n1925 gnd.n1904 9.3005
R11679 gnd.n1926 gnd.n1903 9.3005
R11680 gnd.n1902 gnd.n1900 9.3005
R11681 gnd.n1932 gnd.n1899 9.3005
R11682 gnd.n1933 gnd.n1898 9.3005
R11683 gnd.n1934 gnd.n1897 9.3005
R11684 gnd.n1896 gnd.n1894 9.3005
R11685 gnd.n1940 gnd.n1893 9.3005
R11686 gnd.n1941 gnd.n1892 9.3005
R11687 gnd.n1942 gnd.n1891 9.3005
R11688 gnd.n1890 gnd.n1888 9.3005
R11689 gnd.n1948 gnd.n1887 9.3005
R11690 gnd.n1949 gnd.n1886 9.3005
R11691 gnd.n1950 gnd.n1885 9.3005
R11692 gnd.n1884 gnd.n1882 9.3005
R11693 gnd.n1956 gnd.n1881 9.3005
R11694 gnd.n1877 gnd.n1822 9.3005
R11695 gnd.n1876 gnd.n1875 9.3005
R11696 gnd.n1825 gnd.n1824 9.3005
R11697 gnd.n1866 gnd.n1828 9.3005
R11698 gnd.n1868 gnd.n1867 9.3005
R11699 gnd.n1865 gnd.n1830 9.3005
R11700 gnd.n1864 gnd.n1863 9.3005
R11701 gnd.n1832 gnd.n1831 9.3005
R11702 gnd.n1857 gnd.n1856 9.3005
R11703 gnd.n1855 gnd.n1834 9.3005
R11704 gnd.n1854 gnd.n1853 9.3005
R11705 gnd.n1836 gnd.n1835 9.3005
R11706 gnd.n1847 gnd.n1846 9.3005
R11707 gnd.n1845 gnd.n1838 9.3005
R11708 gnd.n1844 gnd.n1843 9.3005
R11709 gnd.n1840 gnd.n1839 9.3005
R11710 gnd.n1916 gnd.n1910 9.3005
R11711 gnd.n1915 gnd.n1914 9.3005
R11712 gnd.n4358 gnd.n1467 9.3005
R11713 gnd.n4357 gnd.n1468 9.3005
R11714 gnd.n1582 gnd.n1469 9.3005
R11715 gnd.n1584 gnd.n1583 9.3005
R11716 gnd.n1562 gnd.n1561 9.3005
R11717 gnd.n4200 gnd.n4199 9.3005
R11718 gnd.n4201 gnd.n1560 9.3005
R11719 gnd.n4205 gnd.n4202 9.3005
R11720 gnd.n4204 gnd.n4203 9.3005
R11721 gnd.n1537 gnd.n1536 9.3005
R11722 gnd.n4253 gnd.n4252 9.3005
R11723 gnd.n4254 gnd.n1535 9.3005
R11724 gnd.n4258 gnd.n4255 9.3005
R11725 gnd.n4257 gnd.n4256 9.3005
R11726 gnd.n1501 gnd.n224 9.3005
R11727 gnd.n7120 gnd.n7119 9.3005
R11728 gnd.n209 gnd.n208 9.3005
R11729 gnd.n7133 gnd.n7132 9.3005
R11730 gnd.n7134 gnd.n207 9.3005
R11731 gnd.n7136 gnd.n7135 9.3005
R11732 gnd.n193 gnd.n192 9.3005
R11733 gnd.n7149 gnd.n7148 9.3005
R11734 gnd.n7150 gnd.n191 9.3005
R11735 gnd.n7152 gnd.n7151 9.3005
R11736 gnd.n177 gnd.n176 9.3005
R11737 gnd.n7165 gnd.n7164 9.3005
R11738 gnd.n7166 gnd.n175 9.3005
R11739 gnd.n7170 gnd.n7167 9.3005
R11740 gnd.n7169 gnd.n7168 9.3005
R11741 gnd.n88 gnd.n87 9.3005
R11742 gnd.n7324 gnd.n7323 9.3005
R11743 gnd.n4359 gnd.n1466 9.3005
R11744 gnd.n7118 gnd.n223 9.3005
R11745 gnd.n2900 gnd.n2600 9.3005
R11746 gnd.n2904 gnd.n2901 9.3005
R11747 gnd.n2903 gnd.n2902 9.3005
R11748 gnd.n2575 gnd.n2574 9.3005
R11749 gnd.n2964 gnd.n2963 9.3005
R11750 gnd.n2965 gnd.n2573 9.3005
R11751 gnd.n2967 gnd.n2966 9.3005
R11752 gnd.n2571 gnd.n2570 9.3005
R11753 gnd.n2972 gnd.n2971 9.3005
R11754 gnd.n2973 gnd.n2569 9.3005
R11755 gnd.n2975 gnd.n2974 9.3005
R11756 gnd.n2567 gnd.n2566 9.3005
R11757 gnd.n2980 gnd.n2979 9.3005
R11758 gnd.n2981 gnd.n2565 9.3005
R11759 gnd.n2983 gnd.n2982 9.3005
R11760 gnd.n2563 gnd.n2562 9.3005
R11761 gnd.n2988 gnd.n2987 9.3005
R11762 gnd.n2989 gnd.n2561 9.3005
R11763 gnd.n2991 gnd.n2990 9.3005
R11764 gnd.n2557 gnd.n2556 9.3005
R11765 gnd.n3131 gnd.n3130 9.3005
R11766 gnd.n3132 gnd.n2555 9.3005
R11767 gnd.n3134 gnd.n3133 9.3005
R11768 gnd.n2551 gnd.n2550 9.3005
R11769 gnd.n3145 gnd.n3144 9.3005
R11770 gnd.n3146 gnd.n2549 9.3005
R11771 gnd.n3148 gnd.n3147 9.3005
R11772 gnd.n2543 gnd.n2542 9.3005
R11773 gnd.n3159 gnd.n3158 9.3005
R11774 gnd.n3160 gnd.n2541 9.3005
R11775 gnd.n3162 gnd.n3161 9.3005
R11776 gnd.n2535 gnd.n2534 9.3005
R11777 gnd.n3173 gnd.n3172 9.3005
R11778 gnd.n3174 gnd.n2533 9.3005
R11779 gnd.n3176 gnd.n3175 9.3005
R11780 gnd.n2258 gnd.n2257 9.3005
R11781 gnd.n3362 gnd.n3361 9.3005
R11782 gnd.n3363 gnd.n2256 9.3005
R11783 gnd.n3365 gnd.n3364 9.3005
R11784 gnd.n2240 gnd.n2239 9.3005
R11785 gnd.n3453 gnd.n3452 9.3005
R11786 gnd.n3454 gnd.n2238 9.3005
R11787 gnd.n3456 gnd.n3455 9.3005
R11788 gnd.n2219 gnd.n2218 9.3005
R11789 gnd.n3484 gnd.n3483 9.3005
R11790 gnd.n3485 gnd.n2217 9.3005
R11791 gnd.n3487 gnd.n3486 9.3005
R11792 gnd.n2197 gnd.n2196 9.3005
R11793 gnd.n3512 gnd.n3511 9.3005
R11794 gnd.n3513 gnd.n2195 9.3005
R11795 gnd.n3517 gnd.n3514 9.3005
R11796 gnd.n3516 gnd.n3515 9.3005
R11797 gnd.n2168 gnd.n2167 9.3005
R11798 gnd.n3549 gnd.n3548 9.3005
R11799 gnd.n3550 gnd.n2166 9.3005
R11800 gnd.n3552 gnd.n3551 9.3005
R11801 gnd.n2145 gnd.n2144 9.3005
R11802 gnd.n3577 gnd.n3576 9.3005
R11803 gnd.n3578 gnd.n2143 9.3005
R11804 gnd.n3582 gnd.n3579 9.3005
R11805 gnd.n3581 gnd.n3580 9.3005
R11806 gnd.n2116 gnd.n2115 9.3005
R11807 gnd.n3628 gnd.n3627 9.3005
R11808 gnd.n3629 gnd.n2114 9.3005
R11809 gnd.n3631 gnd.n3630 9.3005
R11810 gnd.n2095 gnd.n2094 9.3005
R11811 gnd.n3658 gnd.n3657 9.3005
R11812 gnd.n3659 gnd.n2093 9.3005
R11813 gnd.n3663 gnd.n3660 9.3005
R11814 gnd.n3662 gnd.n3661 9.3005
R11815 gnd.n2065 gnd.n2064 9.3005
R11816 gnd.n3708 gnd.n3707 9.3005
R11817 gnd.n3709 gnd.n2063 9.3005
R11818 gnd.n3711 gnd.n3710 9.3005
R11819 gnd.n2042 gnd.n2041 9.3005
R11820 gnd.n3748 gnd.n3747 9.3005
R11821 gnd.n3749 gnd.n2040 9.3005
R11822 gnd.n3751 gnd.n3750 9.3005
R11823 gnd.n2019 gnd.n2018 9.3005
R11824 gnd.n3787 gnd.n3786 9.3005
R11825 gnd.n3788 gnd.n2017 9.3005
R11826 gnd.n3790 gnd.n3789 9.3005
R11827 gnd.n1997 gnd.n1996 9.3005
R11828 gnd.n3828 gnd.n3827 9.3005
R11829 gnd.n3829 gnd.n1995 9.3005
R11830 gnd.n3831 gnd.n3830 9.3005
R11831 gnd.n1975 gnd.n1974 9.3005
R11832 gnd.n3873 gnd.n3872 9.3005
R11833 gnd.n3874 gnd.n1973 9.3005
R11834 gnd.n3882 gnd.n3875 9.3005
R11835 gnd.n3881 gnd.n3876 9.3005
R11836 gnd.n3880 gnd.n3877 9.3005
R11837 gnd.n1779 gnd.n1778 9.3005
R11838 gnd.n4064 gnd.n4063 9.3005
R11839 gnd.n4065 gnd.n1777 9.3005
R11840 gnd.n4067 gnd.n4066 9.3005
R11841 gnd.n1767 gnd.n1766 9.3005
R11842 gnd.n4085 gnd.n4084 9.3005
R11843 gnd.n4086 gnd.n1765 9.3005
R11844 gnd.n4088 gnd.n4087 9.3005
R11845 gnd.n1755 gnd.n1754 9.3005
R11846 gnd.n4108 gnd.n4107 9.3005
R11847 gnd.n4109 gnd.n1753 9.3005
R11848 gnd.n4112 gnd.n4111 9.3005
R11849 gnd.n4110 gnd.n1444 9.3005
R11850 gnd.n4374 gnd.n1445 9.3005
R11851 gnd.n4373 gnd.n1446 9.3005
R11852 gnd.n4372 gnd.n1447 9.3005
R11853 gnd.n1453 gnd.n1448 9.3005
R11854 gnd.n4366 gnd.n1454 9.3005
R11855 gnd.n4365 gnd.n1455 9.3005
R11856 gnd.n4364 gnd.n1456 9.3005
R11857 gnd.n1576 gnd.n1457 9.3005
R11858 gnd.n1577 gnd.n1575 9.3005
R11859 gnd.n1579 gnd.n1578 9.3005
R11860 gnd.n1573 gnd.n1572 9.3005
R11861 gnd.n4189 gnd.n4188 9.3005
R11862 gnd.n4190 gnd.n1571 9.3005
R11863 gnd.n4194 gnd.n4191 9.3005
R11864 gnd.n4193 gnd.n4192 9.3005
R11865 gnd.n1546 gnd.n1545 9.3005
R11866 gnd.n4226 gnd.n4225 9.3005
R11867 gnd.n4227 gnd.n1544 9.3005
R11868 gnd.n4246 gnd.n4228 9.3005
R11869 gnd.n4245 gnd.n4229 9.3005
R11870 gnd.n4244 gnd.n4230 9.3005
R11871 gnd.n4233 gnd.n4231 9.3005
R11872 gnd.n4240 gnd.n4234 9.3005
R11873 gnd.n7088 gnd.n260 9.3005
R11874 gnd.n274 gnd.n261 9.3005
R11875 gnd.n276 gnd.n275 9.3005
R11876 gnd.n277 gnd.n273 9.3005
R11877 gnd.n281 gnd.n280 9.3005
R11878 gnd.n282 gnd.n272 9.3005
R11879 gnd.n7071 gnd.n283 9.3005
R11880 gnd.n7070 gnd.n284 9.3005
R11881 gnd.n7069 gnd.n285 9.3005
R11882 gnd.n288 gnd.n286 9.3005
R11883 gnd.n7044 gnd.n289 9.3005
R11884 gnd.n7043 gnd.n290 9.3005
R11885 gnd.n7042 gnd.n291 9.3005
R11886 gnd.n294 gnd.n292 9.3005
R11887 gnd.n7038 gnd.n295 9.3005
R11888 gnd.n7037 gnd.n296 9.3005
R11889 gnd.n7036 gnd.n297 9.3005
R11890 gnd.n304 gnd.n298 9.3005
R11891 gnd.n305 gnd.n300 9.3005
R11892 gnd.n306 gnd.n303 9.3005
R11893 gnd.n7027 gnd.n307 9.3005
R11894 gnd.n7026 gnd.n308 9.3005
R11895 gnd.n7025 gnd.n309 9.3005
R11896 gnd.n314 gnd.n310 9.3005
R11897 gnd.n7019 gnd.n315 9.3005
R11898 gnd.n7018 gnd.n316 9.3005
R11899 gnd.n7017 gnd.n317 9.3005
R11900 gnd.n322 gnd.n318 9.3005
R11901 gnd.n7011 gnd.n323 9.3005
R11902 gnd.n7010 gnd.n7009 9.3005
R11903 gnd.n2852 gnd.n2851 9.3005
R11904 gnd.n2730 gnd.n2670 9.3005
R11905 gnd.n2751 gnd.n2731 9.3005
R11906 gnd.n2750 gnd.n2732 9.3005
R11907 gnd.n2749 gnd.n2733 9.3005
R11908 gnd.n2737 gnd.n2734 9.3005
R11909 gnd.n2736 gnd.n2735 9.3005
R11910 gnd.n2651 gnd.n2650 9.3005
R11911 gnd.n2811 gnd.n2810 9.3005
R11912 gnd.n2812 gnd.n2649 9.3005
R11913 gnd.n2814 gnd.n2813 9.3005
R11914 gnd.n2644 gnd.n2643 9.3005
R11915 gnd.n2828 gnd.n2827 9.3005
R11916 gnd.n2829 gnd.n2642 9.3005
R11917 gnd.n2834 gnd.n2830 9.3005
R11918 gnd.n2833 gnd.n2832 9.3005
R11919 gnd.n2831 gnd.n2614 9.3005
R11920 gnd.n2891 gnd.n2615 9.3005
R11921 gnd.n2890 gnd.n2616 9.3005
R11922 gnd.n2889 gnd.n2617 9.3005
R11923 gnd.n2850 gnd.n2618 9.3005
R11924 gnd.n2729 gnd.n2728 9.3005
R11925 gnd.n2724 gnd.n2723 9.3005
R11926 gnd.n2722 gnd.n2675 9.3005
R11927 gnd.n2721 gnd.n2720 9.3005
R11928 gnd.n2717 gnd.n2678 9.3005
R11929 gnd.n2716 gnd.n2713 9.3005
R11930 gnd.n2712 gnd.n2679 9.3005
R11931 gnd.n2711 gnd.n2710 9.3005
R11932 gnd.n2707 gnd.n2680 9.3005
R11933 gnd.n2706 gnd.n2703 9.3005
R11934 gnd.n2702 gnd.n2681 9.3005
R11935 gnd.n2701 gnd.n2700 9.3005
R11936 gnd.n2697 gnd.n2682 9.3005
R11937 gnd.n2696 gnd.n2693 9.3005
R11938 gnd.n2692 gnd.n2683 9.3005
R11939 gnd.n2691 gnd.n2690 9.3005
R11940 gnd.n2687 gnd.n2684 9.3005
R11941 gnd.n2686 gnd.n2685 9.3005
R11942 gnd.n2725 gnd.n2671 9.3005
R11943 gnd.n2727 gnd.n2726 9.3005
R11944 gnd.n4632 gnd.n4631 9.3005
R11945 gnd.n4630 gnd.n1125 9.3005
R11946 gnd.n4629 gnd.n4628 9.3005
R11947 gnd.n1127 gnd.n1126 9.3005
R11948 gnd.n4618 gnd.n1147 9.3005
R11949 gnd.n4617 gnd.n1148 9.3005
R11950 gnd.n4616 gnd.n1149 9.3005
R11951 gnd.n1166 gnd.n1150 9.3005
R11952 gnd.n4606 gnd.n1167 9.3005
R11953 gnd.n4605 gnd.n1168 9.3005
R11954 gnd.n4604 gnd.n1169 9.3005
R11955 gnd.n1188 gnd.n1170 9.3005
R11956 gnd.n4594 gnd.n1189 9.3005
R11957 gnd.n4593 gnd.n1190 9.3005
R11958 gnd.n4592 gnd.n1191 9.3005
R11959 gnd.n1211 gnd.n1192 9.3005
R11960 gnd.n1212 gnd.n1210 9.3005
R11961 gnd.n4580 gnd.n1213 9.3005
R11962 gnd.n4579 gnd.n1214 9.3005
R11963 gnd.n4578 gnd.n1215 9.3005
R11964 gnd.n2636 gnd.n1216 9.3005
R11965 gnd.n4567 gnd.n1229 9.3005
R11966 gnd.n4566 gnd.n1230 9.3005
R11967 gnd.n4565 gnd.n1231 9.3005
R11968 gnd.n1247 gnd.n1232 9.3005
R11969 gnd.n4554 gnd.n1248 9.3005
R11970 gnd.n4553 gnd.n1249 9.3005
R11971 gnd.n4552 gnd.n1250 9.3005
R11972 gnd.n1267 gnd.n1251 9.3005
R11973 gnd.n4542 gnd.n1268 9.3005
R11974 gnd.n4541 gnd.n1269 9.3005
R11975 gnd.n4540 gnd.n1270 9.3005
R11976 gnd.n1289 gnd.n1271 9.3005
R11977 gnd.n4530 gnd.n1290 9.3005
R11978 gnd.n4529 gnd.n1291 9.3005
R11979 gnd.n4528 gnd.n1292 9.3005
R11980 gnd.n1310 gnd.n1293 9.3005
R11981 gnd.n4518 gnd.n1311 9.3005
R11982 gnd.n4517 gnd.n1312 9.3005
R11983 gnd.n4516 gnd.n1313 9.3005
R11984 gnd.n1331 gnd.n1314 9.3005
R11985 gnd.n4506 gnd.n4505 9.3005
R11986 gnd.n4633 gnd.n1124 9.3005
R11987 gnd.n2401 gnd.n2397 9.3005
R11988 gnd.n2434 gnd.n2431 9.3005
R11989 gnd.n2435 gnd.n2430 9.3005
R11990 gnd.n2438 gnd.n2429 9.3005
R11991 gnd.n2439 gnd.n2428 9.3005
R11992 gnd.n2442 gnd.n2427 9.3005
R11993 gnd.n2443 gnd.n2426 9.3005
R11994 gnd.n2446 gnd.n2425 9.3005
R11995 gnd.n2447 gnd.n2424 9.3005
R11996 gnd.n2450 gnd.n2423 9.3005
R11997 gnd.n2451 gnd.n2422 9.3005
R11998 gnd.n2454 gnd.n2421 9.3005
R11999 gnd.n2455 gnd.n2420 9.3005
R12000 gnd.n2456 gnd.n2419 9.3005
R12001 gnd.n2418 gnd.n2415 9.3005
R12002 gnd.n2417 gnd.n2416 9.3005
R12003 gnd.n3281 gnd.n3280 9.3005
R12004 gnd.n2403 gnd.n2402 9.3005
R12005 gnd.n2462 gnd.n2460 9.3005
R12006 gnd.n3273 gnd.n2463 9.3005
R12007 gnd.n3272 gnd.n2464 9.3005
R12008 gnd.n3271 gnd.n2465 9.3005
R12009 gnd.n2469 gnd.n2466 9.3005
R12010 gnd.n3266 gnd.n2470 9.3005
R12011 gnd.n3265 gnd.n2471 9.3005
R12012 gnd.n3264 gnd.n2472 9.3005
R12013 gnd.n2476 gnd.n2473 9.3005
R12014 gnd.n3259 gnd.n2477 9.3005
R12015 gnd.n3258 gnd.n2478 9.3005
R12016 gnd.n3257 gnd.n2479 9.3005
R12017 gnd.n2483 gnd.n2480 9.3005
R12018 gnd.n3252 gnd.n2484 9.3005
R12019 gnd.n3251 gnd.n2485 9.3005
R12020 gnd.n3250 gnd.n2486 9.3005
R12021 gnd.n2491 gnd.n2489 9.3005
R12022 gnd.n3245 gnd.n3244 9.3005
R12023 gnd.n3282 gnd.n2396 9.3005
R12024 gnd.n2740 gnd.n2739 9.3005
R12025 gnd.n2742 gnd.n2741 9.3005
R12026 gnd.n2743 gnd.n2738 9.3005
R12027 gnd.n2745 gnd.n2744 9.3005
R12028 gnd.n2654 gnd.n2653 9.3005
R12029 gnd.n2803 gnd.n2802 9.3005
R12030 gnd.n2804 gnd.n2652 9.3005
R12031 gnd.n2806 gnd.n2805 9.3005
R12032 gnd.n2647 gnd.n2646 9.3005
R12033 gnd.n2819 gnd.n2818 9.3005
R12034 gnd.n2820 gnd.n2645 9.3005
R12035 gnd.n2823 gnd.n2822 9.3005
R12036 gnd.n2821 gnd.n2641 9.3005
R12037 gnd.n2839 gnd.n2640 9.3005
R12038 gnd.n2841 gnd.n2840 9.3005
R12039 gnd.n2842 gnd.n2639 9.3005
R12040 gnd.n2844 gnd.n2843 9.3005
R12041 gnd.n2845 gnd.n2637 9.3005
R12042 gnd.n2847 gnd.n2846 9.3005
R12043 gnd.n2848 gnd.n2635 9.3005
R12044 gnd.n2856 gnd.n2849 9.3005
R12045 gnd.n2857 gnd.n2634 9.3005
R12046 gnd.n2859 gnd.n2858 9.3005
R12047 gnd.n2860 gnd.n2633 9.3005
R12048 gnd.n2866 gnd.n2861 9.3005
R12049 gnd.n2865 gnd.n2862 9.3005
R12050 gnd.n2864 gnd.n2863 9.3005
R12051 gnd.n2593 gnd.n2592 9.3005
R12052 gnd.n2918 gnd.n2917 9.3005
R12053 gnd.n2919 gnd.n2591 9.3005
R12054 gnd.n2921 gnd.n2920 9.3005
R12055 gnd.n2922 gnd.n2590 9.3005
R12056 gnd.n2926 gnd.n2925 9.3005
R12057 gnd.n2927 gnd.n2589 9.3005
R12058 gnd.n2932 gnd.n2928 9.3005
R12059 gnd.n2933 gnd.n2588 9.3005
R12060 gnd.n2937 gnd.n2936 9.3005
R12061 gnd.n2938 gnd.n2587 9.3005
R12062 gnd.n2941 gnd.n2940 9.3005
R12063 gnd.n2939 gnd.n2493 9.3005
R12064 gnd.n3241 gnd.n2492 9.3005
R12065 gnd.n3243 gnd.n3242 9.3005
R12066 gnd.n1118 gnd.n1116 9.3005
R12067 gnd.n4642 gnd.n4641 9.3005
R12068 gnd.n4643 gnd.n1110 9.3005
R12069 gnd.n4646 gnd.n1109 9.3005
R12070 gnd.n4647 gnd.n1108 9.3005
R12071 gnd.n4650 gnd.n1107 9.3005
R12072 gnd.n4651 gnd.n1106 9.3005
R12073 gnd.n4654 gnd.n1105 9.3005
R12074 gnd.n4655 gnd.n1104 9.3005
R12075 gnd.n4658 gnd.n1103 9.3005
R12076 gnd.n4659 gnd.n1102 9.3005
R12077 gnd.n4662 gnd.n1101 9.3005
R12078 gnd.n4663 gnd.n1100 9.3005
R12079 gnd.n4666 gnd.n1099 9.3005
R12080 gnd.n4667 gnd.n1098 9.3005
R12081 gnd.n4670 gnd.n1097 9.3005
R12082 gnd.n4671 gnd.n1096 9.3005
R12083 gnd.n4674 gnd.n1095 9.3005
R12084 gnd.n4675 gnd.n1094 9.3005
R12085 gnd.n4678 gnd.n1093 9.3005
R12086 gnd.n4680 gnd.n1090 9.3005
R12087 gnd.n4683 gnd.n1089 9.3005
R12088 gnd.n4684 gnd.n1088 9.3005
R12089 gnd.n4687 gnd.n1087 9.3005
R12090 gnd.n4688 gnd.n1086 9.3005
R12091 gnd.n4691 gnd.n1085 9.3005
R12092 gnd.n4692 gnd.n1084 9.3005
R12093 gnd.n4695 gnd.n1083 9.3005
R12094 gnd.n4696 gnd.n1082 9.3005
R12095 gnd.n4699 gnd.n1081 9.3005
R12096 gnd.n4700 gnd.n1080 9.3005
R12097 gnd.n4703 gnd.n1079 9.3005
R12098 gnd.n4704 gnd.n1078 9.3005
R12099 gnd.n4707 gnd.n1077 9.3005
R12100 gnd.n4709 gnd.n1076 9.3005
R12101 gnd.n4710 gnd.n1075 9.3005
R12102 gnd.n4711 gnd.n1074 9.3005
R12103 gnd.n4712 gnd.n1073 9.3005
R12104 gnd.n4640 gnd.n1115 9.3005
R12105 gnd.n4639 gnd.n4638 9.3005
R12106 gnd.n2665 gnd.n2664 9.3005
R12107 gnd.n2663 gnd.n1136 9.3005
R12108 gnd.n4624 gnd.n1137 9.3005
R12109 gnd.n4623 gnd.n1138 9.3005
R12110 gnd.n4622 gnd.n1139 9.3005
R12111 gnd.n1156 gnd.n1140 9.3005
R12112 gnd.n4612 gnd.n1157 9.3005
R12113 gnd.n4611 gnd.n1158 9.3005
R12114 gnd.n4610 gnd.n1159 9.3005
R12115 gnd.n1177 gnd.n1160 9.3005
R12116 gnd.n4600 gnd.n1178 9.3005
R12117 gnd.n4599 gnd.n1179 9.3005
R12118 gnd.n4598 gnd.n1180 9.3005
R12119 gnd.n1198 gnd.n1181 9.3005
R12120 gnd.n4588 gnd.n1199 9.3005
R12121 gnd.n1257 gnd.n1240 9.3005
R12122 gnd.n4548 gnd.n1258 9.3005
R12123 gnd.n4547 gnd.n1259 9.3005
R12124 gnd.n4546 gnd.n1260 9.3005
R12125 gnd.n1278 gnd.n1261 9.3005
R12126 gnd.n4536 gnd.n1279 9.3005
R12127 gnd.n4535 gnd.n1280 9.3005
R12128 gnd.n4534 gnd.n1281 9.3005
R12129 gnd.n1299 gnd.n1282 9.3005
R12130 gnd.n4524 gnd.n1300 9.3005
R12131 gnd.n4523 gnd.n1301 9.3005
R12132 gnd.n4522 gnd.n1302 9.3005
R12133 gnd.n1321 gnd.n1303 9.3005
R12134 gnd.n4512 gnd.n1322 9.3005
R12135 gnd.n4511 gnd.n1323 9.3005
R12136 gnd.n4510 gnd.n1324 9.3005
R12137 gnd.n2662 gnd.n2661 9.3005
R12138 gnd.n4558 gnd.n1200 9.3005
R12139 gnd.n4736 gnd.n1021 9.3005
R12140 gnd.n4735 gnd.n1022 9.3005
R12141 gnd.n1027 gnd.n1023 9.3005
R12142 gnd.n4729 gnd.n1028 9.3005
R12143 gnd.n4728 gnd.n1029 9.3005
R12144 gnd.n4727 gnd.n1030 9.3005
R12145 gnd.n1035 gnd.n1031 9.3005
R12146 gnd.n4721 gnd.n1036 9.3005
R12147 gnd.n4720 gnd.n1037 9.3005
R12148 gnd.n4719 gnd.n1038 9.3005
R12149 gnd.n2759 gnd.n1039 9.3005
R12150 gnd.n2761 gnd.n2760 9.3005
R12151 gnd.n2758 gnd.n2757 9.3005
R12152 gnd.n2766 gnd.n2765 9.3005
R12153 gnd.n2767 gnd.n2756 9.3005
R12154 gnd.n2769 gnd.n2768 9.3005
R12155 gnd.n2660 gnd.n2659 9.3005
R12156 gnd.n2774 gnd.n2773 9.3005
R12157 gnd.n2775 gnd.n2658 9.3005
R12158 gnd.n2797 gnd.n2776 9.3005
R12159 gnd.n2796 gnd.n2777 9.3005
R12160 gnd.n2795 gnd.n2778 9.3005
R12161 gnd.n2781 gnd.n2779 9.3005
R12162 gnd.n2791 gnd.n2782 9.3005
R12163 gnd.n2790 gnd.n2783 9.3005
R12164 gnd.n2789 gnd.n2784 9.3005
R12165 gnd.n2786 gnd.n2785 9.3005
R12166 gnd.n2607 gnd.n2606 9.3005
R12167 gnd.n2898 gnd.n2897 9.3005
R12168 gnd.n4737 gnd.n1020 9.3005
R12169 gnd.n6108 gnd.n928 9.3005
R12170 gnd.n6109 gnd.n927 9.3005
R12171 gnd.n6110 gnd.n926 9.3005
R12172 gnd.n925 gnd.n921 9.3005
R12173 gnd.n6116 gnd.n920 9.3005
R12174 gnd.n6117 gnd.n919 9.3005
R12175 gnd.n6118 gnd.n918 9.3005
R12176 gnd.n917 gnd.n913 9.3005
R12177 gnd.n6124 gnd.n912 9.3005
R12178 gnd.n6125 gnd.n911 9.3005
R12179 gnd.n6126 gnd.n910 9.3005
R12180 gnd.n909 gnd.n905 9.3005
R12181 gnd.n6132 gnd.n904 9.3005
R12182 gnd.n6133 gnd.n903 9.3005
R12183 gnd.n6134 gnd.n902 9.3005
R12184 gnd.n901 gnd.n897 9.3005
R12185 gnd.n6140 gnd.n896 9.3005
R12186 gnd.n6141 gnd.n895 9.3005
R12187 gnd.n6142 gnd.n894 9.3005
R12188 gnd.n893 gnd.n889 9.3005
R12189 gnd.n6148 gnd.n888 9.3005
R12190 gnd.n6149 gnd.n887 9.3005
R12191 gnd.n6150 gnd.n886 9.3005
R12192 gnd.n885 gnd.n881 9.3005
R12193 gnd.n6156 gnd.n880 9.3005
R12194 gnd.n6157 gnd.n879 9.3005
R12195 gnd.n6158 gnd.n878 9.3005
R12196 gnd.n877 gnd.n873 9.3005
R12197 gnd.n6164 gnd.n872 9.3005
R12198 gnd.n6165 gnd.n871 9.3005
R12199 gnd.n6166 gnd.n870 9.3005
R12200 gnd.n869 gnd.n865 9.3005
R12201 gnd.n6172 gnd.n864 9.3005
R12202 gnd.n6173 gnd.n863 9.3005
R12203 gnd.n6174 gnd.n862 9.3005
R12204 gnd.n861 gnd.n857 9.3005
R12205 gnd.n6180 gnd.n856 9.3005
R12206 gnd.n6181 gnd.n855 9.3005
R12207 gnd.n6182 gnd.n854 9.3005
R12208 gnd.n853 gnd.n849 9.3005
R12209 gnd.n6188 gnd.n848 9.3005
R12210 gnd.n6189 gnd.n847 9.3005
R12211 gnd.n6190 gnd.n846 9.3005
R12212 gnd.n845 gnd.n841 9.3005
R12213 gnd.n6196 gnd.n840 9.3005
R12214 gnd.n6197 gnd.n839 9.3005
R12215 gnd.n6198 gnd.n838 9.3005
R12216 gnd.n837 gnd.n833 9.3005
R12217 gnd.n6204 gnd.n832 9.3005
R12218 gnd.n6205 gnd.n831 9.3005
R12219 gnd.n6206 gnd.n830 9.3005
R12220 gnd.n829 gnd.n825 9.3005
R12221 gnd.n6212 gnd.n824 9.3005
R12222 gnd.n6213 gnd.n823 9.3005
R12223 gnd.n6214 gnd.n822 9.3005
R12224 gnd.n821 gnd.n817 9.3005
R12225 gnd.n6220 gnd.n816 9.3005
R12226 gnd.n6221 gnd.n815 9.3005
R12227 gnd.n6222 gnd.n814 9.3005
R12228 gnd.n813 gnd.n809 9.3005
R12229 gnd.n6228 gnd.n808 9.3005
R12230 gnd.n6229 gnd.n807 9.3005
R12231 gnd.n6230 gnd.n806 9.3005
R12232 gnd.n805 gnd.n801 9.3005
R12233 gnd.n6236 gnd.n800 9.3005
R12234 gnd.n6237 gnd.n799 9.3005
R12235 gnd.n6238 gnd.n798 9.3005
R12236 gnd.n797 gnd.n793 9.3005
R12237 gnd.n6244 gnd.n792 9.3005
R12238 gnd.n6245 gnd.n791 9.3005
R12239 gnd.n6246 gnd.n790 9.3005
R12240 gnd.n789 gnd.n785 9.3005
R12241 gnd.n6252 gnd.n784 9.3005
R12242 gnd.n6253 gnd.n783 9.3005
R12243 gnd.n6254 gnd.n782 9.3005
R12244 gnd.n781 gnd.n777 9.3005
R12245 gnd.n6260 gnd.n776 9.3005
R12246 gnd.n6261 gnd.n775 9.3005
R12247 gnd.n6262 gnd.n774 9.3005
R12248 gnd.n773 gnd.n769 9.3005
R12249 gnd.n6268 gnd.n768 9.3005
R12250 gnd.n6269 gnd.n767 9.3005
R12251 gnd.n6270 gnd.n766 9.3005
R12252 gnd.n765 gnd.n761 9.3005
R12253 gnd.n1019 gnd.n929 9.3005
R12254 gnd.n1658 gnd.n1657 9.3005
R12255 gnd.n1638 gnd.n1636 9.3005
R12256 gnd.n1665 gnd.n1664 9.3005
R12257 gnd.n1632 gnd.n1631 9.3005
R12258 gnd.n1677 gnd.n1676 9.3005
R12259 gnd.n1629 gnd.n1627 9.3005
R12260 gnd.n1684 gnd.n1683 9.3005
R12261 gnd.n1623 gnd.n1622 9.3005
R12262 gnd.n1696 gnd.n1695 9.3005
R12263 gnd.n1620 gnd.n1618 9.3005
R12264 gnd.n1703 gnd.n1702 9.3005
R12265 gnd.n1614 gnd.n1613 9.3005
R12266 gnd.n1715 gnd.n1714 9.3005
R12267 gnd.n1611 gnd.n1609 9.3005
R12268 gnd.n1722 gnd.n1721 9.3005
R12269 gnd.n1603 gnd.n1602 9.3005
R12270 gnd.n1732 gnd.n1731 9.3005
R12271 gnd.n1600 gnd.n1598 9.3005
R12272 gnd.n1641 gnd.n1640 9.3005
R12273 gnd.n1724 gnd.n1723 9.3005
R12274 gnd.n1713 gnd.n1608 9.3005
R12275 gnd.n1712 gnd.n1711 9.3005
R12276 gnd.n1619 gnd.n1615 9.3005
R12277 gnd.n1705 gnd.n1704 9.3005
R12278 gnd.n1694 gnd.n1617 9.3005
R12279 gnd.n1693 gnd.n1692 9.3005
R12280 gnd.n1628 gnd.n1624 9.3005
R12281 gnd.n1686 gnd.n1685 9.3005
R12282 gnd.n1675 gnd.n1626 9.3005
R12283 gnd.n1674 gnd.n1673 9.3005
R12284 gnd.n1637 gnd.n1633 9.3005
R12285 gnd.n1667 gnd.n1666 9.3005
R12286 gnd.n1656 gnd.n1635 9.3005
R12287 gnd.n1655 gnd.n1654 9.3005
R12288 gnd.n1643 gnd.n1642 9.3005
R12289 gnd.n1610 gnd.n1606 9.3005
R12290 gnd.n1730 gnd.n1729 9.3005
R12291 gnd.n4142 gnd.n4141 9.3005
R12292 gnd.n4140 gnd.n1599 9.3005
R12293 gnd.n4139 gnd.n4138 9.3005
R12294 gnd.n4137 gnd.n1740 9.3005
R12295 gnd.n4136 gnd.n4135 9.3005
R12296 gnd.n4134 gnd.n1741 9.3005
R12297 gnd.n4130 gnd.n4129 9.3005
R12298 gnd.n4128 gnd.n1748 9.3005
R12299 gnd.n4127 gnd.n4126 9.3005
R12300 gnd.n4125 gnd.n4120 9.3005
R12301 gnd.n3214 gnd.n2516 9.3005
R12302 gnd.n3213 gnd.n3212 9.3005
R12303 gnd.n3211 gnd.n2520 9.3005
R12304 gnd.n3210 gnd.n3209 9.3005
R12305 gnd.n3208 gnd.n2521 9.3005
R12306 gnd.n3207 gnd.n3206 9.3005
R12307 gnd.n3205 gnd.n2525 9.3005
R12308 gnd.n3204 gnd.n3203 9.3005
R12309 gnd.n3202 gnd.n2526 9.3005
R12310 gnd.n3201 gnd.n3200 9.3005
R12311 gnd.n3199 gnd.n2530 9.3005
R12312 gnd.n3198 gnd.n3197 9.3005
R12313 gnd.n3196 gnd.n2531 9.3005
R12314 gnd.n3195 gnd.n3194 9.3005
R12315 gnd.n3193 gnd.n3185 9.3005
R12316 gnd.n3192 gnd.n3191 9.3005
R12317 gnd.n3190 gnd.n3186 9.3005
R12318 gnd.n2232 gnd.n2231 9.3005
R12319 gnd.n3463 gnd.n3462 9.3005
R12320 gnd.n3464 gnd.n2230 9.3005
R12321 gnd.n3466 gnd.n3465 9.3005
R12322 gnd.n2212 gnd.n2211 9.3005
R12323 gnd.n3494 gnd.n3493 9.3005
R12324 gnd.n3495 gnd.n2209 9.3005
R12325 gnd.n3498 gnd.n3497 9.3005
R12326 gnd.n3496 gnd.n2210 9.3005
R12327 gnd.n2182 gnd.n2181 9.3005
R12328 gnd.n3530 gnd.n3529 9.3005
R12329 gnd.n3531 gnd.n2180 9.3005
R12330 gnd.n3533 gnd.n3532 9.3005
R12331 gnd.n2161 gnd.n2160 9.3005
R12332 gnd.n3558 gnd.n3557 9.3005
R12333 gnd.n3559 gnd.n2158 9.3005
R12334 gnd.n3562 gnd.n3561 9.3005
R12335 gnd.n3560 gnd.n2159 9.3005
R12336 gnd.n2131 gnd.n2130 9.3005
R12337 gnd.n3596 gnd.n3595 9.3005
R12338 gnd.n3597 gnd.n2128 9.3005
R12339 gnd.n3614 gnd.n3613 9.3005
R12340 gnd.n3612 gnd.n2129 9.3005
R12341 gnd.n3611 gnd.n3610 9.3005
R12342 gnd.n3609 gnd.n3598 9.3005
R12343 gnd.n3608 gnd.n3607 9.3005
R12344 gnd.n3606 gnd.n3602 9.3005
R12345 gnd.n3605 gnd.n3604 9.3005
R12346 gnd.n3603 gnd.n2081 9.3005
R12347 gnd.n3678 gnd.n2080 9.3005
R12348 gnd.n3680 gnd.n3679 9.3005
R12349 gnd.n3681 gnd.n2079 9.3005
R12350 gnd.n3683 gnd.n3682 9.3005
R12351 gnd.n2057 gnd.n2055 9.3005
R12352 gnd.n3732 gnd.n3731 9.3005
R12353 gnd.n3730 gnd.n2056 9.3005
R12354 gnd.n3729 gnd.n3728 9.3005
R12355 gnd.n2034 gnd.n2032 9.3005
R12356 gnd.n3772 gnd.n3771 9.3005
R12357 gnd.n3770 gnd.n2033 9.3005
R12358 gnd.n3769 gnd.n3768 9.3005
R12359 gnd.n2012 gnd.n2010 9.3005
R12360 gnd.n3811 gnd.n3810 9.3005
R12361 gnd.n3809 gnd.n2011 9.3005
R12362 gnd.n3808 gnd.n3807 9.3005
R12363 gnd.n1988 gnd.n1986 9.3005
R12364 gnd.n3859 gnd.n3858 9.3005
R12365 gnd.n3857 gnd.n1987 9.3005
R12366 gnd.n3856 gnd.n3855 9.3005
R12367 gnd.n3854 gnd.n1989 9.3005
R12368 gnd.n1784 gnd.n1783 9.3005
R12369 gnd.n4053 gnd.n4052 9.3005
R12370 gnd.n4054 gnd.n1782 9.3005
R12371 gnd.n4056 gnd.n4055 9.3005
R12372 gnd.n1773 gnd.n1772 9.3005
R12373 gnd.n4074 gnd.n4073 9.3005
R12374 gnd.n4075 gnd.n1771 9.3005
R12375 gnd.n4077 gnd.n4076 9.3005
R12376 gnd.n1761 gnd.n1760 9.3005
R12377 gnd.n4095 gnd.n4094 9.3005
R12378 gnd.n4096 gnd.n1759 9.3005
R12379 gnd.n4099 gnd.n4098 9.3005
R12380 gnd.n4097 gnd.n1750 9.3005
R12381 gnd.n4117 gnd.n1749 9.3005
R12382 gnd.n4119 gnd.n4118 9.3005
R12383 gnd.n3216 gnd.n3215 9.3005
R12384 gnd.n3219 gnd.n3218 9.3005
R12385 gnd.n3220 gnd.n2511 9.3005
R12386 gnd.n3222 gnd.n3221 9.3005
R12387 gnd.n3224 gnd.n3223 9.3005
R12388 gnd.n3225 gnd.n2504 9.3005
R12389 gnd.n3227 gnd.n3226 9.3005
R12390 gnd.n3228 gnd.n2503 9.3005
R12391 gnd.n3230 gnd.n3229 9.3005
R12392 gnd.n3231 gnd.n2497 9.3005
R12393 gnd.n3217 gnd.n2515 9.3005
R12394 gnd.n2632 gnd.n2630 9.3005
R12395 gnd.n2874 gnd.n2873 9.3005
R12396 gnd.n2872 gnd.n2631 9.3005
R12397 gnd.n2871 gnd.n2870 9.3005
R12398 gnd.n2596 gnd.n2595 9.3005
R12399 gnd.n2910 gnd.n2909 9.3005
R12400 gnd.n2911 gnd.n2594 9.3005
R12401 gnd.n2913 gnd.n2912 9.3005
R12402 gnd.n2580 gnd.n2578 9.3005
R12403 gnd.n2958 gnd.n2957 9.3005
R12404 gnd.n2956 gnd.n2579 9.3005
R12405 gnd.n2955 gnd.n2954 9.3005
R12406 gnd.n2953 gnd.n2581 9.3005
R12407 gnd.n2952 gnd.n2951 9.3005
R12408 gnd.n2950 gnd.n2584 9.3005
R12409 gnd.n2949 gnd.n2948 9.3005
R12410 gnd.n2947 gnd.n2585 9.3005
R12411 gnd.n2946 gnd.n2945 9.3005
R12412 gnd.n2496 gnd.n2494 9.3005
R12413 gnd.n3237 gnd.n3236 9.3005
R12414 gnd.n3235 gnd.n2495 9.3005
R12415 gnd.n3233 gnd.n3232 9.3005
R12416 gnd.n2499 gnd.n2498 9.3005
R12417 gnd.n3083 gnd.n3082 9.3005
R12418 gnd.n3085 gnd.n3084 9.3005
R12419 gnd.n3063 gnd.n3062 9.3005
R12420 gnd.n3091 gnd.n3090 9.3005
R12421 gnd.n3093 gnd.n3092 9.3005
R12422 gnd.n3053 gnd.n3052 9.3005
R12423 gnd.n3099 gnd.n3098 9.3005
R12424 gnd.n3101 gnd.n3100 9.3005
R12425 gnd.n3040 gnd.n3039 9.3005
R12426 gnd.n3107 gnd.n3106 9.3005
R12427 gnd.n3109 gnd.n3108 9.3005
R12428 gnd.n3030 gnd.n3029 9.3005
R12429 gnd.n3115 gnd.n3114 9.3005
R12430 gnd.n3117 gnd.n3116 9.3005
R12431 gnd.n3015 gnd.n3013 9.3005
R12432 gnd.n3123 gnd.n3122 9.3005
R12433 gnd.n3124 gnd.n3012 9.3005
R12434 gnd.n3017 gnd.n1333 9.3005
R12435 gnd.n3016 gnd.n3014 9.3005
R12436 gnd.n3121 gnd.n3120 9.3005
R12437 gnd.n3119 gnd.n3118 9.3005
R12438 gnd.n3025 gnd.n3024 9.3005
R12439 gnd.n3113 gnd.n3112 9.3005
R12440 gnd.n3111 gnd.n3110 9.3005
R12441 gnd.n3036 gnd.n3035 9.3005
R12442 gnd.n3105 gnd.n3104 9.3005
R12443 gnd.n3103 gnd.n3102 9.3005
R12444 gnd.n3047 gnd.n3046 9.3005
R12445 gnd.n3097 gnd.n3096 9.3005
R12446 gnd.n3095 gnd.n3094 9.3005
R12447 gnd.n3059 gnd.n3058 9.3005
R12448 gnd.n3089 gnd.n3088 9.3005
R12449 gnd.n3087 gnd.n3086 9.3005
R12450 gnd.n3072 gnd.n3071 9.3005
R12451 gnd.n3081 gnd.n3080 9.3005
R12452 gnd.n4500 gnd.n1334 9.3005
R12453 gnd.n4499 gnd.n4498 9.3005
R12454 gnd.n4497 gnd.n1338 9.3005
R12455 gnd.n4496 gnd.n4495 9.3005
R12456 gnd.n4494 gnd.n1339 9.3005
R12457 gnd.n4493 gnd.n4492 9.3005
R12458 gnd.n4491 gnd.n1343 9.3005
R12459 gnd.n4490 gnd.n4489 9.3005
R12460 gnd.n4488 gnd.n1344 9.3005
R12461 gnd.n4487 gnd.n4486 9.3005
R12462 gnd.n4485 gnd.n1348 9.3005
R12463 gnd.n4484 gnd.n4483 9.3005
R12464 gnd.n4482 gnd.n1349 9.3005
R12465 gnd.n4481 gnd.n4480 9.3005
R12466 gnd.n4479 gnd.n1353 9.3005
R12467 gnd.n4478 gnd.n4477 9.3005
R12468 gnd.n4476 gnd.n1354 9.3005
R12469 gnd.n4475 gnd.n4474 9.3005
R12470 gnd.n4473 gnd.n1358 9.3005
R12471 gnd.n4472 gnd.n4471 9.3005
R12472 gnd.n4470 gnd.n1359 9.3005
R12473 gnd.n4469 gnd.n4468 9.3005
R12474 gnd.n4467 gnd.n1363 9.3005
R12475 gnd.n4466 gnd.n4465 9.3005
R12476 gnd.n4464 gnd.n1364 9.3005
R12477 gnd.n4463 gnd.n4462 9.3005
R12478 gnd.n4461 gnd.n1368 9.3005
R12479 gnd.n4460 gnd.n4459 9.3005
R12480 gnd.n4458 gnd.n1369 9.3005
R12481 gnd.n4457 gnd.n4456 9.3005
R12482 gnd.n4455 gnd.n1373 9.3005
R12483 gnd.n4454 gnd.n4453 9.3005
R12484 gnd.n4452 gnd.n1374 9.3005
R12485 gnd.n4451 gnd.n4450 9.3005
R12486 gnd.n4449 gnd.n1378 9.3005
R12487 gnd.n4448 gnd.n4447 9.3005
R12488 gnd.n4446 gnd.n1379 9.3005
R12489 gnd.n4445 gnd.n4444 9.3005
R12490 gnd.n4443 gnd.n1383 9.3005
R12491 gnd.n4442 gnd.n4441 9.3005
R12492 gnd.n4440 gnd.n1384 9.3005
R12493 gnd.n4439 gnd.n4438 9.3005
R12494 gnd.n4437 gnd.n1388 9.3005
R12495 gnd.n4436 gnd.n4435 9.3005
R12496 gnd.n4434 gnd.n1389 9.3005
R12497 gnd.n4433 gnd.n4432 9.3005
R12498 gnd.n4431 gnd.n1393 9.3005
R12499 gnd.n4430 gnd.n4429 9.3005
R12500 gnd.n4428 gnd.n1394 9.3005
R12501 gnd.n4427 gnd.n4426 9.3005
R12502 gnd.n4425 gnd.n1398 9.3005
R12503 gnd.n4424 gnd.n4423 9.3005
R12504 gnd.n4422 gnd.n1399 9.3005
R12505 gnd.n4421 gnd.n4420 9.3005
R12506 gnd.n4419 gnd.n1403 9.3005
R12507 gnd.n4418 gnd.n4417 9.3005
R12508 gnd.n4416 gnd.n1404 9.3005
R12509 gnd.n4415 gnd.n4414 9.3005
R12510 gnd.n4413 gnd.n1408 9.3005
R12511 gnd.n4412 gnd.n4411 9.3005
R12512 gnd.n4410 gnd.n1409 9.3005
R12513 gnd.n4409 gnd.n4408 9.3005
R12514 gnd.n4407 gnd.n1413 9.3005
R12515 gnd.n4406 gnd.n4405 9.3005
R12516 gnd.n4404 gnd.n1414 9.3005
R12517 gnd.n4403 gnd.n4402 9.3005
R12518 gnd.n4401 gnd.n1418 9.3005
R12519 gnd.n4400 gnd.n4399 9.3005
R12520 gnd.n4398 gnd.n1419 9.3005
R12521 gnd.n4397 gnd.n4396 9.3005
R12522 gnd.n4395 gnd.n1423 9.3005
R12523 gnd.n4394 gnd.n4393 9.3005
R12524 gnd.n4392 gnd.n1424 9.3005
R12525 gnd.n4391 gnd.n4390 9.3005
R12526 gnd.n4389 gnd.n1428 9.3005
R12527 gnd.n4388 gnd.n4387 9.3005
R12528 gnd.n4386 gnd.n1429 9.3005
R12529 gnd.n4385 gnd.n4384 9.3005
R12530 gnd.n4383 gnd.n1433 9.3005
R12531 gnd.n4382 gnd.n4381 9.3005
R12532 gnd.n4380 gnd.n1434 9.3005
R12533 gnd.n4379 gnd.n1437 9.3005
R12534 gnd.n4502 gnd.n4501 9.3005
R12535 gnd.n1479 gnd.n1477 9.3005
R12536 gnd.n4353 gnd.n4352 9.3005
R12537 gnd.n4351 gnd.n1478 9.3005
R12538 gnd.n4350 gnd.n4349 9.3005
R12539 gnd.n4348 gnd.n1480 9.3005
R12540 gnd.n4347 gnd.n4346 9.3005
R12541 gnd.n4345 gnd.n1484 9.3005
R12542 gnd.n4344 gnd.n4343 9.3005
R12543 gnd.n4342 gnd.n1485 9.3005
R12544 gnd.n4341 gnd.n4340 9.3005
R12545 gnd.n4339 gnd.n1489 9.3005
R12546 gnd.n4338 gnd.n4337 9.3005
R12547 gnd.n4336 gnd.n1490 9.3005
R12548 gnd.n4335 gnd.n4334 9.3005
R12549 gnd.n4333 gnd.n1494 9.3005
R12550 gnd.n4332 gnd.n4331 9.3005
R12551 gnd.n241 gnd.n239 9.3005
R12552 gnd.n7111 gnd.n7110 9.3005
R12553 gnd.n7109 gnd.n240 9.3005
R12554 gnd.n7108 gnd.n7107 9.3005
R12555 gnd.n7106 gnd.n242 9.3005
R12556 gnd.n7105 gnd.n7104 9.3005
R12557 gnd.n7103 gnd.n246 9.3005
R12558 gnd.n7102 gnd.n7101 9.3005
R12559 gnd.n7100 gnd.n247 9.3005
R12560 gnd.n218 gnd.n217 9.3005
R12561 gnd.n7125 gnd.n7124 9.3005
R12562 gnd.n7126 gnd.n216 9.3005
R12563 gnd.n7128 gnd.n7127 9.3005
R12564 gnd.n201 gnd.n200 9.3005
R12565 gnd.n7141 gnd.n7140 9.3005
R12566 gnd.n7142 gnd.n199 9.3005
R12567 gnd.n7144 gnd.n7143 9.3005
R12568 gnd.n186 gnd.n185 9.3005
R12569 gnd.n7157 gnd.n7156 9.3005
R12570 gnd.n7158 gnd.n184 9.3005
R12571 gnd.n7160 gnd.n7159 9.3005
R12572 gnd.n167 gnd.n166 9.3005
R12573 gnd.n7175 gnd.n7174 9.3005
R12574 gnd.n7176 gnd.n164 9.3005
R12575 gnd.n7245 gnd.n7244 9.3005
R12576 gnd.n7243 gnd.n165 9.3005
R12577 gnd.n1646 gnd.n1645 9.3005
R12578 gnd.n7240 gnd.n7177 9.3005
R12579 gnd.n7239 gnd.n7238 9.3005
R12580 gnd.n7237 gnd.n7182 9.3005
R12581 gnd.n7236 gnd.n7235 9.3005
R12582 gnd.n7234 gnd.n7183 9.3005
R12583 gnd.n7233 gnd.n7232 9.3005
R12584 gnd.n7231 gnd.n7190 9.3005
R12585 gnd.n7230 gnd.n7229 9.3005
R12586 gnd.n7228 gnd.n7191 9.3005
R12587 gnd.n7227 gnd.n7226 9.3005
R12588 gnd.n7225 gnd.n7198 9.3005
R12589 gnd.n7224 gnd.n7223 9.3005
R12590 gnd.n7222 gnd.n7199 9.3005
R12591 gnd.n7221 gnd.n7220 9.3005
R12592 gnd.n7219 gnd.n7206 9.3005
R12593 gnd.n7218 gnd.n7217 9.3005
R12594 gnd.n7216 gnd.n7207 9.3005
R12595 gnd.n7215 gnd.n78 9.3005
R12596 gnd.n7242 gnd.n7241 9.3005
R12597 gnd.n4146 gnd.n4145 9.3005
R12598 gnd.n1592 gnd.n1591 9.3005
R12599 gnd.n4179 gnd.n4178 9.3005
R12600 gnd.n4180 gnd.n1589 9.3005
R12601 gnd.n4183 gnd.n4182 9.3005
R12602 gnd.n4181 gnd.n1590 9.3005
R12603 gnd.n1553 gnd.n1552 9.3005
R12604 gnd.n4210 gnd.n4209 9.3005
R12605 gnd.n4211 gnd.n1550 9.3005
R12606 gnd.n4220 gnd.n4219 9.3005
R12607 gnd.n4218 gnd.n1551 9.3005
R12608 gnd.n4217 gnd.n4216 9.3005
R12609 gnd.n4215 gnd.n4212 9.3005
R12610 gnd.n1507 gnd.n1505 9.3005
R12611 gnd.n4324 gnd.n4323 9.3005
R12612 gnd.n4322 gnd.n1506 9.3005
R12613 gnd.n4321 gnd.n4320 9.3005
R12614 gnd.n4319 gnd.n1508 9.3005
R12615 gnd.n4318 gnd.n4317 9.3005
R12616 gnd.n4316 gnd.n51 9.3005
R12617 gnd.n7360 gnd.n52 9.3005
R12618 gnd.n7359 gnd.n7358 9.3005
R12619 gnd.n7357 gnd.n53 9.3005
R12620 gnd.n7356 gnd.n7355 9.3005
R12621 gnd.n7354 gnd.n57 9.3005
R12622 gnd.n7353 gnd.n7352 9.3005
R12623 gnd.n7351 gnd.n58 9.3005
R12624 gnd.n7350 gnd.n7349 9.3005
R12625 gnd.n7348 gnd.n62 9.3005
R12626 gnd.n7347 gnd.n7346 9.3005
R12627 gnd.n7345 gnd.n63 9.3005
R12628 gnd.n7344 gnd.n7343 9.3005
R12629 gnd.n7342 gnd.n67 9.3005
R12630 gnd.n7341 gnd.n7340 9.3005
R12631 gnd.n7339 gnd.n68 9.3005
R12632 gnd.n7338 gnd.n7337 9.3005
R12633 gnd.n7336 gnd.n72 9.3005
R12634 gnd.n7335 gnd.n7334 9.3005
R12635 gnd.n7333 gnd.n73 9.3005
R12636 gnd.n7332 gnd.n7331 9.3005
R12637 gnd.n7330 gnd.n77 9.3005
R12638 gnd.n7329 gnd.n7328 9.3005
R12639 gnd.n4144 gnd.n1597 9.3005
R12640 gnd.t21 gnd.n4859 9.24152
R12641 gnd.n6063 gnd.t36 9.24152
R12642 gnd.t90 gnd.n1006 9.24152
R12643 gnd.n2929 gnd.t176 9.24152
R12644 gnd.t228 gnd.n4196 9.24152
R12645 gnd.t157 gnd.t21 8.92286
R12646 gnd.n3432 gnd.n3431 8.92286
R12647 gnd.n3536 gnd.n2177 8.92286
R12648 gnd.n3390 gnd.n2139 8.92286
R12649 gnd.t139 gnd.n3584 8.92286
R12650 gnd.n3665 gnd.t4 8.92286
R12651 gnd.n3645 gnd.n2084 8.92286
R12652 gnd.n3745 gnd.n2044 8.92286
R12653 gnd.n3862 gnd.n1983 8.92286
R12654 gnd.n3852 gnd.t101 8.92286
R12655 gnd.n5917 gnd.n5892 8.92171
R12656 gnd.n5885 gnd.n5860 8.92171
R12657 gnd.n5853 gnd.n5828 8.92171
R12658 gnd.n5822 gnd.n5797 8.92171
R12659 gnd.n5790 gnd.n5765 8.92171
R12660 gnd.n5758 gnd.n5733 8.92171
R12661 gnd.n5726 gnd.n5701 8.92171
R12662 gnd.n5695 gnd.n5670 8.92171
R12663 gnd.n3906 gnd.n3888 8.72777
R12664 gnd.n5491 gnd.t11 8.60421
R12665 gnd.n4923 gnd.n4911 8.43467
R12666 gnd.n38 gnd.n26 8.43467
R12667 gnd.n2851 gnd.n0 8.41456
R12668 gnd.n7361 gnd.n7360 8.41456
R12669 gnd.t104 gnd.n2263 8.28555
R12670 gnd.t127 gnd.n2235 8.28555
R12671 gnd.n2215 gnd.t22 8.28555
R12672 gnd.n3527 gnd.n2184 8.28555
R12673 gnd.n3566 gnd.t149 8.28555
R12674 gnd.n3593 gnd.n3592 8.28555
R12675 gnd.n3668 gnd.n3667 8.28555
R12676 gnd.n3705 gnd.t135 8.28555
R12677 gnd.n3726 gnd.n2038 8.28555
R12678 gnd.t26 gnd.n2015 8.28555
R12679 gnd.n5918 gnd.n5890 8.14595
R12680 gnd.n5886 gnd.n5858 8.14595
R12681 gnd.n5854 gnd.n5826 8.14595
R12682 gnd.n5823 gnd.n5795 8.14595
R12683 gnd.n5791 gnd.n5763 8.14595
R12684 gnd.n5759 gnd.n5731 8.14595
R12685 gnd.n5727 gnd.n5699 8.14595
R12686 gnd.n5696 gnd.n5668 8.14595
R12687 gnd.n5923 gnd.n5922 7.97301
R12688 gnd.t13 gnd.n5006 7.9669
R12689 gnd.n7216 gnd.n7215 7.75808
R12690 gnd.n1729 gnd.n1606 7.75808
R12691 gnd.n3080 gnd.n3071 7.75808
R12692 gnd.n2726 gnd.n2725 7.75808
R12693 gnd.n3440 gnd.t54 7.64824
R12694 gnd.n3471 gnd.n3470 7.64824
R12695 gnd.n3519 gnd.n2184 7.64824
R12696 gnd.n3592 gnd.n2135 7.64824
R12697 gnd.n3668 gnd.n2088 7.64824
R12698 gnd.n3753 gnd.n2038 7.64824
R12699 gnd.n3804 gnd.n2002 7.64824
R12700 gnd.n5400 gnd.t16 7.32958
R12701 gnd.n2285 gnd.n2284 7.30353
R12702 gnd.n3905 gnd.n3904 7.30353
R12703 gnd.n5360 gnd.n5079 7.01093
R12704 gnd.n5082 gnd.n5080 7.01093
R12705 gnd.n5370 gnd.n5369 7.01093
R12706 gnd.n5381 gnd.n5063 7.01093
R12707 gnd.n5380 gnd.n5066 7.01093
R12708 gnd.n5391 gnd.n5054 7.01093
R12709 gnd.n5057 gnd.n5055 7.01093
R12710 gnd.n5401 gnd.n5400 7.01093
R12711 gnd.n5411 gnd.n5035 7.01093
R12712 gnd.n5410 gnd.n5038 7.01093
R12713 gnd.n5419 gnd.n5029 7.01093
R12714 gnd.n5431 gnd.n5019 7.01093
R12715 gnd.n5441 gnd.n5004 7.01093
R12716 gnd.n5457 gnd.n5456 7.01093
R12717 gnd.n5006 gnd.n4943 7.01093
R12718 gnd.n5511 gnd.n4944 7.01093
R12719 gnd.n5505 gnd.n5504 7.01093
R12720 gnd.n4993 gnd.n4955 7.01093
R12721 gnd.n5497 gnd.n4966 7.01093
R12722 gnd.n4984 gnd.n4979 7.01093
R12723 gnd.n5491 gnd.n5490 7.01093
R12724 gnd.n5537 gnd.n4894 7.01093
R12725 gnd.n5536 gnd.n5535 7.01093
R12726 gnd.n5548 gnd.n5547 7.01093
R12727 gnd.n4887 gnd.n4879 7.01093
R12728 gnd.n5577 gnd.n4867 7.01093
R12729 gnd.n5576 gnd.n4870 7.01093
R12730 gnd.n5587 gnd.n4859 7.01093
R12731 gnd.n4860 gnd.n4848 7.01093
R12732 gnd.n5600 gnd.n4849 7.01093
R12733 gnd.n5633 gnd.n4841 7.01093
R12734 gnd.n5632 gnd.n931 7.01093
R12735 gnd.n6098 gnd.n6097 7.01093
R12736 gnd.n5623 gnd.n5622 7.01093
R12737 gnd.n6091 gnd.n952 7.01093
R12738 gnd.n6090 gnd.n955 7.01093
R12739 gnd.n5615 gnd.n964 7.01093
R12740 gnd.n6084 gnd.n6083 7.01093
R12741 gnd.n6077 gnd.n977 7.01093
R12742 gnd.n6076 gnd.n980 7.01093
R12743 gnd.n5955 gnd.n989 7.01093
R12744 gnd.n6070 gnd.n6069 7.01093
R12745 gnd.n5936 gnd.n992 7.01093
R12746 gnd.n6063 gnd.n1003 7.01093
R12747 gnd.n6062 gnd.n1006 7.01093
R12748 gnd.n5966 gnd.n1014 7.01093
R12749 gnd.n6056 gnd.n6055 7.01093
R12750 gnd.n3536 gnd.n3535 7.01093
R12751 gnd.n3390 gnd.n2149 7.01093
R12752 gnd.n3585 gnd.t139 7.01093
R12753 gnd.n3675 gnd.t4 7.01093
R12754 gnd.n3645 gnd.n2074 7.01093
R12755 gnd.n3734 gnd.n2044 7.01093
R12756 gnd.n3862 gnd.n3861 7.01093
R12757 gnd.n3884 gnd.t101 7.01093
R12758 gnd.n5038 gnd.t9 6.69227
R12759 gnd.n4870 gnd.t157 6.69227
R12760 gnd.n6105 gnd.n931 6.69227
R12761 gnd.t8 gnd.n5947 6.69227
R12762 gnd.n2235 gnd.t153 6.69227
R12763 gnd.n3805 gnd.t274 6.69227
R12764 gnd.n4041 gnd.n4040 6.5566
R12765 gnd.n2391 gnd.n2390 6.5566
R12766 gnd.n3293 gnd.n2326 6.5566
R12767 gnd.n3916 gnd.n3915 6.5566
R12768 gnd.n3422 gnd.n3421 6.37362
R12769 gnd.n3509 gnd.n3508 6.37362
R12770 gnd.t136 gnd.n2172 6.37362
R12771 gnd.n3625 gnd.n2118 6.37362
R12772 gnd.n3641 gnd.n2102 6.37362
R12773 gnd.t150 gnd.n3713 6.37362
R12774 gnd.n3784 gnd.n2021 6.37362
R12775 gnd.n3814 gnd.n2007 6.37362
R12776 gnd.n3221 gnd.n2510 6.20656
R12777 gnd.n7291 gnd.n7288 6.20656
R12778 gnd.n4679 gnd.n4678 6.20656
R12779 gnd.n4133 gnd.n4130 6.20656
R12780 gnd.t167 gnd.n5467 6.05496
R12781 gnd.n5468 gnd.t17 6.05496
R12782 gnd.t0 gnd.n4894 6.05496
R12783 gnd.n5642 gnd.t18 6.05496
R12784 gnd.n2754 gnd.t116 6.05496
R12785 gnd.t32 gnd.n162 6.05496
R12786 gnd.n5920 gnd.n5890 5.81868
R12787 gnd.n5888 gnd.n5858 5.81868
R12788 gnd.n5856 gnd.n5826 5.81868
R12789 gnd.n5825 gnd.n5795 5.81868
R12790 gnd.n5793 gnd.n5763 5.81868
R12791 gnd.n5761 gnd.n5731 5.81868
R12792 gnd.n5729 gnd.n5699 5.81868
R12793 gnd.n5698 gnd.n5668 5.81868
R12794 gnd.n2265 gnd.n2254 5.73631
R12795 gnd.n3440 gnd.n2249 5.73631
R12796 gnd.n3555 gnd.n2163 5.73631
R12797 gnd.n3567 gnd.n2153 5.73631
R12798 gnd.n3704 gnd.n2068 5.73631
R12799 gnd.n3685 gnd.n2061 5.73631
R12800 gnd.n3848 gnd.n3847 5.73631
R12801 gnd.n3852 gnd.n3850 5.73631
R12802 gnd.n4045 gnd.n1958 5.62001
R12803 gnd.n3288 gnd.n2395 5.62001
R12804 gnd.n3289 gnd.n3288 5.62001
R12805 gnd.n3911 gnd.n1958 5.62001
R12806 gnd.n5219 gnd.n5214 5.4308
R12807 gnd.n4819 gnd.n4817 5.4308
R12808 gnd.n5535 gnd.t15 5.41765
R12809 gnd.t19 gnd.n5558 5.41765
R12810 gnd.t165 gnd.n941 5.41765
R12811 gnd.t143 gnd.n3500 5.41765
R12812 gnd.t276 gnd.n2023 5.41765
R12813 gnd.n2236 gnd.t127 5.09899
R12814 gnd.n3489 gnd.n2215 5.09899
R12815 gnd.n3502 gnd.n3501 5.09899
R12816 gnd.n3403 gnd.t155 5.09899
R12817 gnd.n3543 gnd.t136 5.09899
R12818 gnd.n3375 gnd.n3374 5.09899
R12819 gnd.n3634 gnd.n3633 5.09899
R12820 gnd.n3716 gnd.t150 5.09899
R12821 gnd.t3 gnd.n2046 5.09899
R12822 gnd.n3765 gnd.n2035 5.09899
R12823 gnd.n3792 gnd.n2015 5.09899
R12824 gnd.n5918 gnd.n5917 5.04292
R12825 gnd.n5886 gnd.n5885 5.04292
R12826 gnd.n5854 gnd.n5853 5.04292
R12827 gnd.n5823 gnd.n5822 5.04292
R12828 gnd.n5791 gnd.n5790 5.04292
R12829 gnd.n5759 gnd.n5758 5.04292
R12830 gnd.n5727 gnd.n5726 5.04292
R12831 gnd.n5696 gnd.n5695 5.04292
R12832 gnd.n4935 gnd.n4934 4.82753
R12833 gnd.n50 gnd.n49 4.82753
R12834 gnd.n5498 gnd.t6 4.78034
R12835 gnd.n4849 gnd.t12 4.78034
R12836 gnd.t272 gnd.n3154 4.78034
R12837 gnd.n4079 gnd.t147 4.78034
R12838 gnd.n4940 gnd.n4937 4.74817
R12839 gnd.n4990 gnd.n4900 4.74817
R12840 gnd.n4977 gnd.n4899 4.74817
R12841 gnd.n4898 gnd.n4897 4.74817
R12842 gnd.n4986 gnd.n4937 4.74817
R12843 gnd.n4987 gnd.n4900 4.74817
R12844 gnd.n4989 gnd.n4899 4.74817
R12845 gnd.n4976 gnd.n4898 4.74817
R12846 gnd.n7117 gnd.n7116 4.74817
R12847 gnd.n4311 gnd.n229 4.74817
R12848 gnd.n1516 gnd.n228 4.74817
R12849 gnd.n253 gnd.n227 4.74817
R12850 gnd.n7096 gnd.n226 4.74817
R12851 gnd.n7117 gnd.n230 4.74817
R12852 gnd.n7115 gnd.n229 4.74817
R12853 gnd.n4312 gnd.n228 4.74817
R12854 gnd.n1515 gnd.n227 4.74817
R12855 gnd.n254 gnd.n226 4.74817
R12856 gnd.n2608 gnd.n2605 4.74817
R12857 gnd.n2884 gnd.n2604 4.74817
R12858 gnd.n2880 gnd.n2603 4.74817
R12859 gnd.n2627 gnd.n2602 4.74817
R12860 gnd.n2623 gnd.n2601 4.74817
R12861 gnd.n4238 gnd.n4237 4.74817
R12862 gnd.n4301 gnd.n1521 4.74817
R12863 gnd.n4306 gnd.n4303 4.74817
R12864 gnd.n4304 gnd.n259 4.74817
R12865 gnd.n7090 gnd.n7089 4.74817
R12866 gnd.n4239 gnd.n4238 4.74817
R12867 gnd.n4235 gnd.n1521 4.74817
R12868 gnd.n4303 gnd.n4302 4.74817
R12869 gnd.n4305 gnd.n4304 4.74817
R12870 gnd.n7091 gnd.n7090 4.74817
R12871 gnd.n4586 gnd.n4585 4.74817
R12872 gnd.n1222 gnd.n1202 4.74817
R12873 gnd.n4573 gnd.n4572 4.74817
R12874 gnd.n1239 gnd.n1223 4.74817
R12875 gnd.n4560 gnd.n4559 4.74817
R12876 gnd.n4587 gnd.n4586 4.74817
R12877 gnd.n4584 gnd.n1202 4.74817
R12878 gnd.n4574 gnd.n4573 4.74817
R12879 gnd.n4571 gnd.n1223 4.74817
R12880 gnd.n4561 gnd.n4560 4.74817
R12881 gnd.n2620 gnd.n2605 4.74817
R12882 gnd.n2621 gnd.n2604 4.74817
R12883 gnd.n2883 gnd.n2603 4.74817
R12884 gnd.n2879 gnd.n2602 4.74817
R12885 gnd.n2626 gnd.n2601 4.74817
R12886 gnd.n4923 gnd.n4922 4.7074
R12887 gnd.n38 gnd.n37 4.7074
R12888 gnd.n4935 gnd.n4923 4.65959
R12889 gnd.n50 gnd.n38 4.65959
R12890 gnd.n1957 gnd.n1878 4.6132
R12891 gnd.n3284 gnd.n3283 4.6132
R12892 gnd.n3358 gnd.n3357 4.46168
R12893 gnd.n3438 gnd.n2242 4.46168
R12894 gnd.n3432 gnd.t81 4.46168
R12895 gnd.n3545 gnd.n3543 4.46168
R12896 gnd.n3565 gnd.n3564 4.46168
R12897 gnd.n3693 gnd.n3692 4.46168
R12898 gnd.n3716 gnd.n3715 4.46168
R12899 gnd.n3979 gnd.n1965 4.46168
R12900 gnd.n3901 gnd.n3888 4.46111
R12901 gnd.n5903 gnd.n5899 4.38594
R12902 gnd.n5871 gnd.n5867 4.38594
R12903 gnd.n5839 gnd.n5835 4.38594
R12904 gnd.n5808 gnd.n5804 4.38594
R12905 gnd.n5776 gnd.n5772 4.38594
R12906 gnd.n5744 gnd.n5740 4.38594
R12907 gnd.n5712 gnd.n5708 4.38594
R12908 gnd.n5681 gnd.n5677 4.38594
R12909 gnd.n5914 gnd.n5892 4.26717
R12910 gnd.n5882 gnd.n5860 4.26717
R12911 gnd.n5850 gnd.n5828 4.26717
R12912 gnd.n5819 gnd.n5797 4.26717
R12913 gnd.n5787 gnd.n5765 4.26717
R12914 gnd.n5755 gnd.n5733 4.26717
R12915 gnd.n5723 gnd.n5701 4.26717
R12916 gnd.n5692 gnd.n5670 4.26717
R12917 gnd.n5442 gnd.t7 4.14303
R12918 gnd.t10 gnd.n955 4.14303
R12919 gnd.t64 gnd.n1319 4.14303
R12920 gnd.t46 gnd.n1471 4.14303
R12921 gnd.n5922 gnd.n5921 4.08274
R12922 gnd.n4040 gnd.n4039 4.05904
R12923 gnd.n2390 gnd.n2389 4.05904
R12924 gnd.n3296 gnd.n2326 4.05904
R12925 gnd.n3917 gnd.n3916 4.05904
R12926 gnd.n15 gnd.n7 3.99943
R12927 gnd.n3481 gnd.n3480 3.82437
R12928 gnd.t156 gnd.n3411 3.82437
R12929 gnd.n3618 gnd.n2124 3.82437
R12930 gnd.n3655 gnd.n2097 3.82437
R12931 gnd.t173 gnd.n2028 3.82437
R12932 gnd.n3825 gnd.n1999 3.82437
R12933 gnd.n3878 gnd.t40 3.82437
R12934 gnd.n5515 gnd.n4936 3.76259
R12935 gnd.n5922 gnd.n5794 3.70378
R12936 gnd.n15 gnd.n14 3.60163
R12937 gnd.n3348 gnd.n2289 3.50571
R12938 gnd.n4048 gnd.n1804 3.50571
R12939 gnd.n5913 gnd.n5894 3.49141
R12940 gnd.n5881 gnd.n5862 3.49141
R12941 gnd.n5849 gnd.n5830 3.49141
R12942 gnd.n5818 gnd.n5799 3.49141
R12943 gnd.n5786 gnd.n5767 3.49141
R12944 gnd.n5754 gnd.n5735 3.49141
R12945 gnd.n5722 gnd.n5703 3.49141
R12946 gnd.n5691 gnd.n5672 3.49141
R12947 gnd.n3183 gnd.t43 3.18706
R12948 gnd.n3460 gnd.n2234 3.18706
R12949 gnd.n3404 gnd.n3403 3.18706
R12950 gnd.t149 gnd.n3565 3.18706
R12951 gnd.n3586 gnd.n3585 3.18706
R12952 gnd.n3675 gnd.n3674 3.18706
R12953 gnd.n3692 gnd.t135 3.18706
R12954 gnd.n3744 gnd.n2046 3.18706
R12955 gnd.n3836 gnd.n3835 3.18706
R12956 gnd.t78 gnd.n1983 3.18706
R12957 gnd.n5021 gnd.t7 2.8684
R12958 gnd.n3367 gnd.t140 2.8684
R12959 gnd.n3884 gnd.t137 2.8684
R12960 gnd.n4924 gnd.t256 2.82907
R12961 gnd.n4924 gnd.t224 2.82907
R12962 gnd.n4926 gnd.t247 2.82907
R12963 gnd.n4926 gnd.t175 2.82907
R12964 gnd.n4928 gnd.t194 2.82907
R12965 gnd.n4928 gnd.t183 2.82907
R12966 gnd.n4930 gnd.t179 2.82907
R12967 gnd.n4930 gnd.t264 2.82907
R12968 gnd.n4932 gnd.t185 2.82907
R12969 gnd.n4932 gnd.t217 2.82907
R12970 gnd.n4901 gnd.t189 2.82907
R12971 gnd.n4901 gnd.t207 2.82907
R12972 gnd.n4903 gnd.t216 2.82907
R12973 gnd.n4903 gnd.t257 2.82907
R12974 gnd.n4905 gnd.t206 2.82907
R12975 gnd.n4905 gnd.t199 2.82907
R12976 gnd.n4907 gnd.t232 2.82907
R12977 gnd.n4907 gnd.t226 2.82907
R12978 gnd.n4909 gnd.t261 2.82907
R12979 gnd.n4909 gnd.t213 2.82907
R12980 gnd.n4912 gnd.t263 2.82907
R12981 gnd.n4912 gnd.t191 2.82907
R12982 gnd.n4914 gnd.t203 2.82907
R12983 gnd.n4914 gnd.t242 2.82907
R12984 gnd.n4916 gnd.t187 2.82907
R12985 gnd.n4916 gnd.t269 2.82907
R12986 gnd.n4918 gnd.t215 2.82907
R12987 gnd.n4918 gnd.t212 2.82907
R12988 gnd.n4920 gnd.t249 2.82907
R12989 gnd.n4920 gnd.t198 2.82907
R12990 gnd.n47 gnd.t193 2.82907
R12991 gnd.n47 gnd.t262 2.82907
R12992 gnd.n45 gnd.t244 2.82907
R12993 gnd.n45 gnd.t253 2.82907
R12994 gnd.n43 gnd.t255 2.82907
R12995 gnd.n43 gnd.t266 2.82907
R12996 gnd.n41 gnd.t250 2.82907
R12997 gnd.n41 gnd.t221 2.82907
R12998 gnd.n39 gnd.t201 2.82907
R12999 gnd.n39 gnd.t241 2.82907
R13000 gnd.n24 gnd.t233 2.82907
R13001 gnd.n24 gnd.t251 2.82907
R13002 gnd.n22 gnd.t248 2.82907
R13003 gnd.n22 gnd.t254 2.82907
R13004 gnd.n20 gnd.t219 2.82907
R13005 gnd.n20 gnd.t196 2.82907
R13006 gnd.n18 gnd.t181 2.82907
R13007 gnd.n18 gnd.t236 2.82907
R13008 gnd.n16 gnd.t227 2.82907
R13009 gnd.n16 gnd.t267 2.82907
R13010 gnd.n35 gnd.t218 2.82907
R13011 gnd.n35 gnd.t238 2.82907
R13012 gnd.n33 gnd.t231 2.82907
R13013 gnd.n33 gnd.t235 2.82907
R13014 gnd.n31 gnd.t205 2.82907
R13015 gnd.n31 gnd.t265 2.82907
R13016 gnd.n29 gnd.t260 2.82907
R13017 gnd.n29 gnd.t222 2.82907
R13018 gnd.n27 gnd.t214 2.82907
R13019 gnd.n27 gnd.t258 2.82907
R13020 gnd.n5910 gnd.n5909 2.71565
R13021 gnd.n5878 gnd.n5877 2.71565
R13022 gnd.n5846 gnd.n5845 2.71565
R13023 gnd.n5815 gnd.n5814 2.71565
R13024 gnd.n5783 gnd.n5782 2.71565
R13025 gnd.n5751 gnd.n5750 2.71565
R13026 gnd.n5719 gnd.n5718 2.71565
R13027 gnd.n5688 gnd.n5687 2.71565
R13028 gnd.t54 gnd.n3439 2.54975
R13029 gnd.t81 gnd.n2244 2.54975
R13030 gnd.n3458 gnd.n2236 2.54975
R13031 gnd.t22 gnd.n2205 2.54975
R13032 gnd.n3526 gnd.n2186 2.54975
R13033 gnd.n3584 gnd.n2133 2.54975
R13034 gnd.n3666 gnd.n3665 2.54975
R13035 gnd.n3725 gnd.n2058 2.54975
R13036 gnd.n3766 gnd.t26 2.54975
R13037 gnd.n3833 gnd.n1993 2.54975
R13038 gnd.t130 gnd.n3868 2.54975
R13039 gnd.n5515 gnd.n4937 2.27742
R13040 gnd.n5515 gnd.n4900 2.27742
R13041 gnd.n5515 gnd.n4899 2.27742
R13042 gnd.n5515 gnd.n4898 2.27742
R13043 gnd.n7118 gnd.n7117 2.27742
R13044 gnd.n7118 gnd.n229 2.27742
R13045 gnd.n7118 gnd.n228 2.27742
R13046 gnd.n7118 gnd.n227 2.27742
R13047 gnd.n7118 gnd.n226 2.27742
R13048 gnd.n4238 gnd.n225 2.27742
R13049 gnd.n1521 gnd.n225 2.27742
R13050 gnd.n4303 gnd.n225 2.27742
R13051 gnd.n4304 gnd.n225 2.27742
R13052 gnd.n7090 gnd.n225 2.27742
R13053 gnd.n4586 gnd.n1200 2.27742
R13054 gnd.n1202 gnd.n1200 2.27742
R13055 gnd.n4573 gnd.n1200 2.27742
R13056 gnd.n1223 gnd.n1200 2.27742
R13057 gnd.n4560 gnd.n1200 2.27742
R13058 gnd.n2899 gnd.n2605 2.27742
R13059 gnd.n2899 gnd.n2604 2.27742
R13060 gnd.n2899 gnd.n2603 2.27742
R13061 gnd.n2899 gnd.n2602 2.27742
R13062 gnd.n2899 gnd.n2601 2.27742
R13063 gnd.n5369 gnd.t50 2.23109
R13064 gnd.n4992 gnd.t6 2.23109
R13065 gnd.n3564 gnd.t159 2.23109
R13066 gnd.t161 gnd.n3693 2.23109
R13067 gnd.n5906 gnd.n5896 1.93989
R13068 gnd.n5874 gnd.n5864 1.93989
R13069 gnd.n5842 gnd.n5832 1.93989
R13070 gnd.n5811 gnd.n5801 1.93989
R13071 gnd.n5779 gnd.n5769 1.93989
R13072 gnd.n5747 gnd.n5737 1.93989
R13073 gnd.n5715 gnd.n5705 1.93989
R13074 gnd.n5684 gnd.n5674 1.93989
R13075 gnd.n2265 gnd.t104 1.91244
R13076 gnd.n3469 gnd.n3468 1.91244
R13077 gnd.n3520 gnd.n2191 1.91244
R13078 gnd.n3383 gnd.n3382 1.91244
R13079 gnd.n3618 gnd.t142 1.91244
R13080 gnd.t25 gnd.n2097 1.91244
R13081 gnd.n3654 gnd.n3653 1.91244
R13082 gnd.n3756 gnd.n3755 1.91244
R13083 gnd.n3824 gnd.n3823 1.91244
R13084 gnd.n3869 gnd.t130 1.91244
R13085 gnd.t169 gnd.n5380 1.59378
R13086 gnd.n5559 gnd.t19 1.59378
R13087 gnd.n4835 gnd.t165 1.59378
R13088 gnd.n3471 gnd.t153 1.59378
R13089 gnd.t151 gnd.n2177 1.59378
R13090 gnd.n3745 gnd.t280 1.59378
R13091 gnd.t274 gnd.n3804 1.59378
R13092 gnd.n3359 gnd.n2260 1.27512
R13093 gnd.t28 gnd.n3438 1.27512
R13094 gnd.n3450 gnd.n3449 1.27512
R13095 gnd.n3481 gnd.t2 1.27512
R13096 gnd.n3546 gnd.n2170 1.27512
R13097 gnd.n3574 gnd.n3573 1.27512
R13098 gnd.n3695 gnd.n3694 1.27512
R13099 gnd.n3735 gnd.n2051 1.27512
R13100 gnd.n3825 gnd.t5 1.27512
R13101 gnd.n3870 gnd.n1977 1.27512
R13102 gnd.n3868 gnd.t57 1.27512
R13103 gnd.n3878 gnd.n1786 1.27512
R13104 gnd.n1804 gnd.t113 1.27512
R13105 gnd.n5222 gnd.n5214 1.16414
R13106 gnd.n5981 gnd.n4817 1.16414
R13107 gnd.n5905 gnd.n5898 1.16414
R13108 gnd.n5873 gnd.n5866 1.16414
R13109 gnd.n5841 gnd.n5834 1.16414
R13110 gnd.n5810 gnd.n5803 1.16414
R13111 gnd.n5778 gnd.n5771 1.16414
R13112 gnd.n5746 gnd.n5739 1.16414
R13113 gnd.n5714 gnd.n5707 1.16414
R13114 gnd.n5683 gnd.n5676 1.16414
R13115 gnd.n1957 gnd.n1956 0.970197
R13116 gnd.n3284 gnd.n2396 0.970197
R13117 gnd.n5889 gnd.n5857 0.962709
R13118 gnd.n5921 gnd.n5889 0.962709
R13119 gnd.n5762 gnd.n5730 0.962709
R13120 gnd.n5794 gnd.n5762 0.962709
R13121 gnd.n5468 gnd.t167 0.956468
R13122 gnd.n6104 gnd.t18 0.956468
R13123 gnd.n2799 gnd.t208 0.956468
R13124 gnd.n4608 gnd.t184 0.956468
R13125 gnd.n2961 gnd.t188 0.956468
R13126 gnd.n2923 gnd.t190 0.956468
R13127 gnd.n3180 gnd.t270 0.956468
R13128 gnd.n4060 gnd.t171 0.956468
R13129 gnd.n4164 gnd.t200 0.956468
R13130 gnd.n4248 gnd.t240 0.956468
R13131 gnd.n7146 gnd.t237 0.956468
R13132 gnd.n7066 gnd.t245 0.956468
R13133 gnd.n4931 gnd.n4929 0.773756
R13134 gnd.n46 gnd.n44 0.773756
R13135 gnd.n4934 gnd.n4933 0.773756
R13136 gnd.n4933 gnd.n4931 0.773756
R13137 gnd.n4929 gnd.n4927 0.773756
R13138 gnd.n4927 gnd.n4925 0.773756
R13139 gnd.n42 gnd.n40 0.773756
R13140 gnd.n44 gnd.n42 0.773756
R13141 gnd.n48 gnd.n46 0.773756
R13142 gnd.n49 gnd.n48 0.773756
R13143 gnd.n2 gnd.n1 0.672012
R13144 gnd.n3 gnd.n2 0.672012
R13145 gnd.n4 gnd.n3 0.672012
R13146 gnd.n5 gnd.n4 0.672012
R13147 gnd.n6 gnd.n5 0.672012
R13148 gnd.n7 gnd.n6 0.672012
R13149 gnd.n9 gnd.n8 0.672012
R13150 gnd.n10 gnd.n9 0.672012
R13151 gnd.n11 gnd.n10 0.672012
R13152 gnd.n12 gnd.n11 0.672012
R13153 gnd.n13 gnd.n12 0.672012
R13154 gnd.n14 gnd.n13 0.672012
R13155 gnd.n3491 gnd.n2214 0.637812
R13156 gnd.n3500 gnd.n2199 0.637812
R13157 gnd.n3624 gnd.n2120 0.637812
R13158 gnd.n2112 gnd.n2111 0.637812
R13159 gnd.n3783 gnd.n2023 0.637812
R13160 gnd.n3795 gnd.n3794 0.637812
R13161 gnd.n4911 gnd.n4910 0.573776
R13162 gnd.n4910 gnd.n4908 0.573776
R13163 gnd.n4908 gnd.n4906 0.573776
R13164 gnd.n4906 gnd.n4904 0.573776
R13165 gnd.n4904 gnd.n4902 0.573776
R13166 gnd.n4922 gnd.n4921 0.573776
R13167 gnd.n4921 gnd.n4919 0.573776
R13168 gnd.n4919 gnd.n4917 0.573776
R13169 gnd.n4917 gnd.n4915 0.573776
R13170 gnd.n4915 gnd.n4913 0.573776
R13171 gnd.n19 gnd.n17 0.573776
R13172 gnd.n21 gnd.n19 0.573776
R13173 gnd.n23 gnd.n21 0.573776
R13174 gnd.n25 gnd.n23 0.573776
R13175 gnd.n26 gnd.n25 0.573776
R13176 gnd.n30 gnd.n28 0.573776
R13177 gnd.n32 gnd.n30 0.573776
R13178 gnd.n34 gnd.n32 0.573776
R13179 gnd.n36 gnd.n34 0.573776
R13180 gnd.n37 gnd.n36 0.573776
R13181 gnd gnd.n0 0.551497
R13182 gnd.n7118 gnd.n225 0.548625
R13183 gnd.n2899 gnd.n1200 0.548625
R13184 gnd.n2729 gnd.n2727 0.532512
R13185 gnd.n2685 gnd.n1124 0.532512
R13186 gnd.n7243 gnd.n7242 0.532512
R13187 gnd.n7329 gnd.n78 0.532512
R13188 gnd.n4503 gnd.n4502 0.523366
R13189 gnd.n1644 gnd.n1437 0.523366
R13190 gnd.n7323 gnd.n7322 0.520317
R13191 gnd.n7252 gnd.n7251 0.520317
R13192 gnd.n1915 gnd.n1595 0.520317
R13193 gnd.n1839 gnd.n1466 0.520317
R13194 gnd.n2417 gnd.n1324 0.520317
R13195 gnd.n3244 gnd.n3243 0.520317
R13196 gnd.n4639 gnd.n1116 0.520317
R13197 gnd.n2662 gnd.n1073 0.520317
R13198 gnd.n4120 gnd.n4119 0.489829
R13199 gnd.n3217 gnd.n3216 0.489829
R13200 gnd.n5971 gnd.n5970 0.486781
R13201 gnd.n5271 gnd.n5270 0.48678
R13202 gnd.n6052 gnd.n6051 0.480683
R13203 gnd.n5355 gnd.n5354 0.480683
R13204 gnd.n7362 gnd.n7361 0.470187
R13205 gnd.n6277 gnd.n761 0.468488
R13206 gnd.n6798 gnd.n450 0.468488
R13207 gnd.n7009 gnd.n7008 0.468488
R13208 gnd.n1020 gnd.n1019 0.468488
R13209 gnd.n4505 gnd.n4504 0.432431
R13210 gnd.n1647 gnd.n1646 0.432431
R13211 gnd.n3224 gnd.n2510 0.388379
R13212 gnd.n5902 gnd.n5901 0.388379
R13213 gnd.n5870 gnd.n5869 0.388379
R13214 gnd.n5838 gnd.n5837 0.388379
R13215 gnd.n5807 gnd.n5806 0.388379
R13216 gnd.n5775 gnd.n5774 0.388379
R13217 gnd.n5743 gnd.n5742 0.388379
R13218 gnd.n5711 gnd.n5710 0.388379
R13219 gnd.n5680 gnd.n5679 0.388379
R13220 gnd.n7292 gnd.n7291 0.388379
R13221 gnd.n4680 gnd.n4679 0.388379
R13222 gnd.n4134 gnd.n4133 0.388379
R13223 gnd.n7362 gnd.n15 0.374463
R13224 gnd.n5948 gnd.t8 0.319156
R13225 gnd.n2836 gnd.t178 0.319156
R13226 gnd.n2893 gnd.t211 0.319156
R13227 gnd.n2877 gnd.t182 0.319156
R13228 gnd.n2868 gnd.t202 0.319156
R13229 gnd.n3142 gnd.t97 0.319156
R13230 gnd.t142 gnd.t282 0.319156
R13231 gnd.t278 gnd.t25 0.319156
R13232 gnd.n4114 gnd.t74 0.319156
R13233 gnd.n4268 gnd.t220 0.319156
R13234 gnd.n4299 gnd.t204 0.319156
R13235 gnd.n7098 gnd.t230 0.319156
R13236 gnd.n7085 gnd.t234 0.319156
R13237 gnd.n5189 gnd.n5167 0.311721
R13238 gnd.n3235 gnd.n3234 0.302329
R13239 gnd.n4144 gnd.n4143 0.302329
R13240 gnd gnd.n7362 0.295112
R13241 gnd.n6021 gnd.n6020 0.268793
R13242 gnd.n6020 gnd.n6019 0.241354
R13243 gnd.n1878 gnd.n1877 0.229039
R13244 gnd.n1881 gnd.n1878 0.229039
R13245 gnd.n3283 gnd.n2401 0.229039
R13246 gnd.n3283 gnd.n3282 0.229039
R13247 gnd.n5343 gnd.n5142 0.206293
R13248 gnd.n5919 gnd.n5891 0.155672
R13249 gnd.n5912 gnd.n5891 0.155672
R13250 gnd.n5912 gnd.n5911 0.155672
R13251 gnd.n5911 gnd.n5895 0.155672
R13252 gnd.n5904 gnd.n5895 0.155672
R13253 gnd.n5904 gnd.n5903 0.155672
R13254 gnd.n5887 gnd.n5859 0.155672
R13255 gnd.n5880 gnd.n5859 0.155672
R13256 gnd.n5880 gnd.n5879 0.155672
R13257 gnd.n5879 gnd.n5863 0.155672
R13258 gnd.n5872 gnd.n5863 0.155672
R13259 gnd.n5872 gnd.n5871 0.155672
R13260 gnd.n5855 gnd.n5827 0.155672
R13261 gnd.n5848 gnd.n5827 0.155672
R13262 gnd.n5848 gnd.n5847 0.155672
R13263 gnd.n5847 gnd.n5831 0.155672
R13264 gnd.n5840 gnd.n5831 0.155672
R13265 gnd.n5840 gnd.n5839 0.155672
R13266 gnd.n5824 gnd.n5796 0.155672
R13267 gnd.n5817 gnd.n5796 0.155672
R13268 gnd.n5817 gnd.n5816 0.155672
R13269 gnd.n5816 gnd.n5800 0.155672
R13270 gnd.n5809 gnd.n5800 0.155672
R13271 gnd.n5809 gnd.n5808 0.155672
R13272 gnd.n5792 gnd.n5764 0.155672
R13273 gnd.n5785 gnd.n5764 0.155672
R13274 gnd.n5785 gnd.n5784 0.155672
R13275 gnd.n5784 gnd.n5768 0.155672
R13276 gnd.n5777 gnd.n5768 0.155672
R13277 gnd.n5777 gnd.n5776 0.155672
R13278 gnd.n5760 gnd.n5732 0.155672
R13279 gnd.n5753 gnd.n5732 0.155672
R13280 gnd.n5753 gnd.n5752 0.155672
R13281 gnd.n5752 gnd.n5736 0.155672
R13282 gnd.n5745 gnd.n5736 0.155672
R13283 gnd.n5745 gnd.n5744 0.155672
R13284 gnd.n5728 gnd.n5700 0.155672
R13285 gnd.n5721 gnd.n5700 0.155672
R13286 gnd.n5721 gnd.n5720 0.155672
R13287 gnd.n5720 gnd.n5704 0.155672
R13288 gnd.n5713 gnd.n5704 0.155672
R13289 gnd.n5713 gnd.n5712 0.155672
R13290 gnd.n5697 gnd.n5669 0.155672
R13291 gnd.n5690 gnd.n5669 0.155672
R13292 gnd.n5690 gnd.n5689 0.155672
R13293 gnd.n5689 gnd.n5673 0.155672
R13294 gnd.n5682 gnd.n5673 0.155672
R13295 gnd.n5682 gnd.n5681 0.155672
R13296 gnd.n6051 gnd.n4747 0.152939
R13297 gnd.n4749 gnd.n4747 0.152939
R13298 gnd.n4753 gnd.n4749 0.152939
R13299 gnd.n4754 gnd.n4753 0.152939
R13300 gnd.n4755 gnd.n4754 0.152939
R13301 gnd.n4756 gnd.n4755 0.152939
R13302 gnd.n4760 gnd.n4756 0.152939
R13303 gnd.n4761 gnd.n4760 0.152939
R13304 gnd.n4762 gnd.n4761 0.152939
R13305 gnd.n4763 gnd.n4762 0.152939
R13306 gnd.n4767 gnd.n4763 0.152939
R13307 gnd.n4768 gnd.n4767 0.152939
R13308 gnd.n4769 gnd.n4768 0.152939
R13309 gnd.n4770 gnd.n4769 0.152939
R13310 gnd.n4775 gnd.n4770 0.152939
R13311 gnd.n6021 gnd.n4775 0.152939
R13312 gnd.n5356 gnd.n5355 0.152939
R13313 gnd.n5356 gnd.n5060 0.152939
R13314 gnd.n5384 gnd.n5060 0.152939
R13315 gnd.n5385 gnd.n5384 0.152939
R13316 gnd.n5386 gnd.n5385 0.152939
R13317 gnd.n5387 gnd.n5386 0.152939
R13318 gnd.n5387 gnd.n5032 0.152939
R13319 gnd.n5414 gnd.n5032 0.152939
R13320 gnd.n5415 gnd.n5414 0.152939
R13321 gnd.n5416 gnd.n5415 0.152939
R13322 gnd.n5416 gnd.n5010 0.152939
R13323 gnd.n5445 gnd.n5010 0.152939
R13324 gnd.n5446 gnd.n5445 0.152939
R13325 gnd.n5447 gnd.n5446 0.152939
R13326 gnd.n5448 gnd.n5447 0.152939
R13327 gnd.n5450 gnd.n5448 0.152939
R13328 gnd.n5450 gnd.n5449 0.152939
R13329 gnd.n5449 gnd.n4959 0.152939
R13330 gnd.n4960 gnd.n4959 0.152939
R13331 gnd.n4961 gnd.n4960 0.152939
R13332 gnd.n4980 gnd.n4961 0.152939
R13333 gnd.n4981 gnd.n4980 0.152939
R13334 gnd.n4981 gnd.n4891 0.152939
R13335 gnd.n5540 gnd.n4891 0.152939
R13336 gnd.n5541 gnd.n5540 0.152939
R13337 gnd.n5542 gnd.n5541 0.152939
R13338 gnd.n5543 gnd.n5542 0.152939
R13339 gnd.n5543 gnd.n4864 0.152939
R13340 gnd.n5580 gnd.n4864 0.152939
R13341 gnd.n5581 gnd.n5580 0.152939
R13342 gnd.n5582 gnd.n5581 0.152939
R13343 gnd.n5583 gnd.n5582 0.152939
R13344 gnd.n5583 gnd.n4838 0.152939
R13345 gnd.n5636 gnd.n4838 0.152939
R13346 gnd.n5637 gnd.n5636 0.152939
R13347 gnd.n5639 gnd.n5637 0.152939
R13348 gnd.n5639 gnd.n5638 0.152939
R13349 gnd.n5638 gnd.n947 0.152939
R13350 gnd.n948 gnd.n947 0.152939
R13351 gnd.n949 gnd.n948 0.152939
R13352 gnd.n970 gnd.n949 0.152939
R13353 gnd.n971 gnd.n970 0.152939
R13354 gnd.n972 gnd.n971 0.152939
R13355 gnd.n973 gnd.n972 0.152939
R13356 gnd.n974 gnd.n973 0.152939
R13357 gnd.n996 gnd.n974 0.152939
R13358 gnd.n997 gnd.n996 0.152939
R13359 gnd.n998 gnd.n997 0.152939
R13360 gnd.n999 gnd.n998 0.152939
R13361 gnd.n1000 gnd.n999 0.152939
R13362 gnd.n4745 gnd.n1000 0.152939
R13363 gnd.n4746 gnd.n4745 0.152939
R13364 gnd.n6052 gnd.n4746 0.152939
R13365 gnd.n5354 gnd.n5084 0.152939
R13366 gnd.n5105 gnd.n5084 0.152939
R13367 gnd.n5106 gnd.n5105 0.152939
R13368 gnd.n5112 gnd.n5106 0.152939
R13369 gnd.n5113 gnd.n5112 0.152939
R13370 gnd.n5114 gnd.n5113 0.152939
R13371 gnd.n5114 gnd.n5103 0.152939
R13372 gnd.n5122 gnd.n5103 0.152939
R13373 gnd.n5123 gnd.n5122 0.152939
R13374 gnd.n5124 gnd.n5123 0.152939
R13375 gnd.n5124 gnd.n5101 0.152939
R13376 gnd.n5132 gnd.n5101 0.152939
R13377 gnd.n5133 gnd.n5132 0.152939
R13378 gnd.n5134 gnd.n5133 0.152939
R13379 gnd.n5134 gnd.n5099 0.152939
R13380 gnd.n5142 gnd.n5099 0.152939
R13381 gnd.n6019 gnd.n4777 0.152939
R13382 gnd.n4779 gnd.n4777 0.152939
R13383 gnd.n4783 gnd.n4779 0.152939
R13384 gnd.n4784 gnd.n4783 0.152939
R13385 gnd.n4785 gnd.n4784 0.152939
R13386 gnd.n4786 gnd.n4785 0.152939
R13387 gnd.n4790 gnd.n4786 0.152939
R13388 gnd.n4791 gnd.n4790 0.152939
R13389 gnd.n4792 gnd.n4791 0.152939
R13390 gnd.n4793 gnd.n4792 0.152939
R13391 gnd.n4797 gnd.n4793 0.152939
R13392 gnd.n4798 gnd.n4797 0.152939
R13393 gnd.n4799 gnd.n4798 0.152939
R13394 gnd.n4800 gnd.n4799 0.152939
R13395 gnd.n4804 gnd.n4800 0.152939
R13396 gnd.n4805 gnd.n4804 0.152939
R13397 gnd.n4806 gnd.n4805 0.152939
R13398 gnd.n4807 gnd.n4806 0.152939
R13399 gnd.n4811 gnd.n4807 0.152939
R13400 gnd.n4812 gnd.n4811 0.152939
R13401 gnd.n4813 gnd.n4812 0.152939
R13402 gnd.n4814 gnd.n4813 0.152939
R13403 gnd.n4821 gnd.n4814 0.152939
R13404 gnd.n4822 gnd.n4821 0.152939
R13405 gnd.n4823 gnd.n4822 0.152939
R13406 gnd.n5971 gnd.n4823 0.152939
R13407 gnd.n5517 gnd.n5516 0.152939
R13408 gnd.n5518 gnd.n5517 0.152939
R13409 gnd.n5519 gnd.n5518 0.152939
R13410 gnd.n5520 gnd.n5519 0.152939
R13411 gnd.n5521 gnd.n5520 0.152939
R13412 gnd.n5522 gnd.n5521 0.152939
R13413 gnd.n5522 gnd.n4845 0.152939
R13414 gnd.n5603 gnd.n4845 0.152939
R13415 gnd.n5604 gnd.n5603 0.152939
R13416 gnd.n5605 gnd.n5604 0.152939
R13417 gnd.n5606 gnd.n5605 0.152939
R13418 gnd.n5607 gnd.n5606 0.152939
R13419 gnd.n5608 gnd.n5607 0.152939
R13420 gnd.n5609 gnd.n5608 0.152939
R13421 gnd.n5610 gnd.n5609 0.152939
R13422 gnd.n5611 gnd.n5610 0.152939
R13423 gnd.n5612 gnd.n5611 0.152939
R13424 gnd.n5613 gnd.n5612 0.152939
R13425 gnd.n5613 gnd.n4828 0.152939
R13426 gnd.n5952 gnd.n4828 0.152939
R13427 gnd.n5953 gnd.n5952 0.152939
R13428 gnd.n5954 gnd.n5953 0.152939
R13429 gnd.n5954 gnd.n4826 0.152939
R13430 gnd.n5962 gnd.n4826 0.152939
R13431 gnd.n5963 gnd.n5962 0.152939
R13432 gnd.n5964 gnd.n5963 0.152939
R13433 gnd.n5964 gnd.n4824 0.152939
R13434 gnd.n5970 gnd.n4824 0.152939
R13435 gnd.n5272 gnd.n5271 0.152939
R13436 gnd.n5272 gnd.n5162 0.152939
R13437 gnd.n5287 gnd.n5162 0.152939
R13438 gnd.n5288 gnd.n5287 0.152939
R13439 gnd.n5289 gnd.n5288 0.152939
R13440 gnd.n5289 gnd.n5150 0.152939
R13441 gnd.n5303 gnd.n5150 0.152939
R13442 gnd.n5304 gnd.n5303 0.152939
R13443 gnd.n5305 gnd.n5304 0.152939
R13444 gnd.n5306 gnd.n5305 0.152939
R13445 gnd.n5307 gnd.n5306 0.152939
R13446 gnd.n5308 gnd.n5307 0.152939
R13447 gnd.n5309 gnd.n5308 0.152939
R13448 gnd.n5310 gnd.n5309 0.152939
R13449 gnd.n5311 gnd.n5310 0.152939
R13450 gnd.n5312 gnd.n5311 0.152939
R13451 gnd.n5313 gnd.n5312 0.152939
R13452 gnd.n5314 gnd.n5313 0.152939
R13453 gnd.n5315 gnd.n5314 0.152939
R13454 gnd.n5316 gnd.n5315 0.152939
R13455 gnd.n5317 gnd.n5316 0.152939
R13456 gnd.n5317 gnd.n5016 0.152939
R13457 gnd.n5434 gnd.n5016 0.152939
R13458 gnd.n5435 gnd.n5434 0.152939
R13459 gnd.n5436 gnd.n5435 0.152939
R13460 gnd.n5437 gnd.n5436 0.152939
R13461 gnd.n5437 gnd.n4938 0.152939
R13462 gnd.n5514 gnd.n4938 0.152939
R13463 gnd.n5190 gnd.n5189 0.152939
R13464 gnd.n5191 gnd.n5190 0.152939
R13465 gnd.n5192 gnd.n5191 0.152939
R13466 gnd.n5193 gnd.n5192 0.152939
R13467 gnd.n5194 gnd.n5193 0.152939
R13468 gnd.n5195 gnd.n5194 0.152939
R13469 gnd.n5196 gnd.n5195 0.152939
R13470 gnd.n5197 gnd.n5196 0.152939
R13471 gnd.n5198 gnd.n5197 0.152939
R13472 gnd.n5199 gnd.n5198 0.152939
R13473 gnd.n5200 gnd.n5199 0.152939
R13474 gnd.n5201 gnd.n5200 0.152939
R13475 gnd.n5202 gnd.n5201 0.152939
R13476 gnd.n5203 gnd.n5202 0.152939
R13477 gnd.n5204 gnd.n5203 0.152939
R13478 gnd.n5205 gnd.n5204 0.152939
R13479 gnd.n5206 gnd.n5205 0.152939
R13480 gnd.n5207 gnd.n5206 0.152939
R13481 gnd.n5208 gnd.n5207 0.152939
R13482 gnd.n5209 gnd.n5208 0.152939
R13483 gnd.n5210 gnd.n5209 0.152939
R13484 gnd.n5211 gnd.n5210 0.152939
R13485 gnd.n5215 gnd.n5211 0.152939
R13486 gnd.n5216 gnd.n5215 0.152939
R13487 gnd.n5216 gnd.n5173 0.152939
R13488 gnd.n5270 gnd.n5173 0.152939
R13489 gnd.n6278 gnd.n6277 0.152939
R13490 gnd.n6279 gnd.n6278 0.152939
R13491 gnd.n6279 gnd.n755 0.152939
R13492 gnd.n6287 gnd.n755 0.152939
R13493 gnd.n6288 gnd.n6287 0.152939
R13494 gnd.n6289 gnd.n6288 0.152939
R13495 gnd.n6289 gnd.n749 0.152939
R13496 gnd.n6297 gnd.n749 0.152939
R13497 gnd.n6298 gnd.n6297 0.152939
R13498 gnd.n6299 gnd.n6298 0.152939
R13499 gnd.n6299 gnd.n743 0.152939
R13500 gnd.n6307 gnd.n743 0.152939
R13501 gnd.n6308 gnd.n6307 0.152939
R13502 gnd.n6309 gnd.n6308 0.152939
R13503 gnd.n6309 gnd.n737 0.152939
R13504 gnd.n6317 gnd.n737 0.152939
R13505 gnd.n6318 gnd.n6317 0.152939
R13506 gnd.n6319 gnd.n6318 0.152939
R13507 gnd.n6319 gnd.n731 0.152939
R13508 gnd.n6327 gnd.n731 0.152939
R13509 gnd.n6328 gnd.n6327 0.152939
R13510 gnd.n6329 gnd.n6328 0.152939
R13511 gnd.n6329 gnd.n725 0.152939
R13512 gnd.n6337 gnd.n725 0.152939
R13513 gnd.n6338 gnd.n6337 0.152939
R13514 gnd.n6339 gnd.n6338 0.152939
R13515 gnd.n6339 gnd.n719 0.152939
R13516 gnd.n6347 gnd.n719 0.152939
R13517 gnd.n6348 gnd.n6347 0.152939
R13518 gnd.n6349 gnd.n6348 0.152939
R13519 gnd.n6349 gnd.n713 0.152939
R13520 gnd.n6357 gnd.n713 0.152939
R13521 gnd.n6358 gnd.n6357 0.152939
R13522 gnd.n6359 gnd.n6358 0.152939
R13523 gnd.n6359 gnd.n707 0.152939
R13524 gnd.n6367 gnd.n707 0.152939
R13525 gnd.n6368 gnd.n6367 0.152939
R13526 gnd.n6369 gnd.n6368 0.152939
R13527 gnd.n6369 gnd.n701 0.152939
R13528 gnd.n6377 gnd.n701 0.152939
R13529 gnd.n6378 gnd.n6377 0.152939
R13530 gnd.n6379 gnd.n6378 0.152939
R13531 gnd.n6379 gnd.n695 0.152939
R13532 gnd.n6387 gnd.n695 0.152939
R13533 gnd.n6388 gnd.n6387 0.152939
R13534 gnd.n6389 gnd.n6388 0.152939
R13535 gnd.n6389 gnd.n689 0.152939
R13536 gnd.n6397 gnd.n689 0.152939
R13537 gnd.n6398 gnd.n6397 0.152939
R13538 gnd.n6399 gnd.n6398 0.152939
R13539 gnd.n6399 gnd.n683 0.152939
R13540 gnd.n6407 gnd.n683 0.152939
R13541 gnd.n6408 gnd.n6407 0.152939
R13542 gnd.n6409 gnd.n6408 0.152939
R13543 gnd.n6409 gnd.n677 0.152939
R13544 gnd.n6417 gnd.n677 0.152939
R13545 gnd.n6418 gnd.n6417 0.152939
R13546 gnd.n6419 gnd.n6418 0.152939
R13547 gnd.n6419 gnd.n671 0.152939
R13548 gnd.n6427 gnd.n671 0.152939
R13549 gnd.n6428 gnd.n6427 0.152939
R13550 gnd.n6429 gnd.n6428 0.152939
R13551 gnd.n6429 gnd.n665 0.152939
R13552 gnd.n6437 gnd.n665 0.152939
R13553 gnd.n6438 gnd.n6437 0.152939
R13554 gnd.n6439 gnd.n6438 0.152939
R13555 gnd.n6439 gnd.n659 0.152939
R13556 gnd.n6447 gnd.n659 0.152939
R13557 gnd.n6448 gnd.n6447 0.152939
R13558 gnd.n6449 gnd.n6448 0.152939
R13559 gnd.n6449 gnd.n653 0.152939
R13560 gnd.n6457 gnd.n653 0.152939
R13561 gnd.n6458 gnd.n6457 0.152939
R13562 gnd.n6459 gnd.n6458 0.152939
R13563 gnd.n6459 gnd.n647 0.152939
R13564 gnd.n6467 gnd.n647 0.152939
R13565 gnd.n6468 gnd.n6467 0.152939
R13566 gnd.n6469 gnd.n6468 0.152939
R13567 gnd.n6469 gnd.n641 0.152939
R13568 gnd.n6477 gnd.n641 0.152939
R13569 gnd.n6478 gnd.n6477 0.152939
R13570 gnd.n6479 gnd.n6478 0.152939
R13571 gnd.n6479 gnd.n635 0.152939
R13572 gnd.n6487 gnd.n635 0.152939
R13573 gnd.n6488 gnd.n6487 0.152939
R13574 gnd.n6489 gnd.n6488 0.152939
R13575 gnd.n6489 gnd.n629 0.152939
R13576 gnd.n6497 gnd.n629 0.152939
R13577 gnd.n6498 gnd.n6497 0.152939
R13578 gnd.n6499 gnd.n6498 0.152939
R13579 gnd.n6499 gnd.n623 0.152939
R13580 gnd.n6507 gnd.n623 0.152939
R13581 gnd.n6508 gnd.n6507 0.152939
R13582 gnd.n6509 gnd.n6508 0.152939
R13583 gnd.n6509 gnd.n617 0.152939
R13584 gnd.n6517 gnd.n617 0.152939
R13585 gnd.n6518 gnd.n6517 0.152939
R13586 gnd.n6519 gnd.n6518 0.152939
R13587 gnd.n6519 gnd.n611 0.152939
R13588 gnd.n6527 gnd.n611 0.152939
R13589 gnd.n6528 gnd.n6527 0.152939
R13590 gnd.n6529 gnd.n6528 0.152939
R13591 gnd.n6529 gnd.n605 0.152939
R13592 gnd.n6537 gnd.n605 0.152939
R13593 gnd.n6538 gnd.n6537 0.152939
R13594 gnd.n6539 gnd.n6538 0.152939
R13595 gnd.n6539 gnd.n599 0.152939
R13596 gnd.n6547 gnd.n599 0.152939
R13597 gnd.n6548 gnd.n6547 0.152939
R13598 gnd.n6549 gnd.n6548 0.152939
R13599 gnd.n6549 gnd.n593 0.152939
R13600 gnd.n6557 gnd.n593 0.152939
R13601 gnd.n6558 gnd.n6557 0.152939
R13602 gnd.n6559 gnd.n6558 0.152939
R13603 gnd.n6559 gnd.n587 0.152939
R13604 gnd.n6567 gnd.n587 0.152939
R13605 gnd.n6568 gnd.n6567 0.152939
R13606 gnd.n6569 gnd.n6568 0.152939
R13607 gnd.n6569 gnd.n581 0.152939
R13608 gnd.n6577 gnd.n581 0.152939
R13609 gnd.n6578 gnd.n6577 0.152939
R13610 gnd.n6579 gnd.n6578 0.152939
R13611 gnd.n6579 gnd.n575 0.152939
R13612 gnd.n6587 gnd.n575 0.152939
R13613 gnd.n6588 gnd.n6587 0.152939
R13614 gnd.n6589 gnd.n6588 0.152939
R13615 gnd.n6589 gnd.n569 0.152939
R13616 gnd.n6597 gnd.n569 0.152939
R13617 gnd.n6598 gnd.n6597 0.152939
R13618 gnd.n6599 gnd.n6598 0.152939
R13619 gnd.n6599 gnd.n563 0.152939
R13620 gnd.n6607 gnd.n563 0.152939
R13621 gnd.n6608 gnd.n6607 0.152939
R13622 gnd.n6609 gnd.n6608 0.152939
R13623 gnd.n6609 gnd.n557 0.152939
R13624 gnd.n6617 gnd.n557 0.152939
R13625 gnd.n6618 gnd.n6617 0.152939
R13626 gnd.n6619 gnd.n6618 0.152939
R13627 gnd.n6619 gnd.n551 0.152939
R13628 gnd.n6627 gnd.n551 0.152939
R13629 gnd.n6628 gnd.n6627 0.152939
R13630 gnd.n6629 gnd.n6628 0.152939
R13631 gnd.n6629 gnd.n545 0.152939
R13632 gnd.n6637 gnd.n545 0.152939
R13633 gnd.n6638 gnd.n6637 0.152939
R13634 gnd.n6639 gnd.n6638 0.152939
R13635 gnd.n6639 gnd.n539 0.152939
R13636 gnd.n6647 gnd.n539 0.152939
R13637 gnd.n6648 gnd.n6647 0.152939
R13638 gnd.n6649 gnd.n6648 0.152939
R13639 gnd.n6649 gnd.n533 0.152939
R13640 gnd.n6657 gnd.n533 0.152939
R13641 gnd.n6658 gnd.n6657 0.152939
R13642 gnd.n6659 gnd.n6658 0.152939
R13643 gnd.n6659 gnd.n527 0.152939
R13644 gnd.n6667 gnd.n527 0.152939
R13645 gnd.n6668 gnd.n6667 0.152939
R13646 gnd.n6669 gnd.n6668 0.152939
R13647 gnd.n6669 gnd.n521 0.152939
R13648 gnd.n6677 gnd.n521 0.152939
R13649 gnd.n6678 gnd.n6677 0.152939
R13650 gnd.n6679 gnd.n6678 0.152939
R13651 gnd.n6679 gnd.n515 0.152939
R13652 gnd.n6687 gnd.n515 0.152939
R13653 gnd.n6688 gnd.n6687 0.152939
R13654 gnd.n6689 gnd.n6688 0.152939
R13655 gnd.n6689 gnd.n509 0.152939
R13656 gnd.n6697 gnd.n509 0.152939
R13657 gnd.n6698 gnd.n6697 0.152939
R13658 gnd.n6699 gnd.n6698 0.152939
R13659 gnd.n6699 gnd.n503 0.152939
R13660 gnd.n6707 gnd.n503 0.152939
R13661 gnd.n6708 gnd.n6707 0.152939
R13662 gnd.n6709 gnd.n6708 0.152939
R13663 gnd.n6709 gnd.n497 0.152939
R13664 gnd.n6717 gnd.n497 0.152939
R13665 gnd.n6718 gnd.n6717 0.152939
R13666 gnd.n6719 gnd.n6718 0.152939
R13667 gnd.n6719 gnd.n491 0.152939
R13668 gnd.n6727 gnd.n491 0.152939
R13669 gnd.n6728 gnd.n6727 0.152939
R13670 gnd.n6729 gnd.n6728 0.152939
R13671 gnd.n6729 gnd.n485 0.152939
R13672 gnd.n6737 gnd.n485 0.152939
R13673 gnd.n6738 gnd.n6737 0.152939
R13674 gnd.n6739 gnd.n6738 0.152939
R13675 gnd.n6739 gnd.n479 0.152939
R13676 gnd.n6747 gnd.n479 0.152939
R13677 gnd.n6748 gnd.n6747 0.152939
R13678 gnd.n6749 gnd.n6748 0.152939
R13679 gnd.n6749 gnd.n473 0.152939
R13680 gnd.n6757 gnd.n473 0.152939
R13681 gnd.n6758 gnd.n6757 0.152939
R13682 gnd.n6759 gnd.n6758 0.152939
R13683 gnd.n6759 gnd.n467 0.152939
R13684 gnd.n6767 gnd.n467 0.152939
R13685 gnd.n6768 gnd.n6767 0.152939
R13686 gnd.n6769 gnd.n6768 0.152939
R13687 gnd.n6769 gnd.n461 0.152939
R13688 gnd.n6777 gnd.n461 0.152939
R13689 gnd.n6778 gnd.n6777 0.152939
R13690 gnd.n6779 gnd.n6778 0.152939
R13691 gnd.n6779 gnd.n455 0.152939
R13692 gnd.n6787 gnd.n455 0.152939
R13693 gnd.n6788 gnd.n6787 0.152939
R13694 gnd.n6789 gnd.n6788 0.152939
R13695 gnd.n6789 gnd.n450 0.152939
R13696 gnd.n6799 gnd.n6798 0.152939
R13697 gnd.n6800 gnd.n6799 0.152939
R13698 gnd.n6800 gnd.n444 0.152939
R13699 gnd.n6808 gnd.n444 0.152939
R13700 gnd.n6809 gnd.n6808 0.152939
R13701 gnd.n6810 gnd.n6809 0.152939
R13702 gnd.n6810 gnd.n438 0.152939
R13703 gnd.n6818 gnd.n438 0.152939
R13704 gnd.n6819 gnd.n6818 0.152939
R13705 gnd.n6820 gnd.n6819 0.152939
R13706 gnd.n6820 gnd.n432 0.152939
R13707 gnd.n6828 gnd.n432 0.152939
R13708 gnd.n6829 gnd.n6828 0.152939
R13709 gnd.n6830 gnd.n6829 0.152939
R13710 gnd.n6830 gnd.n426 0.152939
R13711 gnd.n6838 gnd.n426 0.152939
R13712 gnd.n6839 gnd.n6838 0.152939
R13713 gnd.n6840 gnd.n6839 0.152939
R13714 gnd.n6840 gnd.n420 0.152939
R13715 gnd.n6848 gnd.n420 0.152939
R13716 gnd.n6849 gnd.n6848 0.152939
R13717 gnd.n6850 gnd.n6849 0.152939
R13718 gnd.n6850 gnd.n414 0.152939
R13719 gnd.n6858 gnd.n414 0.152939
R13720 gnd.n6859 gnd.n6858 0.152939
R13721 gnd.n6860 gnd.n6859 0.152939
R13722 gnd.n6860 gnd.n408 0.152939
R13723 gnd.n6868 gnd.n408 0.152939
R13724 gnd.n6869 gnd.n6868 0.152939
R13725 gnd.n6870 gnd.n6869 0.152939
R13726 gnd.n6870 gnd.n402 0.152939
R13727 gnd.n6878 gnd.n402 0.152939
R13728 gnd.n6879 gnd.n6878 0.152939
R13729 gnd.n6880 gnd.n6879 0.152939
R13730 gnd.n6880 gnd.n396 0.152939
R13731 gnd.n6888 gnd.n396 0.152939
R13732 gnd.n6889 gnd.n6888 0.152939
R13733 gnd.n6890 gnd.n6889 0.152939
R13734 gnd.n6890 gnd.n390 0.152939
R13735 gnd.n6898 gnd.n390 0.152939
R13736 gnd.n6899 gnd.n6898 0.152939
R13737 gnd.n6900 gnd.n6899 0.152939
R13738 gnd.n6900 gnd.n384 0.152939
R13739 gnd.n6908 gnd.n384 0.152939
R13740 gnd.n6909 gnd.n6908 0.152939
R13741 gnd.n6910 gnd.n6909 0.152939
R13742 gnd.n6910 gnd.n378 0.152939
R13743 gnd.n6918 gnd.n378 0.152939
R13744 gnd.n6919 gnd.n6918 0.152939
R13745 gnd.n6920 gnd.n6919 0.152939
R13746 gnd.n6920 gnd.n372 0.152939
R13747 gnd.n6928 gnd.n372 0.152939
R13748 gnd.n6929 gnd.n6928 0.152939
R13749 gnd.n6930 gnd.n6929 0.152939
R13750 gnd.n6930 gnd.n366 0.152939
R13751 gnd.n6938 gnd.n366 0.152939
R13752 gnd.n6939 gnd.n6938 0.152939
R13753 gnd.n6940 gnd.n6939 0.152939
R13754 gnd.n6940 gnd.n360 0.152939
R13755 gnd.n6948 gnd.n360 0.152939
R13756 gnd.n6949 gnd.n6948 0.152939
R13757 gnd.n6950 gnd.n6949 0.152939
R13758 gnd.n6950 gnd.n354 0.152939
R13759 gnd.n6958 gnd.n354 0.152939
R13760 gnd.n6959 gnd.n6958 0.152939
R13761 gnd.n6960 gnd.n6959 0.152939
R13762 gnd.n6960 gnd.n348 0.152939
R13763 gnd.n6968 gnd.n348 0.152939
R13764 gnd.n6969 gnd.n6968 0.152939
R13765 gnd.n6970 gnd.n6969 0.152939
R13766 gnd.n6970 gnd.n342 0.152939
R13767 gnd.n6978 gnd.n342 0.152939
R13768 gnd.n6979 gnd.n6978 0.152939
R13769 gnd.n6980 gnd.n6979 0.152939
R13770 gnd.n6980 gnd.n336 0.152939
R13771 gnd.n6988 gnd.n336 0.152939
R13772 gnd.n6989 gnd.n6988 0.152939
R13773 gnd.n6990 gnd.n6989 0.152939
R13774 gnd.n6990 gnd.n330 0.152939
R13775 gnd.n6998 gnd.n330 0.152939
R13776 gnd.n6999 gnd.n6998 0.152939
R13777 gnd.n7000 gnd.n6999 0.152939
R13778 gnd.n7000 gnd.n324 0.152939
R13779 gnd.n7008 gnd.n324 0.152939
R13780 gnd.n274 gnd.n260 0.152939
R13781 gnd.n275 gnd.n274 0.152939
R13782 gnd.n275 gnd.n273 0.152939
R13783 gnd.n281 gnd.n273 0.152939
R13784 gnd.n282 gnd.n281 0.152939
R13785 gnd.n283 gnd.n282 0.152939
R13786 gnd.n284 gnd.n283 0.152939
R13787 gnd.n285 gnd.n284 0.152939
R13788 gnd.n288 gnd.n285 0.152939
R13789 gnd.n289 gnd.n288 0.152939
R13790 gnd.n290 gnd.n289 0.152939
R13791 gnd.n291 gnd.n290 0.152939
R13792 gnd.n294 gnd.n291 0.152939
R13793 gnd.n295 gnd.n294 0.152939
R13794 gnd.n296 gnd.n295 0.152939
R13795 gnd.n297 gnd.n296 0.152939
R13796 gnd.n304 gnd.n297 0.152939
R13797 gnd.n305 gnd.n304 0.152939
R13798 gnd.n306 gnd.n305 0.152939
R13799 gnd.n307 gnd.n306 0.152939
R13800 gnd.n308 gnd.n307 0.152939
R13801 gnd.n309 gnd.n308 0.152939
R13802 gnd.n314 gnd.n309 0.152939
R13803 gnd.n315 gnd.n314 0.152939
R13804 gnd.n316 gnd.n315 0.152939
R13805 gnd.n317 gnd.n316 0.152939
R13806 gnd.n322 gnd.n317 0.152939
R13807 gnd.n323 gnd.n322 0.152939
R13808 gnd.n7009 gnd.n323 0.152939
R13809 gnd.n7119 gnd.n7118 0.152939
R13810 gnd.n7119 gnd.n208 0.152939
R13811 gnd.n7133 gnd.n208 0.152939
R13812 gnd.n7134 gnd.n7133 0.152939
R13813 gnd.n7135 gnd.n7134 0.152939
R13814 gnd.n7135 gnd.n192 0.152939
R13815 gnd.n7149 gnd.n192 0.152939
R13816 gnd.n7150 gnd.n7149 0.152939
R13817 gnd.n7151 gnd.n7150 0.152939
R13818 gnd.n7151 gnd.n176 0.152939
R13819 gnd.n7165 gnd.n176 0.152939
R13820 gnd.n7166 gnd.n7165 0.152939
R13821 gnd.n7167 gnd.n7166 0.152939
R13822 gnd.n7168 gnd.n7167 0.152939
R13823 gnd.n7168 gnd.n88 0.152939
R13824 gnd.n7323 gnd.n88 0.152939
R13825 gnd.n7322 gnd.n89 0.152939
R13826 gnd.n91 gnd.n89 0.152939
R13827 gnd.n96 gnd.n91 0.152939
R13828 gnd.n97 gnd.n96 0.152939
R13829 gnd.n98 gnd.n97 0.152939
R13830 gnd.n99 gnd.n98 0.152939
R13831 gnd.n103 gnd.n99 0.152939
R13832 gnd.n104 gnd.n103 0.152939
R13833 gnd.n105 gnd.n104 0.152939
R13834 gnd.n106 gnd.n105 0.152939
R13835 gnd.n110 gnd.n106 0.152939
R13836 gnd.n111 gnd.n110 0.152939
R13837 gnd.n112 gnd.n111 0.152939
R13838 gnd.n113 gnd.n112 0.152939
R13839 gnd.n117 gnd.n113 0.152939
R13840 gnd.n118 gnd.n117 0.152939
R13841 gnd.n119 gnd.n118 0.152939
R13842 gnd.n120 gnd.n119 0.152939
R13843 gnd.n124 gnd.n120 0.152939
R13844 gnd.n125 gnd.n124 0.152939
R13845 gnd.n126 gnd.n125 0.152939
R13846 gnd.n127 gnd.n126 0.152939
R13847 gnd.n131 gnd.n127 0.152939
R13848 gnd.n132 gnd.n131 0.152939
R13849 gnd.n133 gnd.n132 0.152939
R13850 gnd.n134 gnd.n133 0.152939
R13851 gnd.n138 gnd.n134 0.152939
R13852 gnd.n139 gnd.n138 0.152939
R13853 gnd.n140 gnd.n139 0.152939
R13854 gnd.n141 gnd.n140 0.152939
R13855 gnd.n145 gnd.n141 0.152939
R13856 gnd.n146 gnd.n145 0.152939
R13857 gnd.n147 gnd.n146 0.152939
R13858 gnd.n148 gnd.n147 0.152939
R13859 gnd.n152 gnd.n148 0.152939
R13860 gnd.n153 gnd.n152 0.152939
R13861 gnd.n7253 gnd.n153 0.152939
R13862 gnd.n7253 gnd.n7252 0.152939
R13863 gnd.n4151 gnd.n1595 0.152939
R13864 gnd.n4152 gnd.n4151 0.152939
R13865 gnd.n4153 gnd.n4152 0.152939
R13866 gnd.n4154 gnd.n4153 0.152939
R13867 gnd.n4155 gnd.n4154 0.152939
R13868 gnd.n4156 gnd.n4155 0.152939
R13869 gnd.n4157 gnd.n4156 0.152939
R13870 gnd.n4158 gnd.n4157 0.152939
R13871 gnd.n4159 gnd.n4158 0.152939
R13872 gnd.n4160 gnd.n4159 0.152939
R13873 gnd.n4161 gnd.n4160 0.152939
R13874 gnd.n4161 gnd.n1526 0.152939
R13875 gnd.n4263 gnd.n1526 0.152939
R13876 gnd.n4264 gnd.n4263 0.152939
R13877 gnd.n4265 gnd.n4264 0.152939
R13878 gnd.n4265 gnd.n1524 0.152939
R13879 gnd.n4271 gnd.n1524 0.152939
R13880 gnd.n4272 gnd.n4271 0.152939
R13881 gnd.n4273 gnd.n4272 0.152939
R13882 gnd.n4274 gnd.n4273 0.152939
R13883 gnd.n4275 gnd.n4274 0.152939
R13884 gnd.n4276 gnd.n4275 0.152939
R13885 gnd.n4277 gnd.n4276 0.152939
R13886 gnd.n4278 gnd.n4277 0.152939
R13887 gnd.n4279 gnd.n4278 0.152939
R13888 gnd.n4281 gnd.n4279 0.152939
R13889 gnd.n4281 gnd.n4280 0.152939
R13890 gnd.n4280 gnd.n264 0.152939
R13891 gnd.n265 gnd.n264 0.152939
R13892 gnd.n266 gnd.n265 0.152939
R13893 gnd.n267 gnd.n266 0.152939
R13894 gnd.n268 gnd.n267 0.152939
R13895 gnd.n7047 gnd.n268 0.152939
R13896 gnd.n7051 gnd.n7047 0.152939
R13897 gnd.n7052 gnd.n7051 0.152939
R13898 gnd.n7053 gnd.n7052 0.152939
R13899 gnd.n7054 gnd.n7053 0.152939
R13900 gnd.n7055 gnd.n7054 0.152939
R13901 gnd.n7057 gnd.n7055 0.152939
R13902 gnd.n7057 gnd.n7056 0.152939
R13903 gnd.n7056 gnd.n159 0.152939
R13904 gnd.n7251 gnd.n159 0.152939
R13905 gnd.n1844 gnd.n1839 0.152939
R13906 gnd.n1845 gnd.n1844 0.152939
R13907 gnd.n1846 gnd.n1845 0.152939
R13908 gnd.n1846 gnd.n1835 0.152939
R13909 gnd.n1854 gnd.n1835 0.152939
R13910 gnd.n1855 gnd.n1854 0.152939
R13911 gnd.n1856 gnd.n1855 0.152939
R13912 gnd.n1856 gnd.n1831 0.152939
R13913 gnd.n1864 gnd.n1831 0.152939
R13914 gnd.n1865 gnd.n1864 0.152939
R13915 gnd.n1867 gnd.n1865 0.152939
R13916 gnd.n1867 gnd.n1866 0.152939
R13917 gnd.n1866 gnd.n1824 0.152939
R13918 gnd.n1876 gnd.n1824 0.152939
R13919 gnd.n1877 gnd.n1876 0.152939
R13920 gnd.n1884 gnd.n1881 0.152939
R13921 gnd.n1885 gnd.n1884 0.152939
R13922 gnd.n1886 gnd.n1885 0.152939
R13923 gnd.n1887 gnd.n1886 0.152939
R13924 gnd.n1890 gnd.n1887 0.152939
R13925 gnd.n1891 gnd.n1890 0.152939
R13926 gnd.n1892 gnd.n1891 0.152939
R13927 gnd.n1893 gnd.n1892 0.152939
R13928 gnd.n1896 gnd.n1893 0.152939
R13929 gnd.n1897 gnd.n1896 0.152939
R13930 gnd.n1898 gnd.n1897 0.152939
R13931 gnd.n1899 gnd.n1898 0.152939
R13932 gnd.n1902 gnd.n1899 0.152939
R13933 gnd.n1903 gnd.n1902 0.152939
R13934 gnd.n1904 gnd.n1903 0.152939
R13935 gnd.n1905 gnd.n1904 0.152939
R13936 gnd.n1911 gnd.n1905 0.152939
R13937 gnd.n1917 gnd.n1911 0.152939
R13938 gnd.n1917 gnd.n1916 0.152939
R13939 gnd.n1916 gnd.n1915 0.152939
R13940 gnd.n1467 gnd.n1466 0.152939
R13941 gnd.n1468 gnd.n1467 0.152939
R13942 gnd.n1582 gnd.n1468 0.152939
R13943 gnd.n1583 gnd.n1582 0.152939
R13944 gnd.n1583 gnd.n1561 0.152939
R13945 gnd.n4200 gnd.n1561 0.152939
R13946 gnd.n4201 gnd.n4200 0.152939
R13947 gnd.n4202 gnd.n4201 0.152939
R13948 gnd.n4203 gnd.n4202 0.152939
R13949 gnd.n4203 gnd.n1536 0.152939
R13950 gnd.n4253 gnd.n1536 0.152939
R13951 gnd.n4254 gnd.n4253 0.152939
R13952 gnd.n4255 gnd.n4254 0.152939
R13953 gnd.n4256 gnd.n4255 0.152939
R13954 gnd.n4256 gnd.n224 0.152939
R13955 gnd.n7118 gnd.n224 0.152939
R13956 gnd.n2901 gnd.n2900 0.152939
R13957 gnd.n2902 gnd.n2901 0.152939
R13958 gnd.n2902 gnd.n2574 0.152939
R13959 gnd.n2964 gnd.n2574 0.152939
R13960 gnd.n2965 gnd.n2964 0.152939
R13961 gnd.n2966 gnd.n2965 0.152939
R13962 gnd.n2966 gnd.n2570 0.152939
R13963 gnd.n2972 gnd.n2570 0.152939
R13964 gnd.n2973 gnd.n2972 0.152939
R13965 gnd.n2974 gnd.n2973 0.152939
R13966 gnd.n2974 gnd.n2566 0.152939
R13967 gnd.n2980 gnd.n2566 0.152939
R13968 gnd.n2981 gnd.n2980 0.152939
R13969 gnd.n2982 gnd.n2981 0.152939
R13970 gnd.n2982 gnd.n2562 0.152939
R13971 gnd.n2988 gnd.n2562 0.152939
R13972 gnd.n2989 gnd.n2988 0.152939
R13973 gnd.n2990 gnd.n2989 0.152939
R13974 gnd.n2990 gnd.n2556 0.152939
R13975 gnd.n3131 gnd.n2556 0.152939
R13976 gnd.n3132 gnd.n3131 0.152939
R13977 gnd.n3133 gnd.n3132 0.152939
R13978 gnd.n3133 gnd.n2550 0.152939
R13979 gnd.n3145 gnd.n2550 0.152939
R13980 gnd.n3146 gnd.n3145 0.152939
R13981 gnd.n3147 gnd.n3146 0.152939
R13982 gnd.n3147 gnd.n2542 0.152939
R13983 gnd.n3159 gnd.n2542 0.152939
R13984 gnd.n3160 gnd.n3159 0.152939
R13985 gnd.n3161 gnd.n3160 0.152939
R13986 gnd.n3161 gnd.n2534 0.152939
R13987 gnd.n3173 gnd.n2534 0.152939
R13988 gnd.n3174 gnd.n3173 0.152939
R13989 gnd.n3175 gnd.n3174 0.152939
R13990 gnd.n3175 gnd.n2257 0.152939
R13991 gnd.n3362 gnd.n2257 0.152939
R13992 gnd.n3363 gnd.n3362 0.152939
R13993 gnd.n3364 gnd.n3363 0.152939
R13994 gnd.n3364 gnd.n2239 0.152939
R13995 gnd.n3453 gnd.n2239 0.152939
R13996 gnd.n3454 gnd.n3453 0.152939
R13997 gnd.n3455 gnd.n3454 0.152939
R13998 gnd.n3455 gnd.n2218 0.152939
R13999 gnd.n3484 gnd.n2218 0.152939
R14000 gnd.n3485 gnd.n3484 0.152939
R14001 gnd.n3486 gnd.n3485 0.152939
R14002 gnd.n3486 gnd.n2196 0.152939
R14003 gnd.n3512 gnd.n2196 0.152939
R14004 gnd.n3513 gnd.n3512 0.152939
R14005 gnd.n3514 gnd.n3513 0.152939
R14006 gnd.n3515 gnd.n3514 0.152939
R14007 gnd.n3515 gnd.n2167 0.152939
R14008 gnd.n3549 gnd.n2167 0.152939
R14009 gnd.n3550 gnd.n3549 0.152939
R14010 gnd.n3551 gnd.n3550 0.152939
R14011 gnd.n3551 gnd.n2144 0.152939
R14012 gnd.n3577 gnd.n2144 0.152939
R14013 gnd.n3578 gnd.n3577 0.152939
R14014 gnd.n3579 gnd.n3578 0.152939
R14015 gnd.n3580 gnd.n3579 0.152939
R14016 gnd.n3580 gnd.n2115 0.152939
R14017 gnd.n3628 gnd.n2115 0.152939
R14018 gnd.n3629 gnd.n3628 0.152939
R14019 gnd.n3630 gnd.n3629 0.152939
R14020 gnd.n3630 gnd.n2094 0.152939
R14021 gnd.n3658 gnd.n2094 0.152939
R14022 gnd.n3659 gnd.n3658 0.152939
R14023 gnd.n3660 gnd.n3659 0.152939
R14024 gnd.n3661 gnd.n3660 0.152939
R14025 gnd.n3661 gnd.n2064 0.152939
R14026 gnd.n3708 gnd.n2064 0.152939
R14027 gnd.n3709 gnd.n3708 0.152939
R14028 gnd.n3710 gnd.n3709 0.152939
R14029 gnd.n3710 gnd.n2041 0.152939
R14030 gnd.n3748 gnd.n2041 0.152939
R14031 gnd.n3749 gnd.n3748 0.152939
R14032 gnd.n3750 gnd.n3749 0.152939
R14033 gnd.n3750 gnd.n2018 0.152939
R14034 gnd.n3787 gnd.n2018 0.152939
R14035 gnd.n3788 gnd.n3787 0.152939
R14036 gnd.n3789 gnd.n3788 0.152939
R14037 gnd.n3789 gnd.n1996 0.152939
R14038 gnd.n3828 gnd.n1996 0.152939
R14039 gnd.n3829 gnd.n3828 0.152939
R14040 gnd.n3830 gnd.n3829 0.152939
R14041 gnd.n3830 gnd.n1974 0.152939
R14042 gnd.n3873 gnd.n1974 0.152939
R14043 gnd.n3874 gnd.n3873 0.152939
R14044 gnd.n3875 gnd.n3874 0.152939
R14045 gnd.n3876 gnd.n3875 0.152939
R14046 gnd.n3877 gnd.n3876 0.152939
R14047 gnd.n3877 gnd.n1778 0.152939
R14048 gnd.n4064 gnd.n1778 0.152939
R14049 gnd.n4065 gnd.n4064 0.152939
R14050 gnd.n4066 gnd.n4065 0.152939
R14051 gnd.n4066 gnd.n1766 0.152939
R14052 gnd.n4085 gnd.n1766 0.152939
R14053 gnd.n4086 gnd.n4085 0.152939
R14054 gnd.n4087 gnd.n4086 0.152939
R14055 gnd.n4087 gnd.n1754 0.152939
R14056 gnd.n4108 gnd.n1754 0.152939
R14057 gnd.n4109 gnd.n4108 0.152939
R14058 gnd.n4111 gnd.n4109 0.152939
R14059 gnd.n4111 gnd.n4110 0.152939
R14060 gnd.n4110 gnd.n1445 0.152939
R14061 gnd.n1446 gnd.n1445 0.152939
R14062 gnd.n1447 gnd.n1446 0.152939
R14063 gnd.n1453 gnd.n1447 0.152939
R14064 gnd.n1454 gnd.n1453 0.152939
R14065 gnd.n1455 gnd.n1454 0.152939
R14066 gnd.n1456 gnd.n1455 0.152939
R14067 gnd.n1576 gnd.n1456 0.152939
R14068 gnd.n1577 gnd.n1576 0.152939
R14069 gnd.n1578 gnd.n1577 0.152939
R14070 gnd.n1578 gnd.n1572 0.152939
R14071 gnd.n4189 gnd.n1572 0.152939
R14072 gnd.n4190 gnd.n4189 0.152939
R14073 gnd.n4191 gnd.n4190 0.152939
R14074 gnd.n4192 gnd.n4191 0.152939
R14075 gnd.n4192 gnd.n1545 0.152939
R14076 gnd.n4226 gnd.n1545 0.152939
R14077 gnd.n4227 gnd.n4226 0.152939
R14078 gnd.n4228 gnd.n4227 0.152939
R14079 gnd.n4229 gnd.n4228 0.152939
R14080 gnd.n4230 gnd.n4229 0.152939
R14081 gnd.n4233 gnd.n4230 0.152939
R14082 gnd.n4234 gnd.n4233 0.152939
R14083 gnd.n2730 gnd.n2729 0.152939
R14084 gnd.n2731 gnd.n2730 0.152939
R14085 gnd.n2732 gnd.n2731 0.152939
R14086 gnd.n2733 gnd.n2732 0.152939
R14087 gnd.n2734 gnd.n2733 0.152939
R14088 gnd.n2735 gnd.n2734 0.152939
R14089 gnd.n2735 gnd.n2650 0.152939
R14090 gnd.n2811 gnd.n2650 0.152939
R14091 gnd.n2812 gnd.n2811 0.152939
R14092 gnd.n2813 gnd.n2812 0.152939
R14093 gnd.n2813 gnd.n2643 0.152939
R14094 gnd.n2828 gnd.n2643 0.152939
R14095 gnd.n2829 gnd.n2828 0.152939
R14096 gnd.n2830 gnd.n2829 0.152939
R14097 gnd.n2832 gnd.n2830 0.152939
R14098 gnd.n2832 gnd.n2831 0.152939
R14099 gnd.n2831 gnd.n2615 0.152939
R14100 gnd.n2616 gnd.n2615 0.152939
R14101 gnd.n2617 gnd.n2616 0.152939
R14102 gnd.n2850 gnd.n2617 0.152939
R14103 gnd.n2685 gnd.n2684 0.152939
R14104 gnd.n2691 gnd.n2684 0.152939
R14105 gnd.n2692 gnd.n2691 0.152939
R14106 gnd.n2693 gnd.n2692 0.152939
R14107 gnd.n2693 gnd.n2682 0.152939
R14108 gnd.n2701 gnd.n2682 0.152939
R14109 gnd.n2702 gnd.n2701 0.152939
R14110 gnd.n2703 gnd.n2702 0.152939
R14111 gnd.n2703 gnd.n2680 0.152939
R14112 gnd.n2711 gnd.n2680 0.152939
R14113 gnd.n2712 gnd.n2711 0.152939
R14114 gnd.n2713 gnd.n2712 0.152939
R14115 gnd.n2713 gnd.n2678 0.152939
R14116 gnd.n2721 gnd.n2678 0.152939
R14117 gnd.n2722 gnd.n2721 0.152939
R14118 gnd.n2723 gnd.n2722 0.152939
R14119 gnd.n2723 gnd.n2671 0.152939
R14120 gnd.n2727 gnd.n2671 0.152939
R14121 gnd.n4631 gnd.n1124 0.152939
R14122 gnd.n4631 gnd.n4630 0.152939
R14123 gnd.n4630 gnd.n4629 0.152939
R14124 gnd.n4629 gnd.n1126 0.152939
R14125 gnd.n1147 gnd.n1126 0.152939
R14126 gnd.n1148 gnd.n1147 0.152939
R14127 gnd.n1149 gnd.n1148 0.152939
R14128 gnd.n1166 gnd.n1149 0.152939
R14129 gnd.n1167 gnd.n1166 0.152939
R14130 gnd.n1168 gnd.n1167 0.152939
R14131 gnd.n1169 gnd.n1168 0.152939
R14132 gnd.n1188 gnd.n1169 0.152939
R14133 gnd.n1189 gnd.n1188 0.152939
R14134 gnd.n1190 gnd.n1189 0.152939
R14135 gnd.n1191 gnd.n1190 0.152939
R14136 gnd.n1211 gnd.n1191 0.152939
R14137 gnd.n1212 gnd.n1211 0.152939
R14138 gnd.n1213 gnd.n1212 0.152939
R14139 gnd.n1214 gnd.n1213 0.152939
R14140 gnd.n1215 gnd.n1214 0.152939
R14141 gnd.n2636 gnd.n1215 0.152939
R14142 gnd.n2636 gnd.n1229 0.152939
R14143 gnd.n1230 gnd.n1229 0.152939
R14144 gnd.n1231 gnd.n1230 0.152939
R14145 gnd.n1247 gnd.n1231 0.152939
R14146 gnd.n1248 gnd.n1247 0.152939
R14147 gnd.n1249 gnd.n1248 0.152939
R14148 gnd.n1250 gnd.n1249 0.152939
R14149 gnd.n1267 gnd.n1250 0.152939
R14150 gnd.n1268 gnd.n1267 0.152939
R14151 gnd.n1269 gnd.n1268 0.152939
R14152 gnd.n1270 gnd.n1269 0.152939
R14153 gnd.n1289 gnd.n1270 0.152939
R14154 gnd.n1290 gnd.n1289 0.152939
R14155 gnd.n1291 gnd.n1290 0.152939
R14156 gnd.n1292 gnd.n1291 0.152939
R14157 gnd.n1310 gnd.n1292 0.152939
R14158 gnd.n1311 gnd.n1310 0.152939
R14159 gnd.n1312 gnd.n1311 0.152939
R14160 gnd.n1313 gnd.n1312 0.152939
R14161 gnd.n1331 gnd.n1313 0.152939
R14162 gnd.n4505 gnd.n1331 0.152939
R14163 gnd.n1257 gnd.n1200 0.152939
R14164 gnd.n1258 gnd.n1257 0.152939
R14165 gnd.n1259 gnd.n1258 0.152939
R14166 gnd.n1260 gnd.n1259 0.152939
R14167 gnd.n1278 gnd.n1260 0.152939
R14168 gnd.n1279 gnd.n1278 0.152939
R14169 gnd.n1280 gnd.n1279 0.152939
R14170 gnd.n1281 gnd.n1280 0.152939
R14171 gnd.n1299 gnd.n1281 0.152939
R14172 gnd.n1300 gnd.n1299 0.152939
R14173 gnd.n1301 gnd.n1300 0.152939
R14174 gnd.n1302 gnd.n1301 0.152939
R14175 gnd.n1321 gnd.n1302 0.152939
R14176 gnd.n1322 gnd.n1321 0.152939
R14177 gnd.n1323 gnd.n1322 0.152939
R14178 gnd.n1324 gnd.n1323 0.152939
R14179 gnd.n2418 gnd.n2417 0.152939
R14180 gnd.n2419 gnd.n2418 0.152939
R14181 gnd.n2420 gnd.n2419 0.152939
R14182 gnd.n2421 gnd.n2420 0.152939
R14183 gnd.n2422 gnd.n2421 0.152939
R14184 gnd.n2423 gnd.n2422 0.152939
R14185 gnd.n2424 gnd.n2423 0.152939
R14186 gnd.n2425 gnd.n2424 0.152939
R14187 gnd.n2426 gnd.n2425 0.152939
R14188 gnd.n2427 gnd.n2426 0.152939
R14189 gnd.n2428 gnd.n2427 0.152939
R14190 gnd.n2429 gnd.n2428 0.152939
R14191 gnd.n2430 gnd.n2429 0.152939
R14192 gnd.n2431 gnd.n2430 0.152939
R14193 gnd.n2431 gnd.n2401 0.152939
R14194 gnd.n3282 gnd.n3281 0.152939
R14195 gnd.n3281 gnd.n2402 0.152939
R14196 gnd.n2462 gnd.n2402 0.152939
R14197 gnd.n2463 gnd.n2462 0.152939
R14198 gnd.n2464 gnd.n2463 0.152939
R14199 gnd.n2465 gnd.n2464 0.152939
R14200 gnd.n2469 gnd.n2465 0.152939
R14201 gnd.n2470 gnd.n2469 0.152939
R14202 gnd.n2471 gnd.n2470 0.152939
R14203 gnd.n2472 gnd.n2471 0.152939
R14204 gnd.n2476 gnd.n2472 0.152939
R14205 gnd.n2477 gnd.n2476 0.152939
R14206 gnd.n2478 gnd.n2477 0.152939
R14207 gnd.n2479 gnd.n2478 0.152939
R14208 gnd.n2483 gnd.n2479 0.152939
R14209 gnd.n2484 gnd.n2483 0.152939
R14210 gnd.n2485 gnd.n2484 0.152939
R14211 gnd.n2486 gnd.n2485 0.152939
R14212 gnd.n2491 gnd.n2486 0.152939
R14213 gnd.n3244 gnd.n2491 0.152939
R14214 gnd.n2739 gnd.n1116 0.152939
R14215 gnd.n2742 gnd.n2739 0.152939
R14216 gnd.n2743 gnd.n2742 0.152939
R14217 gnd.n2744 gnd.n2743 0.152939
R14218 gnd.n2744 gnd.n2653 0.152939
R14219 gnd.n2803 gnd.n2653 0.152939
R14220 gnd.n2804 gnd.n2803 0.152939
R14221 gnd.n2805 gnd.n2804 0.152939
R14222 gnd.n2805 gnd.n2646 0.152939
R14223 gnd.n2819 gnd.n2646 0.152939
R14224 gnd.n2820 gnd.n2819 0.152939
R14225 gnd.n2822 gnd.n2820 0.152939
R14226 gnd.n2822 gnd.n2821 0.152939
R14227 gnd.n2821 gnd.n2640 0.152939
R14228 gnd.n2841 gnd.n2640 0.152939
R14229 gnd.n2842 gnd.n2841 0.152939
R14230 gnd.n2843 gnd.n2842 0.152939
R14231 gnd.n2843 gnd.n2637 0.152939
R14232 gnd.n2847 gnd.n2637 0.152939
R14233 gnd.n2848 gnd.n2847 0.152939
R14234 gnd.n2849 gnd.n2848 0.152939
R14235 gnd.n2849 gnd.n2634 0.152939
R14236 gnd.n2859 gnd.n2634 0.152939
R14237 gnd.n2860 gnd.n2859 0.152939
R14238 gnd.n2861 gnd.n2860 0.152939
R14239 gnd.n2862 gnd.n2861 0.152939
R14240 gnd.n2863 gnd.n2862 0.152939
R14241 gnd.n2863 gnd.n2592 0.152939
R14242 gnd.n2918 gnd.n2592 0.152939
R14243 gnd.n2919 gnd.n2918 0.152939
R14244 gnd.n2920 gnd.n2919 0.152939
R14245 gnd.n2920 gnd.n2590 0.152939
R14246 gnd.n2926 gnd.n2590 0.152939
R14247 gnd.n2927 gnd.n2926 0.152939
R14248 gnd.n2928 gnd.n2927 0.152939
R14249 gnd.n2928 gnd.n2588 0.152939
R14250 gnd.n2937 gnd.n2588 0.152939
R14251 gnd.n2938 gnd.n2937 0.152939
R14252 gnd.n2940 gnd.n2938 0.152939
R14253 gnd.n2940 gnd.n2939 0.152939
R14254 gnd.n2939 gnd.n2492 0.152939
R14255 gnd.n3243 gnd.n2492 0.152939
R14256 gnd.n1074 gnd.n1073 0.152939
R14257 gnd.n1075 gnd.n1074 0.152939
R14258 gnd.n1076 gnd.n1075 0.152939
R14259 gnd.n1077 gnd.n1076 0.152939
R14260 gnd.n1078 gnd.n1077 0.152939
R14261 gnd.n1079 gnd.n1078 0.152939
R14262 gnd.n1080 gnd.n1079 0.152939
R14263 gnd.n1081 gnd.n1080 0.152939
R14264 gnd.n1082 gnd.n1081 0.152939
R14265 gnd.n1083 gnd.n1082 0.152939
R14266 gnd.n1084 gnd.n1083 0.152939
R14267 gnd.n1085 gnd.n1084 0.152939
R14268 gnd.n1086 gnd.n1085 0.152939
R14269 gnd.n1087 gnd.n1086 0.152939
R14270 gnd.n1088 gnd.n1087 0.152939
R14271 gnd.n1089 gnd.n1088 0.152939
R14272 gnd.n1090 gnd.n1089 0.152939
R14273 gnd.n1093 gnd.n1090 0.152939
R14274 gnd.n1094 gnd.n1093 0.152939
R14275 gnd.n1095 gnd.n1094 0.152939
R14276 gnd.n1096 gnd.n1095 0.152939
R14277 gnd.n1097 gnd.n1096 0.152939
R14278 gnd.n1098 gnd.n1097 0.152939
R14279 gnd.n1099 gnd.n1098 0.152939
R14280 gnd.n1100 gnd.n1099 0.152939
R14281 gnd.n1101 gnd.n1100 0.152939
R14282 gnd.n1102 gnd.n1101 0.152939
R14283 gnd.n1103 gnd.n1102 0.152939
R14284 gnd.n1104 gnd.n1103 0.152939
R14285 gnd.n1105 gnd.n1104 0.152939
R14286 gnd.n1106 gnd.n1105 0.152939
R14287 gnd.n1107 gnd.n1106 0.152939
R14288 gnd.n1108 gnd.n1107 0.152939
R14289 gnd.n1109 gnd.n1108 0.152939
R14290 gnd.n1110 gnd.n1109 0.152939
R14291 gnd.n4641 gnd.n1110 0.152939
R14292 gnd.n4641 gnd.n4640 0.152939
R14293 gnd.n4640 gnd.n4639 0.152939
R14294 gnd.n2664 gnd.n2662 0.152939
R14295 gnd.n2664 gnd.n2663 0.152939
R14296 gnd.n2663 gnd.n1137 0.152939
R14297 gnd.n1138 gnd.n1137 0.152939
R14298 gnd.n1139 gnd.n1138 0.152939
R14299 gnd.n1156 gnd.n1139 0.152939
R14300 gnd.n1157 gnd.n1156 0.152939
R14301 gnd.n1158 gnd.n1157 0.152939
R14302 gnd.n1159 gnd.n1158 0.152939
R14303 gnd.n1177 gnd.n1159 0.152939
R14304 gnd.n1178 gnd.n1177 0.152939
R14305 gnd.n1179 gnd.n1178 0.152939
R14306 gnd.n1180 gnd.n1179 0.152939
R14307 gnd.n1198 gnd.n1180 0.152939
R14308 gnd.n1199 gnd.n1198 0.152939
R14309 gnd.n1200 gnd.n1199 0.152939
R14310 gnd.n1021 gnd.n1020 0.152939
R14311 gnd.n1022 gnd.n1021 0.152939
R14312 gnd.n1027 gnd.n1022 0.152939
R14313 gnd.n1028 gnd.n1027 0.152939
R14314 gnd.n1029 gnd.n1028 0.152939
R14315 gnd.n1030 gnd.n1029 0.152939
R14316 gnd.n1035 gnd.n1030 0.152939
R14317 gnd.n1036 gnd.n1035 0.152939
R14318 gnd.n1037 gnd.n1036 0.152939
R14319 gnd.n1038 gnd.n1037 0.152939
R14320 gnd.n2759 gnd.n1038 0.152939
R14321 gnd.n2760 gnd.n2759 0.152939
R14322 gnd.n2760 gnd.n2757 0.152939
R14323 gnd.n2766 gnd.n2757 0.152939
R14324 gnd.n2767 gnd.n2766 0.152939
R14325 gnd.n2768 gnd.n2767 0.152939
R14326 gnd.n2768 gnd.n2659 0.152939
R14327 gnd.n2774 gnd.n2659 0.152939
R14328 gnd.n2775 gnd.n2774 0.152939
R14329 gnd.n2776 gnd.n2775 0.152939
R14330 gnd.n2777 gnd.n2776 0.152939
R14331 gnd.n2778 gnd.n2777 0.152939
R14332 gnd.n2781 gnd.n2778 0.152939
R14333 gnd.n2782 gnd.n2781 0.152939
R14334 gnd.n2783 gnd.n2782 0.152939
R14335 gnd.n2784 gnd.n2783 0.152939
R14336 gnd.n2785 gnd.n2784 0.152939
R14337 gnd.n2785 gnd.n2606 0.152939
R14338 gnd.n2898 gnd.n2606 0.152939
R14339 gnd.n766 gnd.n761 0.152939
R14340 gnd.n767 gnd.n766 0.152939
R14341 gnd.n768 gnd.n767 0.152939
R14342 gnd.n773 gnd.n768 0.152939
R14343 gnd.n774 gnd.n773 0.152939
R14344 gnd.n775 gnd.n774 0.152939
R14345 gnd.n776 gnd.n775 0.152939
R14346 gnd.n781 gnd.n776 0.152939
R14347 gnd.n782 gnd.n781 0.152939
R14348 gnd.n783 gnd.n782 0.152939
R14349 gnd.n784 gnd.n783 0.152939
R14350 gnd.n789 gnd.n784 0.152939
R14351 gnd.n790 gnd.n789 0.152939
R14352 gnd.n791 gnd.n790 0.152939
R14353 gnd.n792 gnd.n791 0.152939
R14354 gnd.n797 gnd.n792 0.152939
R14355 gnd.n798 gnd.n797 0.152939
R14356 gnd.n799 gnd.n798 0.152939
R14357 gnd.n800 gnd.n799 0.152939
R14358 gnd.n805 gnd.n800 0.152939
R14359 gnd.n806 gnd.n805 0.152939
R14360 gnd.n807 gnd.n806 0.152939
R14361 gnd.n808 gnd.n807 0.152939
R14362 gnd.n813 gnd.n808 0.152939
R14363 gnd.n814 gnd.n813 0.152939
R14364 gnd.n815 gnd.n814 0.152939
R14365 gnd.n816 gnd.n815 0.152939
R14366 gnd.n821 gnd.n816 0.152939
R14367 gnd.n822 gnd.n821 0.152939
R14368 gnd.n823 gnd.n822 0.152939
R14369 gnd.n824 gnd.n823 0.152939
R14370 gnd.n829 gnd.n824 0.152939
R14371 gnd.n830 gnd.n829 0.152939
R14372 gnd.n831 gnd.n830 0.152939
R14373 gnd.n832 gnd.n831 0.152939
R14374 gnd.n837 gnd.n832 0.152939
R14375 gnd.n838 gnd.n837 0.152939
R14376 gnd.n839 gnd.n838 0.152939
R14377 gnd.n840 gnd.n839 0.152939
R14378 gnd.n845 gnd.n840 0.152939
R14379 gnd.n846 gnd.n845 0.152939
R14380 gnd.n847 gnd.n846 0.152939
R14381 gnd.n848 gnd.n847 0.152939
R14382 gnd.n853 gnd.n848 0.152939
R14383 gnd.n854 gnd.n853 0.152939
R14384 gnd.n855 gnd.n854 0.152939
R14385 gnd.n856 gnd.n855 0.152939
R14386 gnd.n861 gnd.n856 0.152939
R14387 gnd.n862 gnd.n861 0.152939
R14388 gnd.n863 gnd.n862 0.152939
R14389 gnd.n864 gnd.n863 0.152939
R14390 gnd.n869 gnd.n864 0.152939
R14391 gnd.n870 gnd.n869 0.152939
R14392 gnd.n871 gnd.n870 0.152939
R14393 gnd.n872 gnd.n871 0.152939
R14394 gnd.n877 gnd.n872 0.152939
R14395 gnd.n878 gnd.n877 0.152939
R14396 gnd.n879 gnd.n878 0.152939
R14397 gnd.n880 gnd.n879 0.152939
R14398 gnd.n885 gnd.n880 0.152939
R14399 gnd.n886 gnd.n885 0.152939
R14400 gnd.n887 gnd.n886 0.152939
R14401 gnd.n888 gnd.n887 0.152939
R14402 gnd.n893 gnd.n888 0.152939
R14403 gnd.n894 gnd.n893 0.152939
R14404 gnd.n895 gnd.n894 0.152939
R14405 gnd.n896 gnd.n895 0.152939
R14406 gnd.n901 gnd.n896 0.152939
R14407 gnd.n902 gnd.n901 0.152939
R14408 gnd.n903 gnd.n902 0.152939
R14409 gnd.n904 gnd.n903 0.152939
R14410 gnd.n909 gnd.n904 0.152939
R14411 gnd.n910 gnd.n909 0.152939
R14412 gnd.n911 gnd.n910 0.152939
R14413 gnd.n912 gnd.n911 0.152939
R14414 gnd.n917 gnd.n912 0.152939
R14415 gnd.n918 gnd.n917 0.152939
R14416 gnd.n919 gnd.n918 0.152939
R14417 gnd.n920 gnd.n919 0.152939
R14418 gnd.n925 gnd.n920 0.152939
R14419 gnd.n926 gnd.n925 0.152939
R14420 gnd.n927 gnd.n926 0.152939
R14421 gnd.n928 gnd.n927 0.152939
R14422 gnd.n1019 gnd.n928 0.152939
R14423 gnd.n4142 gnd.n1599 0.152939
R14424 gnd.n4138 gnd.n1599 0.152939
R14425 gnd.n4138 gnd.n4137 0.152939
R14426 gnd.n4137 gnd.n4136 0.152939
R14427 gnd.n4136 gnd.n1741 0.152939
R14428 gnd.n4129 gnd.n1741 0.152939
R14429 gnd.n4129 gnd.n4128 0.152939
R14430 gnd.n4128 gnd.n4127 0.152939
R14431 gnd.n4127 gnd.n4120 0.152939
R14432 gnd.n3216 gnd.n2516 0.152939
R14433 gnd.n3212 gnd.n2516 0.152939
R14434 gnd.n3212 gnd.n3211 0.152939
R14435 gnd.n3211 gnd.n3210 0.152939
R14436 gnd.n3210 gnd.n2521 0.152939
R14437 gnd.n3206 gnd.n2521 0.152939
R14438 gnd.n3206 gnd.n3205 0.152939
R14439 gnd.n3205 gnd.n3204 0.152939
R14440 gnd.n3204 gnd.n2526 0.152939
R14441 gnd.n3200 gnd.n2526 0.152939
R14442 gnd.n3200 gnd.n3199 0.152939
R14443 gnd.n3199 gnd.n3198 0.152939
R14444 gnd.n3198 gnd.n2531 0.152939
R14445 gnd.n3194 gnd.n2531 0.152939
R14446 gnd.n3194 gnd.n3193 0.152939
R14447 gnd.n3193 gnd.n3192 0.152939
R14448 gnd.n3192 gnd.n3186 0.152939
R14449 gnd.n3186 gnd.n2231 0.152939
R14450 gnd.n3463 gnd.n2231 0.152939
R14451 gnd.n3464 gnd.n3463 0.152939
R14452 gnd.n3465 gnd.n3464 0.152939
R14453 gnd.n3465 gnd.n2211 0.152939
R14454 gnd.n3494 gnd.n2211 0.152939
R14455 gnd.n3495 gnd.n3494 0.152939
R14456 gnd.n3497 gnd.n3495 0.152939
R14457 gnd.n3497 gnd.n3496 0.152939
R14458 gnd.n3496 gnd.n2181 0.152939
R14459 gnd.n3530 gnd.n2181 0.152939
R14460 gnd.n3531 gnd.n3530 0.152939
R14461 gnd.n3532 gnd.n3531 0.152939
R14462 gnd.n3532 gnd.n2160 0.152939
R14463 gnd.n3558 gnd.n2160 0.152939
R14464 gnd.n3559 gnd.n3558 0.152939
R14465 gnd.n3561 gnd.n3559 0.152939
R14466 gnd.n3561 gnd.n3560 0.152939
R14467 gnd.n3560 gnd.n2130 0.152939
R14468 gnd.n3596 gnd.n2130 0.152939
R14469 gnd.n3597 gnd.n3596 0.152939
R14470 gnd.n3613 gnd.n3597 0.152939
R14471 gnd.n3613 gnd.n3612 0.152939
R14472 gnd.n3612 gnd.n3611 0.152939
R14473 gnd.n3611 gnd.n3598 0.152939
R14474 gnd.n3607 gnd.n3598 0.152939
R14475 gnd.n3607 gnd.n3606 0.152939
R14476 gnd.n3606 gnd.n3605 0.152939
R14477 gnd.n3605 gnd.n3603 0.152939
R14478 gnd.n3603 gnd.n2080 0.152939
R14479 gnd.n3680 gnd.n2080 0.152939
R14480 gnd.n3681 gnd.n3680 0.152939
R14481 gnd.n3682 gnd.n3681 0.152939
R14482 gnd.n3682 gnd.n2057 0.152939
R14483 gnd.n3731 gnd.n2057 0.152939
R14484 gnd.n3731 gnd.n3730 0.152939
R14485 gnd.n3730 gnd.n3729 0.152939
R14486 gnd.n3729 gnd.n2034 0.152939
R14487 gnd.n3771 gnd.n2034 0.152939
R14488 gnd.n3771 gnd.n3770 0.152939
R14489 gnd.n3770 gnd.n3769 0.152939
R14490 gnd.n3769 gnd.n2012 0.152939
R14491 gnd.n3810 gnd.n2012 0.152939
R14492 gnd.n3810 gnd.n3809 0.152939
R14493 gnd.n3809 gnd.n3808 0.152939
R14494 gnd.n3808 gnd.n1988 0.152939
R14495 gnd.n3858 gnd.n1988 0.152939
R14496 gnd.n3858 gnd.n3857 0.152939
R14497 gnd.n3857 gnd.n3856 0.152939
R14498 gnd.n3856 gnd.n1989 0.152939
R14499 gnd.n1989 gnd.n1783 0.152939
R14500 gnd.n4053 gnd.n1783 0.152939
R14501 gnd.n4054 gnd.n4053 0.152939
R14502 gnd.n4055 gnd.n4054 0.152939
R14503 gnd.n4055 gnd.n1772 0.152939
R14504 gnd.n4074 gnd.n1772 0.152939
R14505 gnd.n4075 gnd.n4074 0.152939
R14506 gnd.n4076 gnd.n4075 0.152939
R14507 gnd.n4076 gnd.n1760 0.152939
R14508 gnd.n4095 gnd.n1760 0.152939
R14509 gnd.n4096 gnd.n4095 0.152939
R14510 gnd.n4098 gnd.n4096 0.152939
R14511 gnd.n4098 gnd.n4097 0.152939
R14512 gnd.n4097 gnd.n1749 0.152939
R14513 gnd.n4119 gnd.n1749 0.152939
R14514 gnd.n3229 gnd.n2497 0.152939
R14515 gnd.n3229 gnd.n3228 0.152939
R14516 gnd.n3228 gnd.n3227 0.152939
R14517 gnd.n3227 gnd.n2504 0.152939
R14518 gnd.n3223 gnd.n2504 0.152939
R14519 gnd.n3223 gnd.n3222 0.152939
R14520 gnd.n3222 gnd.n2511 0.152939
R14521 gnd.n3218 gnd.n2511 0.152939
R14522 gnd.n3218 gnd.n3217 0.152939
R14523 gnd.n2873 gnd.n2632 0.152939
R14524 gnd.n2873 gnd.n2872 0.152939
R14525 gnd.n2872 gnd.n2871 0.152939
R14526 gnd.n2871 gnd.n2595 0.152939
R14527 gnd.n2910 gnd.n2595 0.152939
R14528 gnd.n2911 gnd.n2910 0.152939
R14529 gnd.n2912 gnd.n2911 0.152939
R14530 gnd.n2912 gnd.n2580 0.152939
R14531 gnd.n2957 gnd.n2580 0.152939
R14532 gnd.n2957 gnd.n2956 0.152939
R14533 gnd.n2956 gnd.n2955 0.152939
R14534 gnd.n2955 gnd.n2581 0.152939
R14535 gnd.n2951 gnd.n2581 0.152939
R14536 gnd.n2951 gnd.n2950 0.152939
R14537 gnd.n2950 gnd.n2949 0.152939
R14538 gnd.n2949 gnd.n2585 0.152939
R14539 gnd.n2945 gnd.n2585 0.152939
R14540 gnd.n2945 gnd.n2496 0.152939
R14541 gnd.n3236 gnd.n2496 0.152939
R14542 gnd.n3236 gnd.n3235 0.152939
R14543 gnd.n4502 gnd.n1334 0.152939
R14544 gnd.n4498 gnd.n1334 0.152939
R14545 gnd.n4498 gnd.n4497 0.152939
R14546 gnd.n4497 gnd.n4496 0.152939
R14547 gnd.n4496 gnd.n1339 0.152939
R14548 gnd.n4492 gnd.n1339 0.152939
R14549 gnd.n4492 gnd.n4491 0.152939
R14550 gnd.n4491 gnd.n4490 0.152939
R14551 gnd.n4490 gnd.n1344 0.152939
R14552 gnd.n4486 gnd.n1344 0.152939
R14553 gnd.n4486 gnd.n4485 0.152939
R14554 gnd.n4485 gnd.n4484 0.152939
R14555 gnd.n4484 gnd.n1349 0.152939
R14556 gnd.n4480 gnd.n1349 0.152939
R14557 gnd.n4480 gnd.n4479 0.152939
R14558 gnd.n4479 gnd.n4478 0.152939
R14559 gnd.n4478 gnd.n1354 0.152939
R14560 gnd.n4474 gnd.n1354 0.152939
R14561 gnd.n4474 gnd.n4473 0.152939
R14562 gnd.n4473 gnd.n4472 0.152939
R14563 gnd.n4472 gnd.n1359 0.152939
R14564 gnd.n4468 gnd.n1359 0.152939
R14565 gnd.n4468 gnd.n4467 0.152939
R14566 gnd.n4467 gnd.n4466 0.152939
R14567 gnd.n4466 gnd.n1364 0.152939
R14568 gnd.n4462 gnd.n1364 0.152939
R14569 gnd.n4462 gnd.n4461 0.152939
R14570 gnd.n4461 gnd.n4460 0.152939
R14571 gnd.n4460 gnd.n1369 0.152939
R14572 gnd.n4456 gnd.n1369 0.152939
R14573 gnd.n4456 gnd.n4455 0.152939
R14574 gnd.n4455 gnd.n4454 0.152939
R14575 gnd.n4454 gnd.n1374 0.152939
R14576 gnd.n4450 gnd.n1374 0.152939
R14577 gnd.n4450 gnd.n4449 0.152939
R14578 gnd.n4449 gnd.n4448 0.152939
R14579 gnd.n4448 gnd.n1379 0.152939
R14580 gnd.n4444 gnd.n1379 0.152939
R14581 gnd.n4444 gnd.n4443 0.152939
R14582 gnd.n4443 gnd.n4442 0.152939
R14583 gnd.n4442 gnd.n1384 0.152939
R14584 gnd.n4438 gnd.n1384 0.152939
R14585 gnd.n4438 gnd.n4437 0.152939
R14586 gnd.n4437 gnd.n4436 0.152939
R14587 gnd.n4436 gnd.n1389 0.152939
R14588 gnd.n4432 gnd.n1389 0.152939
R14589 gnd.n4432 gnd.n4431 0.152939
R14590 gnd.n4431 gnd.n4430 0.152939
R14591 gnd.n4430 gnd.n1394 0.152939
R14592 gnd.n4426 gnd.n1394 0.152939
R14593 gnd.n4426 gnd.n4425 0.152939
R14594 gnd.n4425 gnd.n4424 0.152939
R14595 gnd.n4424 gnd.n1399 0.152939
R14596 gnd.n4420 gnd.n1399 0.152939
R14597 gnd.n4420 gnd.n4419 0.152939
R14598 gnd.n4419 gnd.n4418 0.152939
R14599 gnd.n4418 gnd.n1404 0.152939
R14600 gnd.n4414 gnd.n1404 0.152939
R14601 gnd.n4414 gnd.n4413 0.152939
R14602 gnd.n4413 gnd.n4412 0.152939
R14603 gnd.n4412 gnd.n1409 0.152939
R14604 gnd.n4408 gnd.n1409 0.152939
R14605 gnd.n4408 gnd.n4407 0.152939
R14606 gnd.n4407 gnd.n4406 0.152939
R14607 gnd.n4406 gnd.n1414 0.152939
R14608 gnd.n4402 gnd.n1414 0.152939
R14609 gnd.n4402 gnd.n4401 0.152939
R14610 gnd.n4401 gnd.n4400 0.152939
R14611 gnd.n4400 gnd.n1419 0.152939
R14612 gnd.n4396 gnd.n1419 0.152939
R14613 gnd.n4396 gnd.n4395 0.152939
R14614 gnd.n4395 gnd.n4394 0.152939
R14615 gnd.n4394 gnd.n1424 0.152939
R14616 gnd.n4390 gnd.n1424 0.152939
R14617 gnd.n4390 gnd.n4389 0.152939
R14618 gnd.n4389 gnd.n4388 0.152939
R14619 gnd.n4388 gnd.n1429 0.152939
R14620 gnd.n4384 gnd.n1429 0.152939
R14621 gnd.n4384 gnd.n4383 0.152939
R14622 gnd.n4383 gnd.n4382 0.152939
R14623 gnd.n4382 gnd.n1434 0.152939
R14624 gnd.n1437 gnd.n1434 0.152939
R14625 gnd.n1646 gnd.n1479 0.152939
R14626 gnd.n4352 gnd.n1479 0.152939
R14627 gnd.n4352 gnd.n4351 0.152939
R14628 gnd.n4351 gnd.n4350 0.152939
R14629 gnd.n4350 gnd.n1480 0.152939
R14630 gnd.n4346 gnd.n1480 0.152939
R14631 gnd.n4346 gnd.n4345 0.152939
R14632 gnd.n4345 gnd.n4344 0.152939
R14633 gnd.n4344 gnd.n1485 0.152939
R14634 gnd.n4340 gnd.n1485 0.152939
R14635 gnd.n4340 gnd.n4339 0.152939
R14636 gnd.n4339 gnd.n4338 0.152939
R14637 gnd.n4338 gnd.n1490 0.152939
R14638 gnd.n4334 gnd.n1490 0.152939
R14639 gnd.n4334 gnd.n4333 0.152939
R14640 gnd.n4333 gnd.n4332 0.152939
R14641 gnd.n4332 gnd.n241 0.152939
R14642 gnd.n7110 gnd.n241 0.152939
R14643 gnd.n7110 gnd.n7109 0.152939
R14644 gnd.n7109 gnd.n7108 0.152939
R14645 gnd.n7108 gnd.n242 0.152939
R14646 gnd.n7104 gnd.n242 0.152939
R14647 gnd.n7104 gnd.n7103 0.152939
R14648 gnd.n7103 gnd.n7102 0.152939
R14649 gnd.n7102 gnd.n247 0.152939
R14650 gnd.n247 gnd.n217 0.152939
R14651 gnd.n7125 gnd.n217 0.152939
R14652 gnd.n7126 gnd.n7125 0.152939
R14653 gnd.n7127 gnd.n7126 0.152939
R14654 gnd.n7127 gnd.n200 0.152939
R14655 gnd.n7141 gnd.n200 0.152939
R14656 gnd.n7142 gnd.n7141 0.152939
R14657 gnd.n7143 gnd.n7142 0.152939
R14658 gnd.n7143 gnd.n185 0.152939
R14659 gnd.n7157 gnd.n185 0.152939
R14660 gnd.n7158 gnd.n7157 0.152939
R14661 gnd.n7159 gnd.n7158 0.152939
R14662 gnd.n7159 gnd.n166 0.152939
R14663 gnd.n7175 gnd.n166 0.152939
R14664 gnd.n7176 gnd.n7175 0.152939
R14665 gnd.n7244 gnd.n7176 0.152939
R14666 gnd.n7244 gnd.n7243 0.152939
R14667 gnd.n7242 gnd.n7177 0.152939
R14668 gnd.n7238 gnd.n7177 0.152939
R14669 gnd.n7238 gnd.n7237 0.152939
R14670 gnd.n7237 gnd.n7236 0.152939
R14671 gnd.n7236 gnd.n7183 0.152939
R14672 gnd.n7232 gnd.n7183 0.152939
R14673 gnd.n7232 gnd.n7231 0.152939
R14674 gnd.n7231 gnd.n7230 0.152939
R14675 gnd.n7230 gnd.n7191 0.152939
R14676 gnd.n7226 gnd.n7191 0.152939
R14677 gnd.n7226 gnd.n7225 0.152939
R14678 gnd.n7225 gnd.n7224 0.152939
R14679 gnd.n7224 gnd.n7199 0.152939
R14680 gnd.n7220 gnd.n7199 0.152939
R14681 gnd.n7220 gnd.n7219 0.152939
R14682 gnd.n7219 gnd.n7218 0.152939
R14683 gnd.n7218 gnd.n7207 0.152939
R14684 gnd.n7207 gnd.n78 0.152939
R14685 gnd.n4145 gnd.n4144 0.152939
R14686 gnd.n4145 gnd.n1591 0.152939
R14687 gnd.n4179 gnd.n1591 0.152939
R14688 gnd.n4180 gnd.n4179 0.152939
R14689 gnd.n4182 gnd.n4180 0.152939
R14690 gnd.n4182 gnd.n4181 0.152939
R14691 gnd.n4181 gnd.n1552 0.152939
R14692 gnd.n4210 gnd.n1552 0.152939
R14693 gnd.n4211 gnd.n4210 0.152939
R14694 gnd.n4219 gnd.n4211 0.152939
R14695 gnd.n4219 gnd.n4218 0.152939
R14696 gnd.n4218 gnd.n4217 0.152939
R14697 gnd.n4217 gnd.n4212 0.152939
R14698 gnd.n4212 gnd.n1507 0.152939
R14699 gnd.n4323 gnd.n1507 0.152939
R14700 gnd.n4323 gnd.n4322 0.152939
R14701 gnd.n4322 gnd.n4321 0.152939
R14702 gnd.n4321 gnd.n1508 0.152939
R14703 gnd.n4317 gnd.n1508 0.152939
R14704 gnd.n4317 gnd.n51 0.152939
R14705 gnd.n7360 gnd.n51 0.152939
R14706 gnd.n7360 gnd.n7359 0.152939
R14707 gnd.n7359 gnd.n53 0.152939
R14708 gnd.n7355 gnd.n53 0.152939
R14709 gnd.n7355 gnd.n7354 0.152939
R14710 gnd.n7354 gnd.n7353 0.152939
R14711 gnd.n7353 gnd.n58 0.152939
R14712 gnd.n7349 gnd.n58 0.152939
R14713 gnd.n7349 gnd.n7348 0.152939
R14714 gnd.n7348 gnd.n7347 0.152939
R14715 gnd.n7347 gnd.n63 0.152939
R14716 gnd.n7343 gnd.n63 0.152939
R14717 gnd.n7343 gnd.n7342 0.152939
R14718 gnd.n7342 gnd.n7341 0.152939
R14719 gnd.n7341 gnd.n68 0.152939
R14720 gnd.n7337 gnd.n68 0.152939
R14721 gnd.n7337 gnd.n7336 0.152939
R14722 gnd.n7336 gnd.n7335 0.152939
R14723 gnd.n7335 gnd.n73 0.152939
R14724 gnd.n7331 gnd.n73 0.152939
R14725 gnd.n7331 gnd.n7330 0.152939
R14726 gnd.n7330 gnd.n7329 0.152939
R14727 gnd.n4143 gnd.n4142 0.151415
R14728 gnd.n3234 gnd.n2497 0.151415
R14729 gnd.n2851 gnd.n2850 0.145814
R14730 gnd.n2851 gnd.n2632 0.145814
R14731 gnd.n4936 gnd.n0 0.127478
R14732 gnd.n260 gnd.n225 0.10111
R14733 gnd.n2899 gnd.n2898 0.10111
R14734 gnd.n5516 gnd.n5515 0.0767195
R14735 gnd.n5515 gnd.n5514 0.0767195
R14736 gnd.n4504 gnd.n4503 0.063
R14737 gnd.n1647 gnd.n1644 0.063
R14738 gnd.n2900 gnd.n2899 0.0523293
R14739 gnd.n4234 gnd.n225 0.0523293
R14740 gnd.n6020 gnd.n4776 0.0477147
R14741 gnd.n5279 gnd.n5167 0.0442063
R14742 gnd.n5280 gnd.n5279 0.0442063
R14743 gnd.n5281 gnd.n5280 0.0442063
R14744 gnd.n5281 gnd.n5156 0.0442063
R14745 gnd.n5295 gnd.n5156 0.0442063
R14746 gnd.n5296 gnd.n5295 0.0442063
R14747 gnd.n5297 gnd.n5296 0.0442063
R14748 gnd.n5297 gnd.n5143 0.0442063
R14749 gnd.n5341 gnd.n5143 0.0442063
R14750 gnd.n5342 gnd.n5341 0.0442063
R14751 gnd.n5344 gnd.n5077 0.0344674
R14752 gnd.n1731 gnd.n1598 0.0344674
R14753 gnd.n3233 gnd.n2498 0.0344674
R14754 gnd.n5364 gnd.n5363 0.0269946
R14755 gnd.n5366 gnd.n5365 0.0269946
R14756 gnd.n5072 gnd.n5070 0.0269946
R14757 gnd.n5376 gnd.n5374 0.0269946
R14758 gnd.n5375 gnd.n5051 0.0269946
R14759 gnd.n5395 gnd.n5394 0.0269946
R14760 gnd.n5397 gnd.n5396 0.0269946
R14761 gnd.n5046 gnd.n5045 0.0269946
R14762 gnd.n5407 gnd.n5041 0.0269946
R14763 gnd.n5406 gnd.n5043 0.0269946
R14764 gnd.n5042 gnd.n5024 0.0269946
R14765 gnd.n5427 gnd.n5025 0.0269946
R14766 gnd.n5426 gnd.n5026 0.0269946
R14767 gnd.n5460 gnd.n5001 0.0269946
R14768 gnd.n5462 gnd.n5461 0.0269946
R14769 gnd.n5463 gnd.n4948 0.0269946
R14770 gnd.n4996 gnd.n4949 0.0269946
R14771 gnd.n4998 gnd.n4950 0.0269946
R14772 gnd.n5473 gnd.n5472 0.0269946
R14773 gnd.n5475 gnd.n5474 0.0269946
R14774 gnd.n5476 gnd.n4970 0.0269946
R14775 gnd.n5478 gnd.n4971 0.0269946
R14776 gnd.n5481 gnd.n4972 0.0269946
R14777 gnd.n5484 gnd.n5483 0.0269946
R14778 gnd.n5486 gnd.n5485 0.0269946
R14779 gnd.n5551 gnd.n4883 0.0269946
R14780 gnd.n5553 gnd.n5552 0.0269946
R14781 gnd.n5562 gnd.n4876 0.0269946
R14782 gnd.n5564 gnd.n5563 0.0269946
R14783 gnd.n5565 gnd.n4874 0.0269946
R14784 gnd.n5572 gnd.n5568 0.0269946
R14785 gnd.n5571 gnd.n5570 0.0269946
R14786 gnd.n5569 gnd.n4853 0.0269946
R14787 gnd.n5596 gnd.n4854 0.0269946
R14788 gnd.n5595 gnd.n4855 0.0269946
R14789 gnd.n5592 gnd.n936 0.0269946
R14790 gnd.n4831 gnd.n937 0.0269946
R14791 gnd.n4833 gnd.n938 0.0269946
R14792 gnd.n5648 gnd.n5647 0.0269946
R14793 gnd.n5650 gnd.n5649 0.0269946
R14794 gnd.n5651 gnd.n959 0.0269946
R14795 gnd.n5653 gnd.n960 0.0269946
R14796 gnd.n5655 gnd.n961 0.0269946
R14797 gnd.n5661 gnd.n5660 0.0269946
R14798 gnd.n5663 gnd.n5662 0.0269946
R14799 gnd.n5664 gnd.n984 0.0269946
R14800 gnd.n5665 gnd.n985 0.0269946
R14801 gnd.n5666 gnd.n986 0.0269946
R14802 gnd.n5926 gnd.n5925 0.0269946
R14803 gnd.n5927 gnd.n1010 0.0269946
R14804 gnd.n5928 gnd.n1011 0.0269946
R14805 gnd.n5929 gnd.n1012 0.0269946
R14806 gnd.n1644 gnd.n1643 0.0246168
R14807 gnd.n4503 gnd.n1333 0.0246168
R14808 gnd.n5344 gnd.n5343 0.0202011
R14809 gnd.n1643 gnd.n1641 0.0174837
R14810 gnd.n1655 gnd.n1641 0.0174837
R14811 gnd.n1657 gnd.n1655 0.0174837
R14812 gnd.n1657 gnd.n1656 0.0174837
R14813 gnd.n1656 gnd.n1636 0.0174837
R14814 gnd.n1666 gnd.n1636 0.0174837
R14815 gnd.n1666 gnd.n1665 0.0174837
R14816 gnd.n1665 gnd.n1637 0.0174837
R14817 gnd.n1637 gnd.n1632 0.0174837
R14818 gnd.n1674 gnd.n1632 0.0174837
R14819 gnd.n1676 gnd.n1674 0.0174837
R14820 gnd.n1676 gnd.n1675 0.0174837
R14821 gnd.n1675 gnd.n1627 0.0174837
R14822 gnd.n1685 gnd.n1627 0.0174837
R14823 gnd.n1685 gnd.n1684 0.0174837
R14824 gnd.n1684 gnd.n1628 0.0174837
R14825 gnd.n1628 gnd.n1623 0.0174837
R14826 gnd.n1693 gnd.n1623 0.0174837
R14827 gnd.n1695 gnd.n1693 0.0174837
R14828 gnd.n1695 gnd.n1694 0.0174837
R14829 gnd.n1694 gnd.n1618 0.0174837
R14830 gnd.n1704 gnd.n1618 0.0174837
R14831 gnd.n1704 gnd.n1703 0.0174837
R14832 gnd.n1703 gnd.n1619 0.0174837
R14833 gnd.n1619 gnd.n1614 0.0174837
R14834 gnd.n1712 gnd.n1614 0.0174837
R14835 gnd.n1714 gnd.n1712 0.0174837
R14836 gnd.n1714 gnd.n1713 0.0174837
R14837 gnd.n1713 gnd.n1609 0.0174837
R14838 gnd.n1723 gnd.n1609 0.0174837
R14839 gnd.n1723 gnd.n1722 0.0174837
R14840 gnd.n1722 gnd.n1610 0.0174837
R14841 gnd.n1610 gnd.n1603 0.0174837
R14842 gnd.n1730 gnd.n1603 0.0174837
R14843 gnd.n1731 gnd.n1730 0.0174837
R14844 gnd.n3012 gnd.n1333 0.0174837
R14845 gnd.n3014 gnd.n3012 0.0174837
R14846 gnd.n3122 gnd.n3014 0.0174837
R14847 gnd.n3122 gnd.n3121 0.0174837
R14848 gnd.n3121 gnd.n3015 0.0174837
R14849 gnd.n3118 gnd.n3015 0.0174837
R14850 gnd.n3118 gnd.n3117 0.0174837
R14851 gnd.n3117 gnd.n3025 0.0174837
R14852 gnd.n3114 gnd.n3025 0.0174837
R14853 gnd.n3114 gnd.n3113 0.0174837
R14854 gnd.n3113 gnd.n3030 0.0174837
R14855 gnd.n3110 gnd.n3030 0.0174837
R14856 gnd.n3110 gnd.n3109 0.0174837
R14857 gnd.n3109 gnd.n3036 0.0174837
R14858 gnd.n3106 gnd.n3036 0.0174837
R14859 gnd.n3106 gnd.n3105 0.0174837
R14860 gnd.n3105 gnd.n3040 0.0174837
R14861 gnd.n3102 gnd.n3040 0.0174837
R14862 gnd.n3102 gnd.n3101 0.0174837
R14863 gnd.n3101 gnd.n3047 0.0174837
R14864 gnd.n3098 gnd.n3047 0.0174837
R14865 gnd.n3098 gnd.n3097 0.0174837
R14866 gnd.n3097 gnd.n3053 0.0174837
R14867 gnd.n3094 gnd.n3053 0.0174837
R14868 gnd.n3094 gnd.n3093 0.0174837
R14869 gnd.n3093 gnd.n3059 0.0174837
R14870 gnd.n3090 gnd.n3059 0.0174837
R14871 gnd.n3090 gnd.n3089 0.0174837
R14872 gnd.n3089 gnd.n3063 0.0174837
R14873 gnd.n3086 gnd.n3063 0.0174837
R14874 gnd.n3086 gnd.n3085 0.0174837
R14875 gnd.n3085 gnd.n3072 0.0174837
R14876 gnd.n3082 gnd.n3072 0.0174837
R14877 gnd.n3082 gnd.n3081 0.0174837
R14878 gnd.n3081 gnd.n2498 0.0174837
R14879 gnd.n5343 gnd.n5342 0.0148637
R14880 gnd.n5923 gnd.n5667 0.0144266
R14881 gnd.n5924 gnd.n5923 0.0130679
R14882 gnd.n5363 gnd.n5077 0.00797283
R14883 gnd.n5365 gnd.n5364 0.00797283
R14884 gnd.n5366 gnd.n5072 0.00797283
R14885 gnd.n5374 gnd.n5070 0.00797283
R14886 gnd.n5376 gnd.n5375 0.00797283
R14887 gnd.n5394 gnd.n5051 0.00797283
R14888 gnd.n5396 gnd.n5395 0.00797283
R14889 gnd.n5397 gnd.n5046 0.00797283
R14890 gnd.n5045 gnd.n5041 0.00797283
R14891 gnd.n5407 gnd.n5406 0.00797283
R14892 gnd.n5043 gnd.n5042 0.00797283
R14893 gnd.n5025 gnd.n5024 0.00797283
R14894 gnd.n5427 gnd.n5426 0.00797283
R14895 gnd.n5026 gnd.n5001 0.00797283
R14896 gnd.n5461 gnd.n5460 0.00797283
R14897 gnd.n5463 gnd.n5462 0.00797283
R14898 gnd.n4996 gnd.n4948 0.00797283
R14899 gnd.n4998 gnd.n4949 0.00797283
R14900 gnd.n5472 gnd.n4950 0.00797283
R14901 gnd.n5474 gnd.n5473 0.00797283
R14902 gnd.n5476 gnd.n5475 0.00797283
R14903 gnd.n5478 gnd.n4970 0.00797283
R14904 gnd.n5481 gnd.n4971 0.00797283
R14905 gnd.n5483 gnd.n4972 0.00797283
R14906 gnd.n5486 gnd.n5484 0.00797283
R14907 gnd.n5485 gnd.n4883 0.00797283
R14908 gnd.n5553 gnd.n5551 0.00797283
R14909 gnd.n5552 gnd.n4876 0.00797283
R14910 gnd.n5563 gnd.n5562 0.00797283
R14911 gnd.n5565 gnd.n5564 0.00797283
R14912 gnd.n5568 gnd.n4874 0.00797283
R14913 gnd.n5572 gnd.n5571 0.00797283
R14914 gnd.n5570 gnd.n5569 0.00797283
R14915 gnd.n4854 gnd.n4853 0.00797283
R14916 gnd.n5596 gnd.n5595 0.00797283
R14917 gnd.n5592 gnd.n4855 0.00797283
R14918 gnd.n4831 gnd.n936 0.00797283
R14919 gnd.n4833 gnd.n937 0.00797283
R14920 gnd.n5647 gnd.n938 0.00797283
R14921 gnd.n5649 gnd.n5648 0.00797283
R14922 gnd.n5651 gnd.n5650 0.00797283
R14923 gnd.n5653 gnd.n959 0.00797283
R14924 gnd.n5655 gnd.n960 0.00797283
R14925 gnd.n5660 gnd.n961 0.00797283
R14926 gnd.n5662 gnd.n5661 0.00797283
R14927 gnd.n5664 gnd.n5663 0.00797283
R14928 gnd.n5665 gnd.n984 0.00797283
R14929 gnd.n5666 gnd.n985 0.00797283
R14930 gnd.n5667 gnd.n986 0.00797283
R14931 gnd.n5925 gnd.n5924 0.00797283
R14932 gnd.n5927 gnd.n5926 0.00797283
R14933 gnd.n5928 gnd.n1010 0.00797283
R14934 gnd.n5929 gnd.n1011 0.00797283
R14935 gnd.n4776 gnd.n1012 0.00797283
R14936 gnd.n4275 gnd.n242 0.00614909
R14937 gnd.n2849 gnd.n2636 0.00614909
R14938 gnd.n4143 gnd.n1598 0.000839674
R14939 gnd.n3234 gnd.n3233 0.000839674
R14940 a_n2982_13878.n14 a_n2982_13878.t102 538.698
R14941 a_n2982_13878.n141 a_n2982_13878.t79 512.366
R14942 a_n2982_13878.n140 a_n2982_13878.t84 512.366
R14943 a_n2982_13878.n93 a_n2982_13878.t72 512.366
R14944 a_n2982_13878.n139 a_n2982_13878.t89 512.366
R14945 a_n2982_13878.n138 a_n2982_13878.t98 512.366
R14946 a_n2982_13878.n94 a_n2982_13878.t99 512.366
R14947 a_n2982_13878.n137 a_n2982_13878.t66 512.366
R14948 a_n2982_13878.n136 a_n2982_13878.t81 512.366
R14949 a_n2982_13878.n95 a_n2982_13878.t69 512.366
R14950 a_n2982_13878.n135 a_n2982_13878.t76 512.366
R14951 a_n2982_13878.n8 a_n2982_13878.t35 538.698
R14952 a_n2982_13878.n148 a_n2982_13878.t59 512.366
R14953 a_n2982_13878.n147 a_n2982_13878.t17 512.366
R14954 a_n2982_13878.n82 a_n2982_13878.t45 512.366
R14955 a_n2982_13878.n146 a_n2982_13878.t61 512.366
R14956 a_n2982_13878.n145 a_n2982_13878.t43 512.366
R14957 a_n2982_13878.n83 a_n2982_13878.t27 512.366
R14958 a_n2982_13878.n144 a_n2982_13878.t37 512.366
R14959 a_n2982_13878.n143 a_n2982_13878.t15 512.366
R14960 a_n2982_13878.n84 a_n2982_13878.t29 512.366
R14961 a_n2982_13878.n142 a_n2982_13878.t53 512.366
R14962 a_n2982_13878.n29 a_n2982_13878.t57 538.698
R14963 a_n2982_13878.n115 a_n2982_13878.t21 512.366
R14964 a_n2982_13878.n104 a_n2982_13878.t39 512.366
R14965 a_n2982_13878.n116 a_n2982_13878.t51 512.366
R14966 a_n2982_13878.n103 a_n2982_13878.t25 512.366
R14967 a_n2982_13878.n117 a_n2982_13878.t19 512.366
R14968 a_n2982_13878.n118 a_n2982_13878.t47 512.366
R14969 a_n2982_13878.n102 a_n2982_13878.t49 512.366
R14970 a_n2982_13878.n119 a_n2982_13878.t23 512.366
R14971 a_n2982_13878.n101 a_n2982_13878.t31 512.366
R14972 a_n2982_13878.n120 a_n2982_13878.t33 512.366
R14973 a_n2982_13878.n35 a_n2982_13878.t101 538.698
R14974 a_n2982_13878.n109 a_n2982_13878.t70 512.366
R14975 a_n2982_13878.n108 a_n2982_13878.t71 512.366
R14976 a_n2982_13878.n110 a_n2982_13878.t96 512.366
R14977 a_n2982_13878.n107 a_n2982_13878.t97 512.366
R14978 a_n2982_13878.n111 a_n2982_13878.t68 512.366
R14979 a_n2982_13878.n112 a_n2982_13878.t92 512.366
R14980 a_n2982_13878.n106 a_n2982_13878.t93 512.366
R14981 a_n2982_13878.n113 a_n2982_13878.t65 512.366
R14982 a_n2982_13878.n105 a_n2982_13878.t78 512.366
R14983 a_n2982_13878.n114 a_n2982_13878.t88 512.366
R14984 a_n2982_13878.n132 a_n2982_13878.t86 512.366
R14985 a_n2982_13878.n122 a_n2982_13878.t75 512.366
R14986 a_n2982_13878.n133 a_n2982_13878.t64 512.366
R14987 a_n2982_13878.n130 a_n2982_13878.t94 512.366
R14988 a_n2982_13878.n123 a_n2982_13878.t83 512.366
R14989 a_n2982_13878.n131 a_n2982_13878.t82 512.366
R14990 a_n2982_13878.n128 a_n2982_13878.t90 512.366
R14991 a_n2982_13878.n124 a_n2982_13878.t73 512.366
R14992 a_n2982_13878.n129 a_n2982_13878.t74 512.366
R14993 a_n2982_13878.n126 a_n2982_13878.t77 512.366
R14994 a_n2982_13878.n125 a_n2982_13878.t87 512.366
R14995 a_n2982_13878.n127 a_n2982_13878.t103 512.366
R14996 a_n2982_13878.n73 a_n2982_13878.n9 70.5844
R14997 a_n2982_13878.n81 a_n2982_13878.n3 70.5844
R14998 a_n2982_13878.n25 a_n2982_13878.n57 70.5844
R14999 a_n2982_13878.n31 a_n2982_13878.n49 70.5844
R15000 a_n2982_13878.n48 a_n2982_13878.n31 70.1674
R15001 a_n2982_13878.n48 a_n2982_13878.n105 20.9683
R15002 a_n2982_13878.n30 a_n2982_13878.n47 74.73
R15003 a_n2982_13878.n113 a_n2982_13878.n47 11.843
R15004 a_n2982_13878.n46 a_n2982_13878.n30 80.4688
R15005 a_n2982_13878.n46 a_n2982_13878.n106 0.365327
R15006 a_n2982_13878.n32 a_n2982_13878.n45 75.0448
R15007 a_n2982_13878.n44 a_n2982_13878.n32 70.1674
R15008 a_n2982_13878.n44 a_n2982_13878.n107 20.9683
R15009 a_n2982_13878.n33 a_n2982_13878.n43 70.3058
R15010 a_n2982_13878.n110 a_n2982_13878.n43 20.6913
R15011 a_n2982_13878.n42 a_n2982_13878.n33 75.3623
R15012 a_n2982_13878.n42 a_n2982_13878.n108 10.5784
R15013 a_n2982_13878.n35 a_n2982_13878.n34 44.7878
R15014 a_n2982_13878.n56 a_n2982_13878.n25 70.1674
R15015 a_n2982_13878.n56 a_n2982_13878.n101 20.9683
R15016 a_n2982_13878.n24 a_n2982_13878.n55 74.73
R15017 a_n2982_13878.n119 a_n2982_13878.n55 11.843
R15018 a_n2982_13878.n54 a_n2982_13878.n24 80.4688
R15019 a_n2982_13878.n54 a_n2982_13878.n102 0.365327
R15020 a_n2982_13878.n26 a_n2982_13878.n53 75.0448
R15021 a_n2982_13878.n52 a_n2982_13878.n26 70.1674
R15022 a_n2982_13878.n52 a_n2982_13878.n103 20.9683
R15023 a_n2982_13878.n27 a_n2982_13878.n51 70.3058
R15024 a_n2982_13878.n116 a_n2982_13878.n51 20.6913
R15025 a_n2982_13878.n50 a_n2982_13878.n27 75.3623
R15026 a_n2982_13878.n50 a_n2982_13878.n104 10.5784
R15027 a_n2982_13878.n29 a_n2982_13878.n28 44.7878
R15028 a_n2982_13878.n15 a_n2982_13878.n65 70.1674
R15029 a_n2982_13878.n17 a_n2982_13878.n63 70.1674
R15030 a_n2982_13878.n19 a_n2982_13878.n61 70.1674
R15031 a_n2982_13878.n22 a_n2982_13878.n59 70.1674
R15032 a_n2982_13878.n127 a_n2982_13878.n59 20.9683
R15033 a_n2982_13878.n58 a_n2982_13878.n23 75.0448
R15034 a_n2982_13878.n58 a_n2982_13878.n125 11.2134
R15035 a_n2982_13878.n23 a_n2982_13878.n126 161.3
R15036 a_n2982_13878.n129 a_n2982_13878.n61 20.9683
R15037 a_n2982_13878.n60 a_n2982_13878.n20 75.0448
R15038 a_n2982_13878.n60 a_n2982_13878.n124 11.2134
R15039 a_n2982_13878.n20 a_n2982_13878.n128 161.3
R15040 a_n2982_13878.n131 a_n2982_13878.n63 20.9683
R15041 a_n2982_13878.n62 a_n2982_13878.n18 75.0448
R15042 a_n2982_13878.n62 a_n2982_13878.n123 11.2134
R15043 a_n2982_13878.n18 a_n2982_13878.n130 161.3
R15044 a_n2982_13878.n133 a_n2982_13878.n65 20.9683
R15045 a_n2982_13878.n64 a_n2982_13878.n16 75.0448
R15046 a_n2982_13878.n64 a_n2982_13878.n122 11.2134
R15047 a_n2982_13878.n16 a_n2982_13878.n132 161.3
R15048 a_n2982_13878.n9 a_n2982_13878.n72 70.1674
R15049 a_n2982_13878.n72 a_n2982_13878.n95 20.9683
R15050 a_n2982_13878.n71 a_n2982_13878.n10 74.73
R15051 a_n2982_13878.n136 a_n2982_13878.n71 11.843
R15052 a_n2982_13878.n70 a_n2982_13878.n10 80.4688
R15053 a_n2982_13878.n70 a_n2982_13878.n137 0.365327
R15054 a_n2982_13878.n11 a_n2982_13878.n69 75.0448
R15055 a_n2982_13878.n68 a_n2982_13878.n11 70.1674
R15056 a_n2982_13878.n139 a_n2982_13878.n68 20.9683
R15057 a_n2982_13878.n13 a_n2982_13878.n67 70.3058
R15058 a_n2982_13878.n67 a_n2982_13878.n93 20.6913
R15059 a_n2982_13878.n66 a_n2982_13878.n13 75.3623
R15060 a_n2982_13878.n140 a_n2982_13878.n66 10.5784
R15061 a_n2982_13878.n12 a_n2982_13878.n14 44.7878
R15062 a_n2982_13878.n3 a_n2982_13878.n80 70.1674
R15063 a_n2982_13878.n80 a_n2982_13878.n84 20.9683
R15064 a_n2982_13878.n79 a_n2982_13878.n4 74.73
R15065 a_n2982_13878.n143 a_n2982_13878.n79 11.843
R15066 a_n2982_13878.n78 a_n2982_13878.n4 80.4688
R15067 a_n2982_13878.n78 a_n2982_13878.n144 0.365327
R15068 a_n2982_13878.n5 a_n2982_13878.n77 75.0448
R15069 a_n2982_13878.n76 a_n2982_13878.n5 70.1674
R15070 a_n2982_13878.n146 a_n2982_13878.n76 20.9683
R15071 a_n2982_13878.n7 a_n2982_13878.n75 70.3058
R15072 a_n2982_13878.n75 a_n2982_13878.n82 20.6913
R15073 a_n2982_13878.n74 a_n2982_13878.n7 75.3623
R15074 a_n2982_13878.n147 a_n2982_13878.n74 10.5784
R15075 a_n2982_13878.n6 a_n2982_13878.n8 44.7878
R15076 a_n2982_13878.n1 a_n2982_13878.n91 81.4626
R15077 a_n2982_13878.n2 a_n2982_13878.n87 81.4626
R15078 a_n2982_13878.n2 a_n2982_13878.n85 81.4626
R15079 a_n2982_13878.n1 a_n2982_13878.n92 80.9324
R15080 a_n2982_13878.n1 a_n2982_13878.n90 80.9324
R15081 a_n2982_13878.n0 a_n2982_13878.n89 80.9324
R15082 a_n2982_13878.n2 a_n2982_13878.n88 80.9324
R15083 a_n2982_13878.n2 a_n2982_13878.n86 80.9324
R15084 a_n2982_13878.n41 a_n2982_13878.t42 74.6477
R15085 a_n2982_13878.n36 a_n2982_13878.t58 74.6477
R15086 a_n2982_13878.n39 a_n2982_13878.t36 74.2899
R15087 a_n2982_13878.n38 a_n2982_13878.t56 74.2897
R15088 a_n2982_13878.n41 a_n2982_13878.n153 70.6783
R15089 a_n2982_13878.n40 a_n2982_13878.n152 70.6783
R15090 a_n2982_13878.n40 a_n2982_13878.n151 70.6783
R15091 a_n2982_13878.n39 a_n2982_13878.n150 70.6783
R15092 a_n2982_13878.n38 a_n2982_13878.n100 70.6783
R15093 a_n2982_13878.n37 a_n2982_13878.n99 70.6783
R15094 a_n2982_13878.n37 a_n2982_13878.n98 70.6783
R15095 a_n2982_13878.n36 a_n2982_13878.n97 70.6783
R15096 a_n2982_13878.n36 a_n2982_13878.n96 70.6783
R15097 a_n2982_13878.n154 a_n2982_13878.n41 70.6782
R15098 a_n2982_13878.n141 a_n2982_13878.n140 48.2005
R15099 a_n2982_13878.n68 a_n2982_13878.n138 20.9683
R15100 a_n2982_13878.n137 a_n2982_13878.n94 48.2005
R15101 a_n2982_13878.n135 a_n2982_13878.n72 20.9683
R15102 a_n2982_13878.n148 a_n2982_13878.n147 48.2005
R15103 a_n2982_13878.n76 a_n2982_13878.n145 20.9683
R15104 a_n2982_13878.n144 a_n2982_13878.n83 48.2005
R15105 a_n2982_13878.n142 a_n2982_13878.n80 20.9683
R15106 a_n2982_13878.n115 a_n2982_13878.n104 48.2005
R15107 a_n2982_13878.n117 a_n2982_13878.n52 20.9683
R15108 a_n2982_13878.n118 a_n2982_13878.n102 48.2005
R15109 a_n2982_13878.n120 a_n2982_13878.n56 20.9683
R15110 a_n2982_13878.n109 a_n2982_13878.n108 48.2005
R15111 a_n2982_13878.n111 a_n2982_13878.n44 20.9683
R15112 a_n2982_13878.n112 a_n2982_13878.n106 48.2005
R15113 a_n2982_13878.n114 a_n2982_13878.n48 20.9683
R15114 a_n2982_13878.n132 a_n2982_13878.n122 48.2005
R15115 a_n2982_13878.t91 a_n2982_13878.n65 533.335
R15116 a_n2982_13878.n130 a_n2982_13878.n123 48.2005
R15117 a_n2982_13878.t100 a_n2982_13878.n63 533.335
R15118 a_n2982_13878.n128 a_n2982_13878.n124 48.2005
R15119 a_n2982_13878.t85 a_n2982_13878.n61 533.335
R15120 a_n2982_13878.n126 a_n2982_13878.n125 48.2005
R15121 a_n2982_13878.t80 a_n2982_13878.n59 533.335
R15122 a_n2982_13878.n139 a_n2982_13878.n67 21.4216
R15123 a_n2982_13878.n146 a_n2982_13878.n75 21.4216
R15124 a_n2982_13878.n103 a_n2982_13878.n51 21.4216
R15125 a_n2982_13878.n107 a_n2982_13878.n43 21.4216
R15126 a_n2982_13878.n73 a_n2982_13878.t95 532.5
R15127 a_n2982_13878.n81 a_n2982_13878.t41 532.5
R15128 a_n2982_13878.t55 a_n2982_13878.n57 532.5
R15129 a_n2982_13878.t67 a_n2982_13878.n49 532.5
R15130 a_n2982_13878.n71 a_n2982_13878.n95 34.4824
R15131 a_n2982_13878.n79 a_n2982_13878.n84 34.4824
R15132 a_n2982_13878.n101 a_n2982_13878.n55 34.4824
R15133 a_n2982_13878.n105 a_n2982_13878.n47 34.4824
R15134 a_n2982_13878.n138 a_n2982_13878.n69 35.3134
R15135 a_n2982_13878.n69 a_n2982_13878.n94 11.2134
R15136 a_n2982_13878.n145 a_n2982_13878.n77 35.3134
R15137 a_n2982_13878.n77 a_n2982_13878.n83 11.2134
R15138 a_n2982_13878.n53 a_n2982_13878.n117 35.3134
R15139 a_n2982_13878.n118 a_n2982_13878.n53 11.2134
R15140 a_n2982_13878.n45 a_n2982_13878.n111 35.3134
R15141 a_n2982_13878.n112 a_n2982_13878.n45 11.2134
R15142 a_n2982_13878.n133 a_n2982_13878.n64 35.3134
R15143 a_n2982_13878.n131 a_n2982_13878.n62 35.3134
R15144 a_n2982_13878.n129 a_n2982_13878.n60 35.3134
R15145 a_n2982_13878.n127 a_n2982_13878.n58 35.3134
R15146 a_n2982_13878.n3 a_n2982_13878.n1 23.891
R15147 a_n2982_13878.n66 a_n2982_13878.n93 36.139
R15148 a_n2982_13878.n74 a_n2982_13878.n82 36.139
R15149 a_n2982_13878.n116 a_n2982_13878.n50 36.139
R15150 a_n2982_13878.n110 a_n2982_13878.n42 36.139
R15151 a_n2982_13878.n34 a_n2982_13878.n21 13.9285
R15152 a_n2982_13878.n9 a_n2982_13878.n134 13.724
R15153 a_n2982_13878.n149 a_n2982_13878.n6 12.4191
R15154 a_n2982_13878.n23 a_n2982_13878.n21 11.2486
R15155 a_n2982_13878.n134 a_n2982_13878.n15 11.2486
R15156 a_n2982_13878.n121 a_n2982_13878.n38 10.5745
R15157 a_n2982_13878.n121 a_n2982_13878.n25 8.58383
R15158 a_n2982_13878.n39 a_n2982_13878.n149 6.7311
R15159 a_n2982_13878.n134 a_n2982_13878.n121 5.3452
R15160 a_n2982_13878.n28 a_n2982_13878.n31 3.94368
R15161 a_n2982_13878.n3 a_n2982_13878.n12 3.94368
R15162 a_n2982_13878.n153 a_n2982_13878.t30 3.61217
R15163 a_n2982_13878.n153 a_n2982_13878.t54 3.61217
R15164 a_n2982_13878.n152 a_n2982_13878.t44 3.61217
R15165 a_n2982_13878.n152 a_n2982_13878.t28 3.61217
R15166 a_n2982_13878.n151 a_n2982_13878.t46 3.61217
R15167 a_n2982_13878.n151 a_n2982_13878.t62 3.61217
R15168 a_n2982_13878.n150 a_n2982_13878.t60 3.61217
R15169 a_n2982_13878.n150 a_n2982_13878.t18 3.61217
R15170 a_n2982_13878.n100 a_n2982_13878.t32 3.61217
R15171 a_n2982_13878.n100 a_n2982_13878.t34 3.61217
R15172 a_n2982_13878.n99 a_n2982_13878.t50 3.61217
R15173 a_n2982_13878.n99 a_n2982_13878.t24 3.61217
R15174 a_n2982_13878.n98 a_n2982_13878.t20 3.61217
R15175 a_n2982_13878.n98 a_n2982_13878.t48 3.61217
R15176 a_n2982_13878.n97 a_n2982_13878.t52 3.61217
R15177 a_n2982_13878.n97 a_n2982_13878.t26 3.61217
R15178 a_n2982_13878.n96 a_n2982_13878.t22 3.61217
R15179 a_n2982_13878.n96 a_n2982_13878.t40 3.61217
R15180 a_n2982_13878.n154 a_n2982_13878.t38 3.61217
R15181 a_n2982_13878.t16 a_n2982_13878.n154 3.61217
R15182 a_n2982_13878.n91 a_n2982_13878.t3 2.82907
R15183 a_n2982_13878.n91 a_n2982_13878.t4 2.82907
R15184 a_n2982_13878.n92 a_n2982_13878.t12 2.82907
R15185 a_n2982_13878.n92 a_n2982_13878.t6 2.82907
R15186 a_n2982_13878.n90 a_n2982_13878.t10 2.82907
R15187 a_n2982_13878.n90 a_n2982_13878.t11 2.82907
R15188 a_n2982_13878.n89 a_n2982_13878.t0 2.82907
R15189 a_n2982_13878.n89 a_n2982_13878.t1 2.82907
R15190 a_n2982_13878.n87 a_n2982_13878.t9 2.82907
R15191 a_n2982_13878.n87 a_n2982_13878.t63 2.82907
R15192 a_n2982_13878.n88 a_n2982_13878.t13 2.82907
R15193 a_n2982_13878.n88 a_n2982_13878.t14 2.82907
R15194 a_n2982_13878.n86 a_n2982_13878.t5 2.82907
R15195 a_n2982_13878.n86 a_n2982_13878.t7 2.82907
R15196 a_n2982_13878.n85 a_n2982_13878.t2 2.82907
R15197 a_n2982_13878.n85 a_n2982_13878.t8 2.82907
R15198 a_n2982_13878.n14 a_n2982_13878.n141 14.1668
R15199 a_n2982_13878.n135 a_n2982_13878.n73 22.3251
R15200 a_n2982_13878.n8 a_n2982_13878.n148 14.1668
R15201 a_n2982_13878.n142 a_n2982_13878.n81 22.3251
R15202 a_n2982_13878.n115 a_n2982_13878.n29 14.1668
R15203 a_n2982_13878.n57 a_n2982_13878.n120 22.3251
R15204 a_n2982_13878.n109 a_n2982_13878.n35 14.1668
R15205 a_n2982_13878.n49 a_n2982_13878.n114 22.3251
R15206 a_n2982_13878.n149 a_n2982_13878.n21 1.30542
R15207 a_n2982_13878.n18 a_n2982_13878.n19 1.04595
R15208 a_n2982_13878.n70 a_n2982_13878.n136 47.835
R15209 a_n2982_13878.n78 a_n2982_13878.n143 47.835
R15210 a_n2982_13878.n119 a_n2982_13878.n54 47.835
R15211 a_n2982_13878.n113 a_n2982_13878.n46 47.835
R15212 a_n2982_13878.n0 a_n2982_13878.n2 32.5247
R15213 a_n2982_13878.n31 a_n2982_13878.n30 1.13686
R15214 a_n2982_13878.n25 a_n2982_13878.n24 1.13686
R15215 a_n2982_13878.n10 a_n2982_13878.n9 1.13686
R15216 a_n2982_13878.n4 a_n2982_13878.n3 1.09898
R15217 a_n2982_13878.n40 a_n2982_13878.n39 1.07378
R15218 a_n2982_13878.n37 a_n2982_13878.n36 1.07378
R15219 a_n2982_13878.n1 a_n2982_13878.n0 1.06084
R15220 a_n2982_13878.n33 a_n2982_13878.n34 0.758076
R15221 a_n2982_13878.n32 a_n2982_13878.n33 0.758076
R15222 a_n2982_13878.n30 a_n2982_13878.n32 0.758076
R15223 a_n2982_13878.n27 a_n2982_13878.n28 0.758076
R15224 a_n2982_13878.n26 a_n2982_13878.n27 0.758076
R15225 a_n2982_13878.n24 a_n2982_13878.n26 0.758076
R15226 a_n2982_13878.n23 a_n2982_13878.n22 0.758076
R15227 a_n2982_13878.n20 a_n2982_13878.n19 0.758076
R15228 a_n2982_13878.n18 a_n2982_13878.n17 0.758076
R15229 a_n2982_13878.n16 a_n2982_13878.n15 0.758076
R15230 a_n2982_13878.n13 a_n2982_13878.n12 0.758076
R15231 a_n2982_13878.n13 a_n2982_13878.n11 0.758076
R15232 a_n2982_13878.n11 a_n2982_13878.n10 0.758076
R15233 a_n2982_13878.n7 a_n2982_13878.n6 0.758076
R15234 a_n2982_13878.n7 a_n2982_13878.n5 0.758076
R15235 a_n2982_13878.n5 a_n2982_13878.n4 0.758076
R15236 a_n2982_13878.n41 a_n2982_13878.n40 0.716017
R15237 a_n2982_13878.n38 a_n2982_13878.n37 0.716017
R15238 a_n2982_13878.n20 a_n2982_13878.n22 0.67853
R15239 a_n2982_13878.n16 a_n2982_13878.n17 0.67853
R15240 vdd.n327 vdd.n291 756.745
R15241 vdd.n268 vdd.n232 756.745
R15242 vdd.n225 vdd.n189 756.745
R15243 vdd.n166 vdd.n130 756.745
R15244 vdd.n124 vdd.n88 756.745
R15245 vdd.n65 vdd.n29 756.745
R15246 vdd.n2201 vdd.n2165 756.745
R15247 vdd.n2260 vdd.n2224 756.745
R15248 vdd.n2099 vdd.n2063 756.745
R15249 vdd.n2158 vdd.n2122 756.745
R15250 vdd.n1998 vdd.n1962 756.745
R15251 vdd.n2057 vdd.n2021 756.745
R15252 vdd.n1315 vdd.t87 640.208
R15253 vdd.n1010 vdd.t128 640.208
R15254 vdd.n1319 vdd.t125 640.208
R15255 vdd.n1001 vdd.t150 640.208
R15256 vdd.n896 vdd.t112 640.208
R15257 vdd.n2823 vdd.t143 640.208
R15258 vdd.n832 vdd.t105 640.208
R15259 vdd.n2820 vdd.t135 640.208
R15260 vdd.n799 vdd.t83 640.208
R15261 vdd.n1071 vdd.t139 640.208
R15262 vdd.n1772 vdd.t153 592.009
R15263 vdd.n1810 vdd.t146 592.009
R15264 vdd.n1706 vdd.t156 592.009
R15265 vdd.n2362 vdd.t116 592.009
R15266 vdd.n1248 vdd.t91 592.009
R15267 vdd.n1208 vdd.t99 592.009
R15268 vdd.n426 vdd.t122 592.009
R15269 vdd.n440 vdd.t95 592.009
R15270 vdd.n452 vdd.t102 592.009
R15271 vdd.n768 vdd.t119 592.009
R15272 vdd.n3456 vdd.t132 592.009
R15273 vdd.n688 vdd.t108 592.009
R15274 vdd.n328 vdd.n327 585
R15275 vdd.n326 vdd.n293 585
R15276 vdd.n325 vdd.n324 585
R15277 vdd.n296 vdd.n294 585
R15278 vdd.n319 vdd.n318 585
R15279 vdd.n317 vdd.n316 585
R15280 vdd.n300 vdd.n299 585
R15281 vdd.n311 vdd.n310 585
R15282 vdd.n309 vdd.n308 585
R15283 vdd.n304 vdd.n303 585
R15284 vdd.n269 vdd.n268 585
R15285 vdd.n267 vdd.n234 585
R15286 vdd.n266 vdd.n265 585
R15287 vdd.n237 vdd.n235 585
R15288 vdd.n260 vdd.n259 585
R15289 vdd.n258 vdd.n257 585
R15290 vdd.n241 vdd.n240 585
R15291 vdd.n252 vdd.n251 585
R15292 vdd.n250 vdd.n249 585
R15293 vdd.n245 vdd.n244 585
R15294 vdd.n226 vdd.n225 585
R15295 vdd.n224 vdd.n191 585
R15296 vdd.n223 vdd.n222 585
R15297 vdd.n194 vdd.n192 585
R15298 vdd.n217 vdd.n216 585
R15299 vdd.n215 vdd.n214 585
R15300 vdd.n198 vdd.n197 585
R15301 vdd.n209 vdd.n208 585
R15302 vdd.n207 vdd.n206 585
R15303 vdd.n202 vdd.n201 585
R15304 vdd.n167 vdd.n166 585
R15305 vdd.n165 vdd.n132 585
R15306 vdd.n164 vdd.n163 585
R15307 vdd.n135 vdd.n133 585
R15308 vdd.n158 vdd.n157 585
R15309 vdd.n156 vdd.n155 585
R15310 vdd.n139 vdd.n138 585
R15311 vdd.n150 vdd.n149 585
R15312 vdd.n148 vdd.n147 585
R15313 vdd.n143 vdd.n142 585
R15314 vdd.n125 vdd.n124 585
R15315 vdd.n123 vdd.n90 585
R15316 vdd.n122 vdd.n121 585
R15317 vdd.n93 vdd.n91 585
R15318 vdd.n116 vdd.n115 585
R15319 vdd.n114 vdd.n113 585
R15320 vdd.n97 vdd.n96 585
R15321 vdd.n108 vdd.n107 585
R15322 vdd.n106 vdd.n105 585
R15323 vdd.n101 vdd.n100 585
R15324 vdd.n66 vdd.n65 585
R15325 vdd.n64 vdd.n31 585
R15326 vdd.n63 vdd.n62 585
R15327 vdd.n34 vdd.n32 585
R15328 vdd.n57 vdd.n56 585
R15329 vdd.n55 vdd.n54 585
R15330 vdd.n38 vdd.n37 585
R15331 vdd.n49 vdd.n48 585
R15332 vdd.n47 vdd.n46 585
R15333 vdd.n42 vdd.n41 585
R15334 vdd.n2202 vdd.n2201 585
R15335 vdd.n2200 vdd.n2167 585
R15336 vdd.n2199 vdd.n2198 585
R15337 vdd.n2170 vdd.n2168 585
R15338 vdd.n2193 vdd.n2192 585
R15339 vdd.n2191 vdd.n2190 585
R15340 vdd.n2174 vdd.n2173 585
R15341 vdd.n2185 vdd.n2184 585
R15342 vdd.n2183 vdd.n2182 585
R15343 vdd.n2178 vdd.n2177 585
R15344 vdd.n2261 vdd.n2260 585
R15345 vdd.n2259 vdd.n2226 585
R15346 vdd.n2258 vdd.n2257 585
R15347 vdd.n2229 vdd.n2227 585
R15348 vdd.n2252 vdd.n2251 585
R15349 vdd.n2250 vdd.n2249 585
R15350 vdd.n2233 vdd.n2232 585
R15351 vdd.n2244 vdd.n2243 585
R15352 vdd.n2242 vdd.n2241 585
R15353 vdd.n2237 vdd.n2236 585
R15354 vdd.n2100 vdd.n2099 585
R15355 vdd.n2098 vdd.n2065 585
R15356 vdd.n2097 vdd.n2096 585
R15357 vdd.n2068 vdd.n2066 585
R15358 vdd.n2091 vdd.n2090 585
R15359 vdd.n2089 vdd.n2088 585
R15360 vdd.n2072 vdd.n2071 585
R15361 vdd.n2083 vdd.n2082 585
R15362 vdd.n2081 vdd.n2080 585
R15363 vdd.n2076 vdd.n2075 585
R15364 vdd.n2159 vdd.n2158 585
R15365 vdd.n2157 vdd.n2124 585
R15366 vdd.n2156 vdd.n2155 585
R15367 vdd.n2127 vdd.n2125 585
R15368 vdd.n2150 vdd.n2149 585
R15369 vdd.n2148 vdd.n2147 585
R15370 vdd.n2131 vdd.n2130 585
R15371 vdd.n2142 vdd.n2141 585
R15372 vdd.n2140 vdd.n2139 585
R15373 vdd.n2135 vdd.n2134 585
R15374 vdd.n1999 vdd.n1998 585
R15375 vdd.n1997 vdd.n1964 585
R15376 vdd.n1996 vdd.n1995 585
R15377 vdd.n1967 vdd.n1965 585
R15378 vdd.n1990 vdd.n1989 585
R15379 vdd.n1988 vdd.n1987 585
R15380 vdd.n1971 vdd.n1970 585
R15381 vdd.n1982 vdd.n1981 585
R15382 vdd.n1980 vdd.n1979 585
R15383 vdd.n1975 vdd.n1974 585
R15384 vdd.n2058 vdd.n2057 585
R15385 vdd.n2056 vdd.n2023 585
R15386 vdd.n2055 vdd.n2054 585
R15387 vdd.n2026 vdd.n2024 585
R15388 vdd.n2049 vdd.n2048 585
R15389 vdd.n2047 vdd.n2046 585
R15390 vdd.n2030 vdd.n2029 585
R15391 vdd.n2041 vdd.n2040 585
R15392 vdd.n2039 vdd.n2038 585
R15393 vdd.n2034 vdd.n2033 585
R15394 vdd.n3628 vdd.n392 509.269
R15395 vdd.n3624 vdd.n393 509.269
R15396 vdd.n3496 vdd.n685 509.269
R15397 vdd.n3493 vdd.n684 509.269
R15398 vdd.n2357 vdd.n1530 509.269
R15399 vdd.n2360 vdd.n2359 509.269
R15400 vdd.n1679 vdd.n1643 509.269
R15401 vdd.n1875 vdd.n1644 509.269
R15402 vdd.n305 vdd.t210 329.043
R15403 vdd.n246 vdd.t65 329.043
R15404 vdd.n203 vdd.t185 329.043
R15405 vdd.n144 vdd.t81 329.043
R15406 vdd.n102 vdd.t202 329.043
R15407 vdd.n43 vdd.t32 329.043
R15408 vdd.n2179 vdd.t211 329.043
R15409 vdd.n2238 vdd.t38 329.043
R15410 vdd.n2077 vdd.t165 329.043
R15411 vdd.n2136 vdd.t60 329.043
R15412 vdd.n1976 vdd.t48 329.043
R15413 vdd.n2035 vdd.t225 329.043
R15414 vdd.n1772 vdd.t155 319.788
R15415 vdd.n1810 vdd.t149 319.788
R15416 vdd.n1706 vdd.t158 319.788
R15417 vdd.n2362 vdd.t117 319.788
R15418 vdd.n1248 vdd.t93 319.788
R15419 vdd.n1208 vdd.t100 319.788
R15420 vdd.n426 vdd.t123 319.788
R15421 vdd.n440 vdd.t97 319.788
R15422 vdd.n452 vdd.t103 319.788
R15423 vdd.n768 vdd.t121 319.788
R15424 vdd.n3456 vdd.t134 319.788
R15425 vdd.n688 vdd.t111 319.788
R15426 vdd.n1773 vdd.t154 303.69
R15427 vdd.n1811 vdd.t148 303.69
R15428 vdd.n1707 vdd.t157 303.69
R15429 vdd.n2363 vdd.t118 303.69
R15430 vdd.n1249 vdd.t94 303.69
R15431 vdd.n1209 vdd.t101 303.69
R15432 vdd.n427 vdd.t124 303.69
R15433 vdd.n441 vdd.t98 303.69
R15434 vdd.n453 vdd.t104 303.69
R15435 vdd.n769 vdd.t120 303.69
R15436 vdd.n3457 vdd.t133 303.69
R15437 vdd.n689 vdd.t110 303.69
R15438 vdd.n3090 vdd.n960 279.512
R15439 vdd.n3330 vdd.n809 279.512
R15440 vdd.n3267 vdd.n806 279.512
R15441 vdd.n3022 vdd.n3021 279.512
R15442 vdd.n2783 vdd.n998 279.512
R15443 vdd.n2714 vdd.n2713 279.512
R15444 vdd.n1355 vdd.n1354 279.512
R15445 vdd.n2508 vdd.n1138 279.512
R15446 vdd.n3246 vdd.n807 279.512
R15447 vdd.n3333 vdd.n3332 279.512
R15448 vdd.n2895 vdd.n2818 279.512
R15449 vdd.n2826 vdd.n956 279.512
R15450 vdd.n2711 vdd.n1008 279.512
R15451 vdd.n1006 vdd.n980 279.512
R15452 vdd.n1480 vdd.n1175 279.512
R15453 vdd.n1280 vdd.n1133 279.512
R15454 vdd.n2506 vdd.n1141 254.619
R15455 vdd.n3495 vdd.n692 254.619
R15456 vdd.n3248 vdd.n807 185
R15457 vdd.n3331 vdd.n807 185
R15458 vdd.n3250 vdd.n3249 185
R15459 vdd.n3249 vdd.n805 185
R15460 vdd.n3251 vdd.n839 185
R15461 vdd.n3261 vdd.n839 185
R15462 vdd.n3252 vdd.n848 185
R15463 vdd.n848 vdd.n846 185
R15464 vdd.n3254 vdd.n3253 185
R15465 vdd.n3255 vdd.n3254 185
R15466 vdd.n3207 vdd.n847 185
R15467 vdd.n847 vdd.n843 185
R15468 vdd.n3206 vdd.n3205 185
R15469 vdd.n3205 vdd.n3204 185
R15470 vdd.n850 vdd.n849 185
R15471 vdd.n851 vdd.n850 185
R15472 vdd.n3197 vdd.n3196 185
R15473 vdd.n3198 vdd.n3197 185
R15474 vdd.n3195 vdd.n859 185
R15475 vdd.n864 vdd.n859 185
R15476 vdd.n3194 vdd.n3193 185
R15477 vdd.n3193 vdd.n3192 185
R15478 vdd.n861 vdd.n860 185
R15479 vdd.n870 vdd.n861 185
R15480 vdd.n3185 vdd.n3184 185
R15481 vdd.n3186 vdd.n3185 185
R15482 vdd.n3183 vdd.n871 185
R15483 vdd.n877 vdd.n871 185
R15484 vdd.n3182 vdd.n3181 185
R15485 vdd.n3181 vdd.n3180 185
R15486 vdd.n873 vdd.n872 185
R15487 vdd.n874 vdd.n873 185
R15488 vdd.n3173 vdd.n3172 185
R15489 vdd.n3174 vdd.n3173 185
R15490 vdd.n3171 vdd.n884 185
R15491 vdd.n884 vdd.n881 185
R15492 vdd.n3170 vdd.n3169 185
R15493 vdd.n3169 vdd.n3168 185
R15494 vdd.n886 vdd.n885 185
R15495 vdd.n887 vdd.n886 185
R15496 vdd.n3161 vdd.n3160 185
R15497 vdd.n3162 vdd.n3161 185
R15498 vdd.n3159 vdd.n895 185
R15499 vdd.n901 vdd.n895 185
R15500 vdd.n3158 vdd.n3157 185
R15501 vdd.n3157 vdd.n3156 185
R15502 vdd.n3147 vdd.n898 185
R15503 vdd.n908 vdd.n898 185
R15504 vdd.n3149 vdd.n3148 185
R15505 vdd.n3150 vdd.n3149 185
R15506 vdd.n3146 vdd.n909 185
R15507 vdd.n909 vdd.n905 185
R15508 vdd.n3145 vdd.n3144 185
R15509 vdd.n3144 vdd.n3143 185
R15510 vdd.n911 vdd.n910 185
R15511 vdd.n912 vdd.n911 185
R15512 vdd.n3136 vdd.n3135 185
R15513 vdd.n3137 vdd.n3136 185
R15514 vdd.n3134 vdd.n920 185
R15515 vdd.n925 vdd.n920 185
R15516 vdd.n3133 vdd.n3132 185
R15517 vdd.n3132 vdd.n3131 185
R15518 vdd.n922 vdd.n921 185
R15519 vdd.n931 vdd.n922 185
R15520 vdd.n3124 vdd.n3123 185
R15521 vdd.n3125 vdd.n3124 185
R15522 vdd.n3122 vdd.n932 185
R15523 vdd.n2998 vdd.n932 185
R15524 vdd.n3121 vdd.n3120 185
R15525 vdd.n3120 vdd.n3119 185
R15526 vdd.n934 vdd.n933 185
R15527 vdd.n3004 vdd.n934 185
R15528 vdd.n3112 vdd.n3111 185
R15529 vdd.n3113 vdd.n3112 185
R15530 vdd.n3110 vdd.n943 185
R15531 vdd.n943 vdd.n940 185
R15532 vdd.n3109 vdd.n3108 185
R15533 vdd.n3108 vdd.n3107 185
R15534 vdd.n945 vdd.n944 185
R15535 vdd.n946 vdd.n945 185
R15536 vdd.n3100 vdd.n3099 185
R15537 vdd.n3101 vdd.n3100 185
R15538 vdd.n3098 vdd.n954 185
R15539 vdd.n3016 vdd.n954 185
R15540 vdd.n3097 vdd.n3096 185
R15541 vdd.n3096 vdd.n3095 185
R15542 vdd.n956 vdd.n955 185
R15543 vdd.n957 vdd.n956 185
R15544 vdd.n2827 vdd.n2826 185
R15545 vdd.n2829 vdd.n2828 185
R15546 vdd.n2831 vdd.n2830 185
R15547 vdd.n2833 vdd.n2832 185
R15548 vdd.n2835 vdd.n2834 185
R15549 vdd.n2837 vdd.n2836 185
R15550 vdd.n2839 vdd.n2838 185
R15551 vdd.n2841 vdd.n2840 185
R15552 vdd.n2843 vdd.n2842 185
R15553 vdd.n2845 vdd.n2844 185
R15554 vdd.n2847 vdd.n2846 185
R15555 vdd.n2849 vdd.n2848 185
R15556 vdd.n2851 vdd.n2850 185
R15557 vdd.n2853 vdd.n2852 185
R15558 vdd.n2855 vdd.n2854 185
R15559 vdd.n2857 vdd.n2856 185
R15560 vdd.n2859 vdd.n2858 185
R15561 vdd.n2861 vdd.n2860 185
R15562 vdd.n2863 vdd.n2862 185
R15563 vdd.n2865 vdd.n2864 185
R15564 vdd.n2867 vdd.n2866 185
R15565 vdd.n2869 vdd.n2868 185
R15566 vdd.n2871 vdd.n2870 185
R15567 vdd.n2873 vdd.n2872 185
R15568 vdd.n2875 vdd.n2874 185
R15569 vdd.n2877 vdd.n2876 185
R15570 vdd.n2879 vdd.n2878 185
R15571 vdd.n2881 vdd.n2880 185
R15572 vdd.n2883 vdd.n2882 185
R15573 vdd.n2885 vdd.n2884 185
R15574 vdd.n2887 vdd.n2886 185
R15575 vdd.n2889 vdd.n2888 185
R15576 vdd.n2891 vdd.n2890 185
R15577 vdd.n2893 vdd.n2892 185
R15578 vdd.n2894 vdd.n2818 185
R15579 vdd.n3088 vdd.n2818 185
R15580 vdd.n3334 vdd.n3333 185
R15581 vdd.n3335 vdd.n798 185
R15582 vdd.n3337 vdd.n3336 185
R15583 vdd.n3339 vdd.n796 185
R15584 vdd.n3341 vdd.n3340 185
R15585 vdd.n3342 vdd.n795 185
R15586 vdd.n3344 vdd.n3343 185
R15587 vdd.n3346 vdd.n793 185
R15588 vdd.n3348 vdd.n3347 185
R15589 vdd.n3349 vdd.n792 185
R15590 vdd.n3351 vdd.n3350 185
R15591 vdd.n3353 vdd.n790 185
R15592 vdd.n3355 vdd.n3354 185
R15593 vdd.n3356 vdd.n789 185
R15594 vdd.n3358 vdd.n3357 185
R15595 vdd.n3360 vdd.n788 185
R15596 vdd.n3361 vdd.n786 185
R15597 vdd.n3364 vdd.n3363 185
R15598 vdd.n787 vdd.n785 185
R15599 vdd.n3220 vdd.n3219 185
R15600 vdd.n3222 vdd.n3221 185
R15601 vdd.n3224 vdd.n3216 185
R15602 vdd.n3226 vdd.n3225 185
R15603 vdd.n3227 vdd.n3215 185
R15604 vdd.n3229 vdd.n3228 185
R15605 vdd.n3231 vdd.n3213 185
R15606 vdd.n3233 vdd.n3232 185
R15607 vdd.n3234 vdd.n3212 185
R15608 vdd.n3236 vdd.n3235 185
R15609 vdd.n3238 vdd.n3210 185
R15610 vdd.n3240 vdd.n3239 185
R15611 vdd.n3241 vdd.n3209 185
R15612 vdd.n3243 vdd.n3242 185
R15613 vdd.n3245 vdd.n3208 185
R15614 vdd.n3247 vdd.n3246 185
R15615 vdd.n3246 vdd.n692 185
R15616 vdd.n3332 vdd.n802 185
R15617 vdd.n3332 vdd.n3331 185
R15618 vdd.n2949 vdd.n804 185
R15619 vdd.n805 vdd.n804 185
R15620 vdd.n2950 vdd.n838 185
R15621 vdd.n3261 vdd.n838 185
R15622 vdd.n2952 vdd.n2951 185
R15623 vdd.n2951 vdd.n846 185
R15624 vdd.n2953 vdd.n845 185
R15625 vdd.n3255 vdd.n845 185
R15626 vdd.n2955 vdd.n2954 185
R15627 vdd.n2954 vdd.n843 185
R15628 vdd.n2956 vdd.n853 185
R15629 vdd.n3204 vdd.n853 185
R15630 vdd.n2958 vdd.n2957 185
R15631 vdd.n2957 vdd.n851 185
R15632 vdd.n2959 vdd.n858 185
R15633 vdd.n3198 vdd.n858 185
R15634 vdd.n2961 vdd.n2960 185
R15635 vdd.n2960 vdd.n864 185
R15636 vdd.n2962 vdd.n863 185
R15637 vdd.n3192 vdd.n863 185
R15638 vdd.n2964 vdd.n2963 185
R15639 vdd.n2963 vdd.n870 185
R15640 vdd.n2965 vdd.n869 185
R15641 vdd.n3186 vdd.n869 185
R15642 vdd.n2967 vdd.n2966 185
R15643 vdd.n2966 vdd.n877 185
R15644 vdd.n2968 vdd.n876 185
R15645 vdd.n3180 vdd.n876 185
R15646 vdd.n2970 vdd.n2969 185
R15647 vdd.n2969 vdd.n874 185
R15648 vdd.n2971 vdd.n883 185
R15649 vdd.n3174 vdd.n883 185
R15650 vdd.n2973 vdd.n2972 185
R15651 vdd.n2972 vdd.n881 185
R15652 vdd.n2974 vdd.n889 185
R15653 vdd.n3168 vdd.n889 185
R15654 vdd.n2976 vdd.n2975 185
R15655 vdd.n2975 vdd.n887 185
R15656 vdd.n2977 vdd.n894 185
R15657 vdd.n3162 vdd.n894 185
R15658 vdd.n2979 vdd.n2978 185
R15659 vdd.n2978 vdd.n901 185
R15660 vdd.n2980 vdd.n900 185
R15661 vdd.n3156 vdd.n900 185
R15662 vdd.n2982 vdd.n2981 185
R15663 vdd.n2981 vdd.n908 185
R15664 vdd.n2983 vdd.n907 185
R15665 vdd.n3150 vdd.n907 185
R15666 vdd.n2985 vdd.n2984 185
R15667 vdd.n2984 vdd.n905 185
R15668 vdd.n2986 vdd.n914 185
R15669 vdd.n3143 vdd.n914 185
R15670 vdd.n2988 vdd.n2987 185
R15671 vdd.n2987 vdd.n912 185
R15672 vdd.n2989 vdd.n919 185
R15673 vdd.n3137 vdd.n919 185
R15674 vdd.n2991 vdd.n2990 185
R15675 vdd.n2990 vdd.n925 185
R15676 vdd.n2992 vdd.n924 185
R15677 vdd.n3131 vdd.n924 185
R15678 vdd.n2994 vdd.n2993 185
R15679 vdd.n2993 vdd.n931 185
R15680 vdd.n2995 vdd.n930 185
R15681 vdd.n3125 vdd.n930 185
R15682 vdd.n2997 vdd.n2996 185
R15683 vdd.n2998 vdd.n2997 185
R15684 vdd.n2898 vdd.n936 185
R15685 vdd.n3119 vdd.n936 185
R15686 vdd.n3006 vdd.n3005 185
R15687 vdd.n3005 vdd.n3004 185
R15688 vdd.n3007 vdd.n942 185
R15689 vdd.n3113 vdd.n942 185
R15690 vdd.n3009 vdd.n3008 185
R15691 vdd.n3008 vdd.n940 185
R15692 vdd.n3010 vdd.n948 185
R15693 vdd.n3107 vdd.n948 185
R15694 vdd.n3012 vdd.n3011 185
R15695 vdd.n3011 vdd.n946 185
R15696 vdd.n3013 vdd.n953 185
R15697 vdd.n3101 vdd.n953 185
R15698 vdd.n3015 vdd.n3014 185
R15699 vdd.n3016 vdd.n3015 185
R15700 vdd.n2897 vdd.n959 185
R15701 vdd.n3095 vdd.n959 185
R15702 vdd.n2896 vdd.n2895 185
R15703 vdd.n2895 vdd.n957 185
R15704 vdd.n2357 vdd.n2356 185
R15705 vdd.n2358 vdd.n2357 185
R15706 vdd.n1531 vdd.n1529 185
R15707 vdd.n2349 vdd.n1529 185
R15708 vdd.n2352 vdd.n2351 185
R15709 vdd.n2351 vdd.n2350 185
R15710 vdd.n1534 vdd.n1533 185
R15711 vdd.n1535 vdd.n1534 185
R15712 vdd.n2338 vdd.n2337 185
R15713 vdd.n2339 vdd.n2338 185
R15714 vdd.n1543 vdd.n1542 185
R15715 vdd.n2330 vdd.n1542 185
R15716 vdd.n2333 vdd.n2332 185
R15717 vdd.n2332 vdd.n2331 185
R15718 vdd.n1546 vdd.n1545 185
R15719 vdd.n1553 vdd.n1546 185
R15720 vdd.n2321 vdd.n2320 185
R15721 vdd.n2322 vdd.n2321 185
R15722 vdd.n1555 vdd.n1554 185
R15723 vdd.n1554 vdd.n1552 185
R15724 vdd.n2316 vdd.n2315 185
R15725 vdd.n2315 vdd.n2314 185
R15726 vdd.n1558 vdd.n1557 185
R15727 vdd.n1559 vdd.n1558 185
R15728 vdd.n2305 vdd.n2304 185
R15729 vdd.n2306 vdd.n2305 185
R15730 vdd.n1566 vdd.n1565 185
R15731 vdd.n2297 vdd.n1565 185
R15732 vdd.n2300 vdd.n2299 185
R15733 vdd.n2299 vdd.n2298 185
R15734 vdd.n1569 vdd.n1568 185
R15735 vdd.n1575 vdd.n1569 185
R15736 vdd.n2288 vdd.n2287 185
R15737 vdd.n2289 vdd.n2288 185
R15738 vdd.n1577 vdd.n1576 185
R15739 vdd.n2280 vdd.n1576 185
R15740 vdd.n2283 vdd.n2282 185
R15741 vdd.n2282 vdd.n2281 185
R15742 vdd.n1580 vdd.n1579 185
R15743 vdd.n1581 vdd.n1580 185
R15744 vdd.n2271 vdd.n2270 185
R15745 vdd.n2272 vdd.n2271 185
R15746 vdd.n1589 vdd.n1588 185
R15747 vdd.n1588 vdd.n1587 185
R15748 vdd.n1959 vdd.n1958 185
R15749 vdd.n1958 vdd.n1957 185
R15750 vdd.n1592 vdd.n1591 185
R15751 vdd.n1598 vdd.n1592 185
R15752 vdd.n1948 vdd.n1947 185
R15753 vdd.n1949 vdd.n1948 185
R15754 vdd.n1600 vdd.n1599 185
R15755 vdd.n1940 vdd.n1599 185
R15756 vdd.n1943 vdd.n1942 185
R15757 vdd.n1942 vdd.n1941 185
R15758 vdd.n1603 vdd.n1602 185
R15759 vdd.n1610 vdd.n1603 185
R15760 vdd.n1931 vdd.n1930 185
R15761 vdd.n1932 vdd.n1931 185
R15762 vdd.n1612 vdd.n1611 185
R15763 vdd.n1611 vdd.n1609 185
R15764 vdd.n1926 vdd.n1925 185
R15765 vdd.n1925 vdd.n1924 185
R15766 vdd.n1615 vdd.n1614 185
R15767 vdd.n1616 vdd.n1615 185
R15768 vdd.n1915 vdd.n1914 185
R15769 vdd.n1916 vdd.n1915 185
R15770 vdd.n1623 vdd.n1622 185
R15771 vdd.n1907 vdd.n1622 185
R15772 vdd.n1910 vdd.n1909 185
R15773 vdd.n1909 vdd.n1908 185
R15774 vdd.n1626 vdd.n1625 185
R15775 vdd.n1632 vdd.n1626 185
R15776 vdd.n1898 vdd.n1897 185
R15777 vdd.n1899 vdd.n1898 185
R15778 vdd.n1634 vdd.n1633 185
R15779 vdd.n1890 vdd.n1633 185
R15780 vdd.n1893 vdd.n1892 185
R15781 vdd.n1892 vdd.n1891 185
R15782 vdd.n1637 vdd.n1636 185
R15783 vdd.n1638 vdd.n1637 185
R15784 vdd.n1881 vdd.n1880 185
R15785 vdd.n1882 vdd.n1881 185
R15786 vdd.n1645 vdd.n1644 185
R15787 vdd.n1680 vdd.n1644 185
R15788 vdd.n1876 vdd.n1875 185
R15789 vdd.n1648 vdd.n1647 185
R15790 vdd.n1872 vdd.n1871 185
R15791 vdd.n1873 vdd.n1872 185
R15792 vdd.n1682 vdd.n1681 185
R15793 vdd.n1867 vdd.n1684 185
R15794 vdd.n1866 vdd.n1685 185
R15795 vdd.n1865 vdd.n1686 185
R15796 vdd.n1688 vdd.n1687 185
R15797 vdd.n1861 vdd.n1690 185
R15798 vdd.n1860 vdd.n1691 185
R15799 vdd.n1859 vdd.n1692 185
R15800 vdd.n1694 vdd.n1693 185
R15801 vdd.n1855 vdd.n1696 185
R15802 vdd.n1854 vdd.n1697 185
R15803 vdd.n1853 vdd.n1698 185
R15804 vdd.n1700 vdd.n1699 185
R15805 vdd.n1849 vdd.n1702 185
R15806 vdd.n1848 vdd.n1703 185
R15807 vdd.n1847 vdd.n1704 185
R15808 vdd.n1708 vdd.n1705 185
R15809 vdd.n1843 vdd.n1710 185
R15810 vdd.n1842 vdd.n1711 185
R15811 vdd.n1841 vdd.n1712 185
R15812 vdd.n1714 vdd.n1713 185
R15813 vdd.n1837 vdd.n1716 185
R15814 vdd.n1836 vdd.n1717 185
R15815 vdd.n1835 vdd.n1718 185
R15816 vdd.n1720 vdd.n1719 185
R15817 vdd.n1831 vdd.n1722 185
R15818 vdd.n1830 vdd.n1723 185
R15819 vdd.n1829 vdd.n1724 185
R15820 vdd.n1726 vdd.n1725 185
R15821 vdd.n1825 vdd.n1728 185
R15822 vdd.n1824 vdd.n1729 185
R15823 vdd.n1823 vdd.n1730 185
R15824 vdd.n1732 vdd.n1731 185
R15825 vdd.n1819 vdd.n1734 185
R15826 vdd.n1818 vdd.n1735 185
R15827 vdd.n1817 vdd.n1736 185
R15828 vdd.n1738 vdd.n1737 185
R15829 vdd.n1813 vdd.n1740 185
R15830 vdd.n1812 vdd.n1809 185
R15831 vdd.n1808 vdd.n1741 185
R15832 vdd.n1743 vdd.n1742 185
R15833 vdd.n1804 vdd.n1745 185
R15834 vdd.n1803 vdd.n1746 185
R15835 vdd.n1802 vdd.n1747 185
R15836 vdd.n1749 vdd.n1748 185
R15837 vdd.n1798 vdd.n1751 185
R15838 vdd.n1797 vdd.n1752 185
R15839 vdd.n1796 vdd.n1753 185
R15840 vdd.n1755 vdd.n1754 185
R15841 vdd.n1792 vdd.n1757 185
R15842 vdd.n1791 vdd.n1758 185
R15843 vdd.n1790 vdd.n1759 185
R15844 vdd.n1761 vdd.n1760 185
R15845 vdd.n1786 vdd.n1763 185
R15846 vdd.n1785 vdd.n1764 185
R15847 vdd.n1784 vdd.n1765 185
R15848 vdd.n1767 vdd.n1766 185
R15849 vdd.n1780 vdd.n1769 185
R15850 vdd.n1779 vdd.n1770 185
R15851 vdd.n1778 vdd.n1771 185
R15852 vdd.n1775 vdd.n1679 185
R15853 vdd.n1873 vdd.n1679 185
R15854 vdd.n2361 vdd.n2360 185
R15855 vdd.n2365 vdd.n1525 185
R15856 vdd.n1524 vdd.n1518 185
R15857 vdd.n1522 vdd.n1521 185
R15858 vdd.n1520 vdd.n1279 185
R15859 vdd.n2369 vdd.n1276 185
R15860 vdd.n2371 vdd.n2370 185
R15861 vdd.n2373 vdd.n1274 185
R15862 vdd.n2375 vdd.n2374 185
R15863 vdd.n2376 vdd.n1269 185
R15864 vdd.n2378 vdd.n2377 185
R15865 vdd.n2380 vdd.n1267 185
R15866 vdd.n2382 vdd.n2381 185
R15867 vdd.n2383 vdd.n1262 185
R15868 vdd.n2385 vdd.n2384 185
R15869 vdd.n2387 vdd.n1260 185
R15870 vdd.n2389 vdd.n2388 185
R15871 vdd.n2390 vdd.n1256 185
R15872 vdd.n2392 vdd.n2391 185
R15873 vdd.n2394 vdd.n1253 185
R15874 vdd.n2396 vdd.n2395 185
R15875 vdd.n1254 vdd.n1247 185
R15876 vdd.n2400 vdd.n1251 185
R15877 vdd.n2401 vdd.n1243 185
R15878 vdd.n2403 vdd.n2402 185
R15879 vdd.n2405 vdd.n1241 185
R15880 vdd.n2407 vdd.n2406 185
R15881 vdd.n2408 vdd.n1236 185
R15882 vdd.n2410 vdd.n2409 185
R15883 vdd.n2412 vdd.n1234 185
R15884 vdd.n2414 vdd.n2413 185
R15885 vdd.n2415 vdd.n1229 185
R15886 vdd.n2417 vdd.n2416 185
R15887 vdd.n2419 vdd.n1227 185
R15888 vdd.n2421 vdd.n2420 185
R15889 vdd.n2422 vdd.n1222 185
R15890 vdd.n2424 vdd.n2423 185
R15891 vdd.n2426 vdd.n1220 185
R15892 vdd.n2428 vdd.n2427 185
R15893 vdd.n2429 vdd.n1216 185
R15894 vdd.n2431 vdd.n2430 185
R15895 vdd.n2433 vdd.n1213 185
R15896 vdd.n2435 vdd.n2434 185
R15897 vdd.n1214 vdd.n1207 185
R15898 vdd.n2439 vdd.n1211 185
R15899 vdd.n2440 vdd.n1203 185
R15900 vdd.n2442 vdd.n2441 185
R15901 vdd.n2444 vdd.n1201 185
R15902 vdd.n2446 vdd.n2445 185
R15903 vdd.n2447 vdd.n1196 185
R15904 vdd.n2449 vdd.n2448 185
R15905 vdd.n2451 vdd.n1194 185
R15906 vdd.n2453 vdd.n2452 185
R15907 vdd.n2454 vdd.n1189 185
R15908 vdd.n2456 vdd.n2455 185
R15909 vdd.n2458 vdd.n1187 185
R15910 vdd.n2460 vdd.n2459 185
R15911 vdd.n2461 vdd.n1185 185
R15912 vdd.n2463 vdd.n2462 185
R15913 vdd.n2466 vdd.n2465 185
R15914 vdd.n2468 vdd.n2467 185
R15915 vdd.n2470 vdd.n1183 185
R15916 vdd.n2472 vdd.n2471 185
R15917 vdd.n1530 vdd.n1182 185
R15918 vdd.n2359 vdd.n1528 185
R15919 vdd.n2359 vdd.n2358 185
R15920 vdd.n1538 vdd.n1527 185
R15921 vdd.n2349 vdd.n1527 185
R15922 vdd.n2348 vdd.n2347 185
R15923 vdd.n2350 vdd.n2348 185
R15924 vdd.n1537 vdd.n1536 185
R15925 vdd.n1536 vdd.n1535 185
R15926 vdd.n2341 vdd.n2340 185
R15927 vdd.n2340 vdd.n2339 185
R15928 vdd.n1541 vdd.n1540 185
R15929 vdd.n2330 vdd.n1541 185
R15930 vdd.n2329 vdd.n2328 185
R15931 vdd.n2331 vdd.n2329 185
R15932 vdd.n1548 vdd.n1547 185
R15933 vdd.n1553 vdd.n1547 185
R15934 vdd.n2324 vdd.n2323 185
R15935 vdd.n2323 vdd.n2322 185
R15936 vdd.n1551 vdd.n1550 185
R15937 vdd.n1552 vdd.n1551 185
R15938 vdd.n2313 vdd.n2312 185
R15939 vdd.n2314 vdd.n2313 185
R15940 vdd.n1561 vdd.n1560 185
R15941 vdd.n1560 vdd.n1559 185
R15942 vdd.n2308 vdd.n2307 185
R15943 vdd.n2307 vdd.n2306 185
R15944 vdd.n1564 vdd.n1563 185
R15945 vdd.n2297 vdd.n1564 185
R15946 vdd.n2296 vdd.n2295 185
R15947 vdd.n2298 vdd.n2296 185
R15948 vdd.n1571 vdd.n1570 185
R15949 vdd.n1575 vdd.n1570 185
R15950 vdd.n2291 vdd.n2290 185
R15951 vdd.n2290 vdd.n2289 185
R15952 vdd.n1574 vdd.n1573 185
R15953 vdd.n2280 vdd.n1574 185
R15954 vdd.n2279 vdd.n2278 185
R15955 vdd.n2281 vdd.n2279 185
R15956 vdd.n1583 vdd.n1582 185
R15957 vdd.n1582 vdd.n1581 185
R15958 vdd.n2274 vdd.n2273 185
R15959 vdd.n2273 vdd.n2272 185
R15960 vdd.n1586 vdd.n1585 185
R15961 vdd.n1587 vdd.n1586 185
R15962 vdd.n1956 vdd.n1955 185
R15963 vdd.n1957 vdd.n1956 185
R15964 vdd.n1594 vdd.n1593 185
R15965 vdd.n1598 vdd.n1593 185
R15966 vdd.n1951 vdd.n1950 185
R15967 vdd.n1950 vdd.n1949 185
R15968 vdd.n1597 vdd.n1596 185
R15969 vdd.n1940 vdd.n1597 185
R15970 vdd.n1939 vdd.n1938 185
R15971 vdd.n1941 vdd.n1939 185
R15972 vdd.n1605 vdd.n1604 185
R15973 vdd.n1610 vdd.n1604 185
R15974 vdd.n1934 vdd.n1933 185
R15975 vdd.n1933 vdd.n1932 185
R15976 vdd.n1608 vdd.n1607 185
R15977 vdd.n1609 vdd.n1608 185
R15978 vdd.n1923 vdd.n1922 185
R15979 vdd.n1924 vdd.n1923 185
R15980 vdd.n1618 vdd.n1617 185
R15981 vdd.n1617 vdd.n1616 185
R15982 vdd.n1918 vdd.n1917 185
R15983 vdd.n1917 vdd.n1916 185
R15984 vdd.n1621 vdd.n1620 185
R15985 vdd.n1907 vdd.n1621 185
R15986 vdd.n1906 vdd.n1905 185
R15987 vdd.n1908 vdd.n1906 185
R15988 vdd.n1628 vdd.n1627 185
R15989 vdd.n1632 vdd.n1627 185
R15990 vdd.n1901 vdd.n1900 185
R15991 vdd.n1900 vdd.n1899 185
R15992 vdd.n1631 vdd.n1630 185
R15993 vdd.n1890 vdd.n1631 185
R15994 vdd.n1889 vdd.n1888 185
R15995 vdd.n1891 vdd.n1889 185
R15996 vdd.n1640 vdd.n1639 185
R15997 vdd.n1639 vdd.n1638 185
R15998 vdd.n1884 vdd.n1883 185
R15999 vdd.n1883 vdd.n1882 185
R16000 vdd.n1643 vdd.n1642 185
R16001 vdd.n1680 vdd.n1643 185
R16002 vdd.n1000 vdd.n998 185
R16003 vdd.n2712 vdd.n998 185
R16004 vdd.n2634 vdd.n1018 185
R16005 vdd.n1018 vdd.n1005 185
R16006 vdd.n2636 vdd.n2635 185
R16007 vdd.n2637 vdd.n2636 185
R16008 vdd.n2633 vdd.n1017 185
R16009 vdd.n1399 vdd.n1017 185
R16010 vdd.n2632 vdd.n2631 185
R16011 vdd.n2631 vdd.n2630 185
R16012 vdd.n1020 vdd.n1019 185
R16013 vdd.n1021 vdd.n1020 185
R16014 vdd.n2621 vdd.n2620 185
R16015 vdd.n2622 vdd.n2621 185
R16016 vdd.n2619 vdd.n1031 185
R16017 vdd.n1031 vdd.n1028 185
R16018 vdd.n2618 vdd.n2617 185
R16019 vdd.n2617 vdd.n2616 185
R16020 vdd.n1033 vdd.n1032 185
R16021 vdd.n1425 vdd.n1033 185
R16022 vdd.n2609 vdd.n2608 185
R16023 vdd.n2610 vdd.n2609 185
R16024 vdd.n2607 vdd.n1041 185
R16025 vdd.n1046 vdd.n1041 185
R16026 vdd.n2606 vdd.n2605 185
R16027 vdd.n2605 vdd.n2604 185
R16028 vdd.n1043 vdd.n1042 185
R16029 vdd.n1052 vdd.n1043 185
R16030 vdd.n2597 vdd.n2596 185
R16031 vdd.n2598 vdd.n2597 185
R16032 vdd.n2595 vdd.n1053 185
R16033 vdd.n1437 vdd.n1053 185
R16034 vdd.n2594 vdd.n2593 185
R16035 vdd.n2593 vdd.n2592 185
R16036 vdd.n1055 vdd.n1054 185
R16037 vdd.n1056 vdd.n1055 185
R16038 vdd.n2585 vdd.n2584 185
R16039 vdd.n2586 vdd.n2585 185
R16040 vdd.n2583 vdd.n1065 185
R16041 vdd.n1065 vdd.n1062 185
R16042 vdd.n2582 vdd.n2581 185
R16043 vdd.n2581 vdd.n2580 185
R16044 vdd.n1067 vdd.n1066 185
R16045 vdd.n1076 vdd.n1067 185
R16046 vdd.n2572 vdd.n2571 185
R16047 vdd.n2573 vdd.n2572 185
R16048 vdd.n2570 vdd.n1077 185
R16049 vdd.n1083 vdd.n1077 185
R16050 vdd.n2569 vdd.n2568 185
R16051 vdd.n2568 vdd.n2567 185
R16052 vdd.n1079 vdd.n1078 185
R16053 vdd.n1080 vdd.n1079 185
R16054 vdd.n2560 vdd.n2559 185
R16055 vdd.n2561 vdd.n2560 185
R16056 vdd.n2558 vdd.n1090 185
R16057 vdd.n1090 vdd.n1087 185
R16058 vdd.n2557 vdd.n2556 185
R16059 vdd.n2556 vdd.n2555 185
R16060 vdd.n1092 vdd.n1091 185
R16061 vdd.n1093 vdd.n1092 185
R16062 vdd.n2548 vdd.n2547 185
R16063 vdd.n2549 vdd.n2548 185
R16064 vdd.n2546 vdd.n1101 185
R16065 vdd.n1106 vdd.n1101 185
R16066 vdd.n2545 vdd.n2544 185
R16067 vdd.n2544 vdd.n2543 185
R16068 vdd.n1103 vdd.n1102 185
R16069 vdd.n1112 vdd.n1103 185
R16070 vdd.n2536 vdd.n2535 185
R16071 vdd.n2537 vdd.n2536 185
R16072 vdd.n2534 vdd.n1113 185
R16073 vdd.n1119 vdd.n1113 185
R16074 vdd.n2533 vdd.n2532 185
R16075 vdd.n2532 vdd.n2531 185
R16076 vdd.n1115 vdd.n1114 185
R16077 vdd.n1116 vdd.n1115 185
R16078 vdd.n2524 vdd.n2523 185
R16079 vdd.n2525 vdd.n2524 185
R16080 vdd.n2522 vdd.n1126 185
R16081 vdd.n1126 vdd.n1123 185
R16082 vdd.n2521 vdd.n2520 185
R16083 vdd.n2520 vdd.n2519 185
R16084 vdd.n1128 vdd.n1127 185
R16085 vdd.n1137 vdd.n1128 185
R16086 vdd.n2512 vdd.n2511 185
R16087 vdd.n2513 vdd.n2512 185
R16088 vdd.n2510 vdd.n1138 185
R16089 vdd.n1138 vdd.n1134 185
R16090 vdd.n2509 vdd.n2508 185
R16091 vdd.n1140 vdd.n1139 185
R16092 vdd.n2505 vdd.n2504 185
R16093 vdd.n2506 vdd.n2505 185
R16094 vdd.n2503 vdd.n1176 185
R16095 vdd.n2502 vdd.n2501 185
R16096 vdd.n2500 vdd.n2499 185
R16097 vdd.n2498 vdd.n2497 185
R16098 vdd.n2496 vdd.n2495 185
R16099 vdd.n2494 vdd.n2493 185
R16100 vdd.n2492 vdd.n2491 185
R16101 vdd.n2490 vdd.n2489 185
R16102 vdd.n2488 vdd.n2487 185
R16103 vdd.n2486 vdd.n2485 185
R16104 vdd.n2484 vdd.n2483 185
R16105 vdd.n2482 vdd.n2481 185
R16106 vdd.n2480 vdd.n2479 185
R16107 vdd.n2478 vdd.n2477 185
R16108 vdd.n2476 vdd.n2475 185
R16109 vdd.n1321 vdd.n1177 185
R16110 vdd.n1323 vdd.n1322 185
R16111 vdd.n1325 vdd.n1324 185
R16112 vdd.n1327 vdd.n1326 185
R16113 vdd.n1329 vdd.n1328 185
R16114 vdd.n1331 vdd.n1330 185
R16115 vdd.n1333 vdd.n1332 185
R16116 vdd.n1335 vdd.n1334 185
R16117 vdd.n1337 vdd.n1336 185
R16118 vdd.n1339 vdd.n1338 185
R16119 vdd.n1341 vdd.n1340 185
R16120 vdd.n1343 vdd.n1342 185
R16121 vdd.n1345 vdd.n1344 185
R16122 vdd.n1347 vdd.n1346 185
R16123 vdd.n1350 vdd.n1349 185
R16124 vdd.n1352 vdd.n1351 185
R16125 vdd.n1354 vdd.n1353 185
R16126 vdd.n2715 vdd.n2714 185
R16127 vdd.n2717 vdd.n2716 185
R16128 vdd.n2719 vdd.n2718 185
R16129 vdd.n2722 vdd.n2721 185
R16130 vdd.n2724 vdd.n2723 185
R16131 vdd.n2726 vdd.n2725 185
R16132 vdd.n2728 vdd.n2727 185
R16133 vdd.n2730 vdd.n2729 185
R16134 vdd.n2732 vdd.n2731 185
R16135 vdd.n2734 vdd.n2733 185
R16136 vdd.n2736 vdd.n2735 185
R16137 vdd.n2738 vdd.n2737 185
R16138 vdd.n2740 vdd.n2739 185
R16139 vdd.n2742 vdd.n2741 185
R16140 vdd.n2744 vdd.n2743 185
R16141 vdd.n2746 vdd.n2745 185
R16142 vdd.n2748 vdd.n2747 185
R16143 vdd.n2750 vdd.n2749 185
R16144 vdd.n2752 vdd.n2751 185
R16145 vdd.n2754 vdd.n2753 185
R16146 vdd.n2756 vdd.n2755 185
R16147 vdd.n2758 vdd.n2757 185
R16148 vdd.n2760 vdd.n2759 185
R16149 vdd.n2762 vdd.n2761 185
R16150 vdd.n2764 vdd.n2763 185
R16151 vdd.n2766 vdd.n2765 185
R16152 vdd.n2768 vdd.n2767 185
R16153 vdd.n2770 vdd.n2769 185
R16154 vdd.n2772 vdd.n2771 185
R16155 vdd.n2774 vdd.n2773 185
R16156 vdd.n2776 vdd.n2775 185
R16157 vdd.n2778 vdd.n2777 185
R16158 vdd.n2780 vdd.n2779 185
R16159 vdd.n2781 vdd.n999 185
R16160 vdd.n2783 vdd.n2782 185
R16161 vdd.n2784 vdd.n2783 185
R16162 vdd.n2713 vdd.n1003 185
R16163 vdd.n2713 vdd.n2712 185
R16164 vdd.n1397 vdd.n1004 185
R16165 vdd.n1005 vdd.n1004 185
R16166 vdd.n1398 vdd.n1015 185
R16167 vdd.n2637 vdd.n1015 185
R16168 vdd.n1401 vdd.n1400 185
R16169 vdd.n1400 vdd.n1399 185
R16170 vdd.n1402 vdd.n1022 185
R16171 vdd.n2630 vdd.n1022 185
R16172 vdd.n1404 vdd.n1403 185
R16173 vdd.n1403 vdd.n1021 185
R16174 vdd.n1405 vdd.n1029 185
R16175 vdd.n2622 vdd.n1029 185
R16176 vdd.n1407 vdd.n1406 185
R16177 vdd.n1406 vdd.n1028 185
R16178 vdd.n1408 vdd.n1034 185
R16179 vdd.n2616 vdd.n1034 185
R16180 vdd.n1427 vdd.n1426 185
R16181 vdd.n1426 vdd.n1425 185
R16182 vdd.n1428 vdd.n1039 185
R16183 vdd.n2610 vdd.n1039 185
R16184 vdd.n1430 vdd.n1429 185
R16185 vdd.n1429 vdd.n1046 185
R16186 vdd.n1431 vdd.n1044 185
R16187 vdd.n2604 vdd.n1044 185
R16188 vdd.n1433 vdd.n1432 185
R16189 vdd.n1432 vdd.n1052 185
R16190 vdd.n1434 vdd.n1050 185
R16191 vdd.n2598 vdd.n1050 185
R16192 vdd.n1436 vdd.n1435 185
R16193 vdd.n1437 vdd.n1436 185
R16194 vdd.n1396 vdd.n1057 185
R16195 vdd.n2592 vdd.n1057 185
R16196 vdd.n1395 vdd.n1394 185
R16197 vdd.n1394 vdd.n1056 185
R16198 vdd.n1393 vdd.n1063 185
R16199 vdd.n2586 vdd.n1063 185
R16200 vdd.n1392 vdd.n1391 185
R16201 vdd.n1391 vdd.n1062 185
R16202 vdd.n1390 vdd.n1068 185
R16203 vdd.n2580 vdd.n1068 185
R16204 vdd.n1389 vdd.n1388 185
R16205 vdd.n1388 vdd.n1076 185
R16206 vdd.n1387 vdd.n1074 185
R16207 vdd.n2573 vdd.n1074 185
R16208 vdd.n1386 vdd.n1385 185
R16209 vdd.n1385 vdd.n1083 185
R16210 vdd.n1384 vdd.n1081 185
R16211 vdd.n2567 vdd.n1081 185
R16212 vdd.n1383 vdd.n1382 185
R16213 vdd.n1382 vdd.n1080 185
R16214 vdd.n1381 vdd.n1088 185
R16215 vdd.n2561 vdd.n1088 185
R16216 vdd.n1380 vdd.n1379 185
R16217 vdd.n1379 vdd.n1087 185
R16218 vdd.n1378 vdd.n1094 185
R16219 vdd.n2555 vdd.n1094 185
R16220 vdd.n1377 vdd.n1376 185
R16221 vdd.n1376 vdd.n1093 185
R16222 vdd.n1375 vdd.n1099 185
R16223 vdd.n2549 vdd.n1099 185
R16224 vdd.n1374 vdd.n1373 185
R16225 vdd.n1373 vdd.n1106 185
R16226 vdd.n1372 vdd.n1104 185
R16227 vdd.n2543 vdd.n1104 185
R16228 vdd.n1371 vdd.n1370 185
R16229 vdd.n1370 vdd.n1112 185
R16230 vdd.n1369 vdd.n1110 185
R16231 vdd.n2537 vdd.n1110 185
R16232 vdd.n1368 vdd.n1367 185
R16233 vdd.n1367 vdd.n1119 185
R16234 vdd.n1366 vdd.n1117 185
R16235 vdd.n2531 vdd.n1117 185
R16236 vdd.n1365 vdd.n1364 185
R16237 vdd.n1364 vdd.n1116 185
R16238 vdd.n1363 vdd.n1124 185
R16239 vdd.n2525 vdd.n1124 185
R16240 vdd.n1362 vdd.n1361 185
R16241 vdd.n1361 vdd.n1123 185
R16242 vdd.n1360 vdd.n1129 185
R16243 vdd.n2519 vdd.n1129 185
R16244 vdd.n1359 vdd.n1358 185
R16245 vdd.n1358 vdd.n1137 185
R16246 vdd.n1357 vdd.n1135 185
R16247 vdd.n2513 vdd.n1135 185
R16248 vdd.n1356 vdd.n1355 185
R16249 vdd.n1355 vdd.n1134 185
R16250 vdd.n3629 vdd.n3628 185
R16251 vdd.n3628 vdd.n3627 185
R16252 vdd.n3630 vdd.n387 185
R16253 vdd.n387 vdd.n386 185
R16254 vdd.n3632 vdd.n3631 185
R16255 vdd.n3633 vdd.n3632 185
R16256 vdd.n382 vdd.n381 185
R16257 vdd.n3634 vdd.n382 185
R16258 vdd.n3637 vdd.n3636 185
R16259 vdd.n3636 vdd.n3635 185
R16260 vdd.n3638 vdd.n376 185
R16261 vdd.n376 vdd.n375 185
R16262 vdd.n3640 vdd.n3639 185
R16263 vdd.n3641 vdd.n3640 185
R16264 vdd.n371 vdd.n370 185
R16265 vdd.n3642 vdd.n371 185
R16266 vdd.n3645 vdd.n3644 185
R16267 vdd.n3644 vdd.n3643 185
R16268 vdd.n3646 vdd.n365 185
R16269 vdd.n3603 vdd.n365 185
R16270 vdd.n3648 vdd.n3647 185
R16271 vdd.n3649 vdd.n3648 185
R16272 vdd.n360 vdd.n359 185
R16273 vdd.n3650 vdd.n360 185
R16274 vdd.n3653 vdd.n3652 185
R16275 vdd.n3652 vdd.n3651 185
R16276 vdd.n3654 vdd.n354 185
R16277 vdd.n361 vdd.n354 185
R16278 vdd.n3656 vdd.n3655 185
R16279 vdd.n3657 vdd.n3656 185
R16280 vdd.n350 vdd.n349 185
R16281 vdd.n3658 vdd.n350 185
R16282 vdd.n3661 vdd.n3660 185
R16283 vdd.n3660 vdd.n3659 185
R16284 vdd.n3662 vdd.n345 185
R16285 vdd.n345 vdd.n344 185
R16286 vdd.n3664 vdd.n3663 185
R16287 vdd.n3665 vdd.n3664 185
R16288 vdd.n339 vdd.n337 185
R16289 vdd.n3666 vdd.n339 185
R16290 vdd.n3669 vdd.n3668 185
R16291 vdd.n3668 vdd.n3667 185
R16292 vdd.n338 vdd.n336 185
R16293 vdd.n340 vdd.n338 185
R16294 vdd.n3579 vdd.n3578 185
R16295 vdd.n3580 vdd.n3579 185
R16296 vdd.n635 vdd.n634 185
R16297 vdd.n634 vdd.n633 185
R16298 vdd.n3574 vdd.n3573 185
R16299 vdd.n3573 vdd.n3572 185
R16300 vdd.n638 vdd.n637 185
R16301 vdd.n644 vdd.n638 185
R16302 vdd.n3560 vdd.n3559 185
R16303 vdd.n3561 vdd.n3560 185
R16304 vdd.n646 vdd.n645 185
R16305 vdd.n3552 vdd.n645 185
R16306 vdd.n3555 vdd.n3554 185
R16307 vdd.n3554 vdd.n3553 185
R16308 vdd.n649 vdd.n648 185
R16309 vdd.n656 vdd.n649 185
R16310 vdd.n3543 vdd.n3542 185
R16311 vdd.n3544 vdd.n3543 185
R16312 vdd.n658 vdd.n657 185
R16313 vdd.n657 vdd.n655 185
R16314 vdd.n3538 vdd.n3537 185
R16315 vdd.n3537 vdd.n3536 185
R16316 vdd.n661 vdd.n660 185
R16317 vdd.n662 vdd.n661 185
R16318 vdd.n3527 vdd.n3526 185
R16319 vdd.n3528 vdd.n3527 185
R16320 vdd.n669 vdd.n668 185
R16321 vdd.n3519 vdd.n668 185
R16322 vdd.n3522 vdd.n3521 185
R16323 vdd.n3521 vdd.n3520 185
R16324 vdd.n672 vdd.n671 185
R16325 vdd.n679 vdd.n672 185
R16326 vdd.n3510 vdd.n3509 185
R16327 vdd.n3511 vdd.n3510 185
R16328 vdd.n681 vdd.n680 185
R16329 vdd.n680 vdd.n678 185
R16330 vdd.n3505 vdd.n3504 185
R16331 vdd.n3504 vdd.n3503 185
R16332 vdd.n684 vdd.n683 185
R16333 vdd.n723 vdd.n684 185
R16334 vdd.n3493 vdd.n3492 185
R16335 vdd.n3491 vdd.n725 185
R16336 vdd.n3490 vdd.n724 185
R16337 vdd.n3495 vdd.n724 185
R16338 vdd.n729 vdd.n728 185
R16339 vdd.n733 vdd.n732 185
R16340 vdd.n3486 vdd.n734 185
R16341 vdd.n3485 vdd.n3484 185
R16342 vdd.n3483 vdd.n3482 185
R16343 vdd.n3481 vdd.n3480 185
R16344 vdd.n3479 vdd.n3478 185
R16345 vdd.n3477 vdd.n3476 185
R16346 vdd.n3475 vdd.n3474 185
R16347 vdd.n3473 vdd.n3472 185
R16348 vdd.n3471 vdd.n3470 185
R16349 vdd.n3469 vdd.n3468 185
R16350 vdd.n3467 vdd.n3466 185
R16351 vdd.n3465 vdd.n3464 185
R16352 vdd.n3463 vdd.n3462 185
R16353 vdd.n3461 vdd.n3460 185
R16354 vdd.n3459 vdd.n3458 185
R16355 vdd.n3450 vdd.n747 185
R16356 vdd.n3452 vdd.n3451 185
R16357 vdd.n3449 vdd.n3448 185
R16358 vdd.n3447 vdd.n3446 185
R16359 vdd.n3445 vdd.n3444 185
R16360 vdd.n3443 vdd.n3442 185
R16361 vdd.n3441 vdd.n3440 185
R16362 vdd.n3439 vdd.n3438 185
R16363 vdd.n3437 vdd.n3436 185
R16364 vdd.n3435 vdd.n3434 185
R16365 vdd.n3433 vdd.n3432 185
R16366 vdd.n3431 vdd.n3430 185
R16367 vdd.n3429 vdd.n3428 185
R16368 vdd.n3427 vdd.n3426 185
R16369 vdd.n3425 vdd.n3424 185
R16370 vdd.n3423 vdd.n3422 185
R16371 vdd.n3421 vdd.n3420 185
R16372 vdd.n3419 vdd.n3418 185
R16373 vdd.n3417 vdd.n3416 185
R16374 vdd.n3415 vdd.n3414 185
R16375 vdd.n3413 vdd.n3412 185
R16376 vdd.n3411 vdd.n3410 185
R16377 vdd.n3404 vdd.n767 185
R16378 vdd.n3406 vdd.n3405 185
R16379 vdd.n3403 vdd.n3402 185
R16380 vdd.n3401 vdd.n3400 185
R16381 vdd.n3399 vdd.n3398 185
R16382 vdd.n3397 vdd.n3396 185
R16383 vdd.n3395 vdd.n3394 185
R16384 vdd.n3393 vdd.n3392 185
R16385 vdd.n3391 vdd.n3390 185
R16386 vdd.n3389 vdd.n3388 185
R16387 vdd.n3387 vdd.n3386 185
R16388 vdd.n3385 vdd.n3384 185
R16389 vdd.n3383 vdd.n3382 185
R16390 vdd.n3381 vdd.n3380 185
R16391 vdd.n3379 vdd.n3378 185
R16392 vdd.n3377 vdd.n3376 185
R16393 vdd.n3375 vdd.n3374 185
R16394 vdd.n3373 vdd.n3372 185
R16395 vdd.n3371 vdd.n3370 185
R16396 vdd.n3369 vdd.n3368 185
R16397 vdd.n3367 vdd.n691 185
R16398 vdd.n3497 vdd.n3496 185
R16399 vdd.n3496 vdd.n3495 185
R16400 vdd.n3624 vdd.n3623 185
R16401 vdd.n618 vdd.n425 185
R16402 vdd.n617 vdd.n616 185
R16403 vdd.n615 vdd.n614 185
R16404 vdd.n613 vdd.n430 185
R16405 vdd.n609 vdd.n608 185
R16406 vdd.n607 vdd.n606 185
R16407 vdd.n605 vdd.n604 185
R16408 vdd.n603 vdd.n432 185
R16409 vdd.n599 vdd.n598 185
R16410 vdd.n597 vdd.n596 185
R16411 vdd.n595 vdd.n594 185
R16412 vdd.n593 vdd.n434 185
R16413 vdd.n589 vdd.n588 185
R16414 vdd.n587 vdd.n586 185
R16415 vdd.n585 vdd.n584 185
R16416 vdd.n583 vdd.n436 185
R16417 vdd.n579 vdd.n578 185
R16418 vdd.n577 vdd.n576 185
R16419 vdd.n575 vdd.n574 185
R16420 vdd.n573 vdd.n438 185
R16421 vdd.n569 vdd.n568 185
R16422 vdd.n567 vdd.n566 185
R16423 vdd.n565 vdd.n564 185
R16424 vdd.n563 vdd.n442 185
R16425 vdd.n559 vdd.n558 185
R16426 vdd.n557 vdd.n556 185
R16427 vdd.n555 vdd.n554 185
R16428 vdd.n553 vdd.n444 185
R16429 vdd.n549 vdd.n548 185
R16430 vdd.n547 vdd.n546 185
R16431 vdd.n545 vdd.n544 185
R16432 vdd.n543 vdd.n446 185
R16433 vdd.n539 vdd.n538 185
R16434 vdd.n537 vdd.n536 185
R16435 vdd.n535 vdd.n534 185
R16436 vdd.n533 vdd.n448 185
R16437 vdd.n529 vdd.n528 185
R16438 vdd.n527 vdd.n526 185
R16439 vdd.n525 vdd.n524 185
R16440 vdd.n523 vdd.n450 185
R16441 vdd.n519 vdd.n518 185
R16442 vdd.n517 vdd.n516 185
R16443 vdd.n515 vdd.n514 185
R16444 vdd.n513 vdd.n454 185
R16445 vdd.n509 vdd.n508 185
R16446 vdd.n507 vdd.n506 185
R16447 vdd.n505 vdd.n504 185
R16448 vdd.n503 vdd.n456 185
R16449 vdd.n499 vdd.n498 185
R16450 vdd.n497 vdd.n496 185
R16451 vdd.n495 vdd.n494 185
R16452 vdd.n493 vdd.n458 185
R16453 vdd.n489 vdd.n488 185
R16454 vdd.n487 vdd.n486 185
R16455 vdd.n485 vdd.n484 185
R16456 vdd.n483 vdd.n460 185
R16457 vdd.n479 vdd.n478 185
R16458 vdd.n477 vdd.n476 185
R16459 vdd.n475 vdd.n474 185
R16460 vdd.n473 vdd.n462 185
R16461 vdd.n469 vdd.n468 185
R16462 vdd.n467 vdd.n466 185
R16463 vdd.n465 vdd.n392 185
R16464 vdd.n3620 vdd.n393 185
R16465 vdd.n3627 vdd.n393 185
R16466 vdd.n3619 vdd.n3618 185
R16467 vdd.n3618 vdd.n386 185
R16468 vdd.n3617 vdd.n385 185
R16469 vdd.n3633 vdd.n385 185
R16470 vdd.n621 vdd.n384 185
R16471 vdd.n3634 vdd.n384 185
R16472 vdd.n3613 vdd.n383 185
R16473 vdd.n3635 vdd.n383 185
R16474 vdd.n3612 vdd.n3611 185
R16475 vdd.n3611 vdd.n375 185
R16476 vdd.n3610 vdd.n374 185
R16477 vdd.n3641 vdd.n374 185
R16478 vdd.n623 vdd.n373 185
R16479 vdd.n3642 vdd.n373 185
R16480 vdd.n3606 vdd.n372 185
R16481 vdd.n3643 vdd.n372 185
R16482 vdd.n3605 vdd.n3604 185
R16483 vdd.n3604 vdd.n3603 185
R16484 vdd.n3602 vdd.n364 185
R16485 vdd.n3649 vdd.n364 185
R16486 vdd.n625 vdd.n363 185
R16487 vdd.n3650 vdd.n363 185
R16488 vdd.n3598 vdd.n362 185
R16489 vdd.n3651 vdd.n362 185
R16490 vdd.n3597 vdd.n3596 185
R16491 vdd.n3596 vdd.n361 185
R16492 vdd.n3595 vdd.n353 185
R16493 vdd.n3657 vdd.n353 185
R16494 vdd.n627 vdd.n352 185
R16495 vdd.n3658 vdd.n352 185
R16496 vdd.n3591 vdd.n351 185
R16497 vdd.n3659 vdd.n351 185
R16498 vdd.n3590 vdd.n3589 185
R16499 vdd.n3589 vdd.n344 185
R16500 vdd.n3588 vdd.n343 185
R16501 vdd.n3665 vdd.n343 185
R16502 vdd.n629 vdd.n342 185
R16503 vdd.n3666 vdd.n342 185
R16504 vdd.n3584 vdd.n341 185
R16505 vdd.n3667 vdd.n341 185
R16506 vdd.n3583 vdd.n3582 185
R16507 vdd.n3582 vdd.n340 185
R16508 vdd.n3581 vdd.n631 185
R16509 vdd.n3581 vdd.n3580 185
R16510 vdd.n3569 vdd.n632 185
R16511 vdd.n633 vdd.n632 185
R16512 vdd.n3571 vdd.n3570 185
R16513 vdd.n3572 vdd.n3571 185
R16514 vdd.n640 vdd.n639 185
R16515 vdd.n644 vdd.n639 185
R16516 vdd.n3563 vdd.n3562 185
R16517 vdd.n3562 vdd.n3561 185
R16518 vdd.n643 vdd.n642 185
R16519 vdd.n3552 vdd.n643 185
R16520 vdd.n3551 vdd.n3550 185
R16521 vdd.n3553 vdd.n3551 185
R16522 vdd.n651 vdd.n650 185
R16523 vdd.n656 vdd.n650 185
R16524 vdd.n3546 vdd.n3545 185
R16525 vdd.n3545 vdd.n3544 185
R16526 vdd.n654 vdd.n653 185
R16527 vdd.n655 vdd.n654 185
R16528 vdd.n3535 vdd.n3534 185
R16529 vdd.n3536 vdd.n3535 185
R16530 vdd.n664 vdd.n663 185
R16531 vdd.n663 vdd.n662 185
R16532 vdd.n3530 vdd.n3529 185
R16533 vdd.n3529 vdd.n3528 185
R16534 vdd.n667 vdd.n666 185
R16535 vdd.n3519 vdd.n667 185
R16536 vdd.n3518 vdd.n3517 185
R16537 vdd.n3520 vdd.n3518 185
R16538 vdd.n674 vdd.n673 185
R16539 vdd.n679 vdd.n673 185
R16540 vdd.n3513 vdd.n3512 185
R16541 vdd.n3512 vdd.n3511 185
R16542 vdd.n677 vdd.n676 185
R16543 vdd.n678 vdd.n677 185
R16544 vdd.n3502 vdd.n3501 185
R16545 vdd.n3503 vdd.n3502 185
R16546 vdd.n686 vdd.n685 185
R16547 vdd.n723 vdd.n685 185
R16548 vdd.n3091 vdd.n3090 185
R16549 vdd.n962 vdd.n961 185
R16550 vdd.n3087 vdd.n3086 185
R16551 vdd.n3088 vdd.n3087 185
R16552 vdd.n3085 vdd.n2819 185
R16553 vdd.n3084 vdd.n3083 185
R16554 vdd.n3082 vdd.n3081 185
R16555 vdd.n3080 vdd.n3079 185
R16556 vdd.n3078 vdd.n3077 185
R16557 vdd.n3076 vdd.n3075 185
R16558 vdd.n3074 vdd.n3073 185
R16559 vdd.n3072 vdd.n3071 185
R16560 vdd.n3070 vdd.n3069 185
R16561 vdd.n3068 vdd.n3067 185
R16562 vdd.n3066 vdd.n3065 185
R16563 vdd.n3064 vdd.n3063 185
R16564 vdd.n3062 vdd.n3061 185
R16565 vdd.n3060 vdd.n3059 185
R16566 vdd.n3058 vdd.n3057 185
R16567 vdd.n3056 vdd.n3055 185
R16568 vdd.n3054 vdd.n3053 185
R16569 vdd.n3052 vdd.n3051 185
R16570 vdd.n3050 vdd.n3049 185
R16571 vdd.n3048 vdd.n3047 185
R16572 vdd.n3046 vdd.n3045 185
R16573 vdd.n3044 vdd.n3043 185
R16574 vdd.n3042 vdd.n3041 185
R16575 vdd.n3040 vdd.n3039 185
R16576 vdd.n3038 vdd.n3037 185
R16577 vdd.n3036 vdd.n3035 185
R16578 vdd.n3034 vdd.n3033 185
R16579 vdd.n3032 vdd.n3031 185
R16580 vdd.n3030 vdd.n3029 185
R16581 vdd.n3027 vdd.n3026 185
R16582 vdd.n3025 vdd.n3024 185
R16583 vdd.n3023 vdd.n3022 185
R16584 vdd.n3267 vdd.n3266 185
R16585 vdd.n3269 vdd.n834 185
R16586 vdd.n3271 vdd.n3270 185
R16587 vdd.n3273 vdd.n831 185
R16588 vdd.n3275 vdd.n3274 185
R16589 vdd.n3277 vdd.n829 185
R16590 vdd.n3279 vdd.n3278 185
R16591 vdd.n3280 vdd.n828 185
R16592 vdd.n3282 vdd.n3281 185
R16593 vdd.n3284 vdd.n826 185
R16594 vdd.n3286 vdd.n3285 185
R16595 vdd.n3287 vdd.n825 185
R16596 vdd.n3289 vdd.n3288 185
R16597 vdd.n3291 vdd.n823 185
R16598 vdd.n3293 vdd.n3292 185
R16599 vdd.n3294 vdd.n822 185
R16600 vdd.n3296 vdd.n3295 185
R16601 vdd.n3298 vdd.n731 185
R16602 vdd.n3300 vdd.n3299 185
R16603 vdd.n3302 vdd.n820 185
R16604 vdd.n3304 vdd.n3303 185
R16605 vdd.n3305 vdd.n819 185
R16606 vdd.n3307 vdd.n3306 185
R16607 vdd.n3309 vdd.n817 185
R16608 vdd.n3311 vdd.n3310 185
R16609 vdd.n3312 vdd.n816 185
R16610 vdd.n3314 vdd.n3313 185
R16611 vdd.n3316 vdd.n814 185
R16612 vdd.n3318 vdd.n3317 185
R16613 vdd.n3319 vdd.n813 185
R16614 vdd.n3321 vdd.n3320 185
R16615 vdd.n3323 vdd.n812 185
R16616 vdd.n3324 vdd.n811 185
R16617 vdd.n3327 vdd.n3326 185
R16618 vdd.n3328 vdd.n809 185
R16619 vdd.n809 vdd.n692 185
R16620 vdd.n3265 vdd.n806 185
R16621 vdd.n3331 vdd.n806 185
R16622 vdd.n3264 vdd.n3263 185
R16623 vdd.n3263 vdd.n805 185
R16624 vdd.n3262 vdd.n836 185
R16625 vdd.n3262 vdd.n3261 185
R16626 vdd.n2905 vdd.n837 185
R16627 vdd.n846 vdd.n837 185
R16628 vdd.n2906 vdd.n844 185
R16629 vdd.n3255 vdd.n844 185
R16630 vdd.n2908 vdd.n2907 185
R16631 vdd.n2907 vdd.n843 185
R16632 vdd.n2909 vdd.n852 185
R16633 vdd.n3204 vdd.n852 185
R16634 vdd.n2911 vdd.n2910 185
R16635 vdd.n2910 vdd.n851 185
R16636 vdd.n2912 vdd.n857 185
R16637 vdd.n3198 vdd.n857 185
R16638 vdd.n2914 vdd.n2913 185
R16639 vdd.n2913 vdd.n864 185
R16640 vdd.n2915 vdd.n862 185
R16641 vdd.n3192 vdd.n862 185
R16642 vdd.n2917 vdd.n2916 185
R16643 vdd.n2916 vdd.n870 185
R16644 vdd.n2918 vdd.n868 185
R16645 vdd.n3186 vdd.n868 185
R16646 vdd.n2920 vdd.n2919 185
R16647 vdd.n2919 vdd.n877 185
R16648 vdd.n2921 vdd.n875 185
R16649 vdd.n3180 vdd.n875 185
R16650 vdd.n2923 vdd.n2922 185
R16651 vdd.n2922 vdd.n874 185
R16652 vdd.n2924 vdd.n882 185
R16653 vdd.n3174 vdd.n882 185
R16654 vdd.n2926 vdd.n2925 185
R16655 vdd.n2925 vdd.n881 185
R16656 vdd.n2927 vdd.n888 185
R16657 vdd.n3168 vdd.n888 185
R16658 vdd.n2929 vdd.n2928 185
R16659 vdd.n2928 vdd.n887 185
R16660 vdd.n2930 vdd.n893 185
R16661 vdd.n3162 vdd.n893 185
R16662 vdd.n2932 vdd.n2931 185
R16663 vdd.n2931 vdd.n901 185
R16664 vdd.n2933 vdd.n899 185
R16665 vdd.n3156 vdd.n899 185
R16666 vdd.n2935 vdd.n2934 185
R16667 vdd.n2934 vdd.n908 185
R16668 vdd.n2936 vdd.n906 185
R16669 vdd.n3150 vdd.n906 185
R16670 vdd.n2938 vdd.n2937 185
R16671 vdd.n2937 vdd.n905 185
R16672 vdd.n2939 vdd.n913 185
R16673 vdd.n3143 vdd.n913 185
R16674 vdd.n2941 vdd.n2940 185
R16675 vdd.n2940 vdd.n912 185
R16676 vdd.n2942 vdd.n918 185
R16677 vdd.n3137 vdd.n918 185
R16678 vdd.n2944 vdd.n2943 185
R16679 vdd.n2943 vdd.n925 185
R16680 vdd.n2945 vdd.n923 185
R16681 vdd.n3131 vdd.n923 185
R16682 vdd.n2947 vdd.n2946 185
R16683 vdd.n2946 vdd.n931 185
R16684 vdd.n2948 vdd.n929 185
R16685 vdd.n3125 vdd.n929 185
R16686 vdd.n3000 vdd.n2999 185
R16687 vdd.n2999 vdd.n2998 185
R16688 vdd.n3001 vdd.n935 185
R16689 vdd.n3119 vdd.n935 185
R16690 vdd.n3003 vdd.n3002 185
R16691 vdd.n3004 vdd.n3003 185
R16692 vdd.n2904 vdd.n941 185
R16693 vdd.n3113 vdd.n941 185
R16694 vdd.n2903 vdd.n2902 185
R16695 vdd.n2902 vdd.n940 185
R16696 vdd.n2901 vdd.n947 185
R16697 vdd.n3107 vdd.n947 185
R16698 vdd.n2900 vdd.n2899 185
R16699 vdd.n2899 vdd.n946 185
R16700 vdd.n2822 vdd.n952 185
R16701 vdd.n3101 vdd.n952 185
R16702 vdd.n3018 vdd.n3017 185
R16703 vdd.n3017 vdd.n3016 185
R16704 vdd.n3019 vdd.n958 185
R16705 vdd.n3095 vdd.n958 185
R16706 vdd.n3021 vdd.n3020 185
R16707 vdd.n3021 vdd.n957 185
R16708 vdd.n3092 vdd.n960 185
R16709 vdd.n960 vdd.n957 185
R16710 vdd.n3094 vdd.n3093 185
R16711 vdd.n3095 vdd.n3094 185
R16712 vdd.n951 vdd.n950 185
R16713 vdd.n3016 vdd.n951 185
R16714 vdd.n3103 vdd.n3102 185
R16715 vdd.n3102 vdd.n3101 185
R16716 vdd.n3104 vdd.n949 185
R16717 vdd.n949 vdd.n946 185
R16718 vdd.n3106 vdd.n3105 185
R16719 vdd.n3107 vdd.n3106 185
R16720 vdd.n939 vdd.n938 185
R16721 vdd.n940 vdd.n939 185
R16722 vdd.n3115 vdd.n3114 185
R16723 vdd.n3114 vdd.n3113 185
R16724 vdd.n3116 vdd.n937 185
R16725 vdd.n3004 vdd.n937 185
R16726 vdd.n3118 vdd.n3117 185
R16727 vdd.n3119 vdd.n3118 185
R16728 vdd.n928 vdd.n927 185
R16729 vdd.n2998 vdd.n928 185
R16730 vdd.n3127 vdd.n3126 185
R16731 vdd.n3126 vdd.n3125 185
R16732 vdd.n3128 vdd.n926 185
R16733 vdd.n931 vdd.n926 185
R16734 vdd.n3130 vdd.n3129 185
R16735 vdd.n3131 vdd.n3130 185
R16736 vdd.n917 vdd.n916 185
R16737 vdd.n925 vdd.n917 185
R16738 vdd.n3139 vdd.n3138 185
R16739 vdd.n3138 vdd.n3137 185
R16740 vdd.n3140 vdd.n915 185
R16741 vdd.n915 vdd.n912 185
R16742 vdd.n3142 vdd.n3141 185
R16743 vdd.n3143 vdd.n3142 185
R16744 vdd.n904 vdd.n903 185
R16745 vdd.n905 vdd.n904 185
R16746 vdd.n3152 vdd.n3151 185
R16747 vdd.n3151 vdd.n3150 185
R16748 vdd.n3153 vdd.n902 185
R16749 vdd.n908 vdd.n902 185
R16750 vdd.n3155 vdd.n3154 185
R16751 vdd.n3156 vdd.n3155 185
R16752 vdd.n892 vdd.n891 185
R16753 vdd.n901 vdd.n892 185
R16754 vdd.n3164 vdd.n3163 185
R16755 vdd.n3163 vdd.n3162 185
R16756 vdd.n3165 vdd.n890 185
R16757 vdd.n890 vdd.n887 185
R16758 vdd.n3167 vdd.n3166 185
R16759 vdd.n3168 vdd.n3167 185
R16760 vdd.n880 vdd.n879 185
R16761 vdd.n881 vdd.n880 185
R16762 vdd.n3176 vdd.n3175 185
R16763 vdd.n3175 vdd.n3174 185
R16764 vdd.n3177 vdd.n878 185
R16765 vdd.n878 vdd.n874 185
R16766 vdd.n3179 vdd.n3178 185
R16767 vdd.n3180 vdd.n3179 185
R16768 vdd.n867 vdd.n866 185
R16769 vdd.n877 vdd.n867 185
R16770 vdd.n3188 vdd.n3187 185
R16771 vdd.n3187 vdd.n3186 185
R16772 vdd.n3189 vdd.n865 185
R16773 vdd.n870 vdd.n865 185
R16774 vdd.n3191 vdd.n3190 185
R16775 vdd.n3192 vdd.n3191 185
R16776 vdd.n856 vdd.n855 185
R16777 vdd.n864 vdd.n856 185
R16778 vdd.n3200 vdd.n3199 185
R16779 vdd.n3199 vdd.n3198 185
R16780 vdd.n3201 vdd.n854 185
R16781 vdd.n854 vdd.n851 185
R16782 vdd.n3203 vdd.n3202 185
R16783 vdd.n3204 vdd.n3203 185
R16784 vdd.n842 vdd.n841 185
R16785 vdd.n843 vdd.n842 185
R16786 vdd.n3257 vdd.n3256 185
R16787 vdd.n3256 vdd.n3255 185
R16788 vdd.n3258 vdd.n840 185
R16789 vdd.n846 vdd.n840 185
R16790 vdd.n3260 vdd.n3259 185
R16791 vdd.n3261 vdd.n3260 185
R16792 vdd.n810 vdd.n808 185
R16793 vdd.n808 vdd.n805 185
R16794 vdd.n3330 vdd.n3329 185
R16795 vdd.n3331 vdd.n3330 185
R16796 vdd.n2711 vdd.n2710 185
R16797 vdd.n2712 vdd.n2711 185
R16798 vdd.n1009 vdd.n1007 185
R16799 vdd.n1007 vdd.n1005 185
R16800 vdd.n2626 vdd.n1016 185
R16801 vdd.n2637 vdd.n1016 185
R16802 vdd.n2627 vdd.n1025 185
R16803 vdd.n1399 vdd.n1025 185
R16804 vdd.n2629 vdd.n2628 185
R16805 vdd.n2630 vdd.n2629 185
R16806 vdd.n2625 vdd.n1024 185
R16807 vdd.n1024 vdd.n1021 185
R16808 vdd.n2624 vdd.n2623 185
R16809 vdd.n2623 vdd.n2622 185
R16810 vdd.n1027 vdd.n1026 185
R16811 vdd.n1028 vdd.n1027 185
R16812 vdd.n2615 vdd.n2614 185
R16813 vdd.n2616 vdd.n2615 185
R16814 vdd.n2613 vdd.n1036 185
R16815 vdd.n1425 vdd.n1036 185
R16816 vdd.n2612 vdd.n2611 185
R16817 vdd.n2611 vdd.n2610 185
R16818 vdd.n1038 vdd.n1037 185
R16819 vdd.n1046 vdd.n1038 185
R16820 vdd.n2603 vdd.n2602 185
R16821 vdd.n2604 vdd.n2603 185
R16822 vdd.n2601 vdd.n1047 185
R16823 vdd.n1052 vdd.n1047 185
R16824 vdd.n2600 vdd.n2599 185
R16825 vdd.n2599 vdd.n2598 185
R16826 vdd.n1049 vdd.n1048 185
R16827 vdd.n1437 vdd.n1049 185
R16828 vdd.n2591 vdd.n2590 185
R16829 vdd.n2592 vdd.n2591 185
R16830 vdd.n2589 vdd.n1059 185
R16831 vdd.n1059 vdd.n1056 185
R16832 vdd.n2588 vdd.n2587 185
R16833 vdd.n2587 vdd.n2586 185
R16834 vdd.n1061 vdd.n1060 185
R16835 vdd.n1062 vdd.n1061 185
R16836 vdd.n2579 vdd.n2578 185
R16837 vdd.n2580 vdd.n2579 185
R16838 vdd.n2576 vdd.n1070 185
R16839 vdd.n1076 vdd.n1070 185
R16840 vdd.n2575 vdd.n2574 185
R16841 vdd.n2574 vdd.n2573 185
R16842 vdd.n1073 vdd.n1072 185
R16843 vdd.n1083 vdd.n1073 185
R16844 vdd.n2566 vdd.n2565 185
R16845 vdd.n2567 vdd.n2566 185
R16846 vdd.n2564 vdd.n1084 185
R16847 vdd.n1084 vdd.n1080 185
R16848 vdd.n2563 vdd.n2562 185
R16849 vdd.n2562 vdd.n2561 185
R16850 vdd.n1086 vdd.n1085 185
R16851 vdd.n1087 vdd.n1086 185
R16852 vdd.n2554 vdd.n2553 185
R16853 vdd.n2555 vdd.n2554 185
R16854 vdd.n2552 vdd.n1096 185
R16855 vdd.n1096 vdd.n1093 185
R16856 vdd.n2551 vdd.n2550 185
R16857 vdd.n2550 vdd.n2549 185
R16858 vdd.n1098 vdd.n1097 185
R16859 vdd.n1106 vdd.n1098 185
R16860 vdd.n2542 vdd.n2541 185
R16861 vdd.n2543 vdd.n2542 185
R16862 vdd.n2540 vdd.n1107 185
R16863 vdd.n1112 vdd.n1107 185
R16864 vdd.n2539 vdd.n2538 185
R16865 vdd.n2538 vdd.n2537 185
R16866 vdd.n1109 vdd.n1108 185
R16867 vdd.n1119 vdd.n1109 185
R16868 vdd.n2530 vdd.n2529 185
R16869 vdd.n2531 vdd.n2530 185
R16870 vdd.n2528 vdd.n1120 185
R16871 vdd.n1120 vdd.n1116 185
R16872 vdd.n2527 vdd.n2526 185
R16873 vdd.n2526 vdd.n2525 185
R16874 vdd.n1122 vdd.n1121 185
R16875 vdd.n1123 vdd.n1122 185
R16876 vdd.n2518 vdd.n2517 185
R16877 vdd.n2519 vdd.n2518 185
R16878 vdd.n2516 vdd.n1131 185
R16879 vdd.n1137 vdd.n1131 185
R16880 vdd.n2515 vdd.n2514 185
R16881 vdd.n2514 vdd.n2513 185
R16882 vdd.n1133 vdd.n1132 185
R16883 vdd.n1134 vdd.n1133 185
R16884 vdd.n2642 vdd.n980 185
R16885 vdd.n2784 vdd.n980 185
R16886 vdd.n2644 vdd.n2643 185
R16887 vdd.n2646 vdd.n2645 185
R16888 vdd.n2648 vdd.n2647 185
R16889 vdd.n2650 vdd.n2649 185
R16890 vdd.n2652 vdd.n2651 185
R16891 vdd.n2654 vdd.n2653 185
R16892 vdd.n2656 vdd.n2655 185
R16893 vdd.n2658 vdd.n2657 185
R16894 vdd.n2660 vdd.n2659 185
R16895 vdd.n2662 vdd.n2661 185
R16896 vdd.n2664 vdd.n2663 185
R16897 vdd.n2666 vdd.n2665 185
R16898 vdd.n2668 vdd.n2667 185
R16899 vdd.n2670 vdd.n2669 185
R16900 vdd.n2672 vdd.n2671 185
R16901 vdd.n2674 vdd.n2673 185
R16902 vdd.n2676 vdd.n2675 185
R16903 vdd.n2678 vdd.n2677 185
R16904 vdd.n2680 vdd.n2679 185
R16905 vdd.n2682 vdd.n2681 185
R16906 vdd.n2684 vdd.n2683 185
R16907 vdd.n2686 vdd.n2685 185
R16908 vdd.n2688 vdd.n2687 185
R16909 vdd.n2690 vdd.n2689 185
R16910 vdd.n2692 vdd.n2691 185
R16911 vdd.n2694 vdd.n2693 185
R16912 vdd.n2696 vdd.n2695 185
R16913 vdd.n2698 vdd.n2697 185
R16914 vdd.n2700 vdd.n2699 185
R16915 vdd.n2702 vdd.n2701 185
R16916 vdd.n2704 vdd.n2703 185
R16917 vdd.n2706 vdd.n2705 185
R16918 vdd.n2708 vdd.n2707 185
R16919 vdd.n2709 vdd.n1008 185
R16920 vdd.n2641 vdd.n1006 185
R16921 vdd.n2712 vdd.n1006 185
R16922 vdd.n2640 vdd.n2639 185
R16923 vdd.n2639 vdd.n1005 185
R16924 vdd.n2638 vdd.n1013 185
R16925 vdd.n2638 vdd.n2637 185
R16926 vdd.n1415 vdd.n1014 185
R16927 vdd.n1399 vdd.n1014 185
R16928 vdd.n1416 vdd.n1023 185
R16929 vdd.n2630 vdd.n1023 185
R16930 vdd.n1418 vdd.n1417 185
R16931 vdd.n1417 vdd.n1021 185
R16932 vdd.n1419 vdd.n1030 185
R16933 vdd.n2622 vdd.n1030 185
R16934 vdd.n1421 vdd.n1420 185
R16935 vdd.n1420 vdd.n1028 185
R16936 vdd.n1422 vdd.n1035 185
R16937 vdd.n2616 vdd.n1035 185
R16938 vdd.n1424 vdd.n1423 185
R16939 vdd.n1425 vdd.n1424 185
R16940 vdd.n1414 vdd.n1040 185
R16941 vdd.n2610 vdd.n1040 185
R16942 vdd.n1413 vdd.n1412 185
R16943 vdd.n1412 vdd.n1046 185
R16944 vdd.n1411 vdd.n1045 185
R16945 vdd.n2604 vdd.n1045 185
R16946 vdd.n1410 vdd.n1409 185
R16947 vdd.n1409 vdd.n1052 185
R16948 vdd.n1318 vdd.n1051 185
R16949 vdd.n2598 vdd.n1051 185
R16950 vdd.n1439 vdd.n1438 185
R16951 vdd.n1438 vdd.n1437 185
R16952 vdd.n1440 vdd.n1058 185
R16953 vdd.n2592 vdd.n1058 185
R16954 vdd.n1442 vdd.n1441 185
R16955 vdd.n1441 vdd.n1056 185
R16956 vdd.n1443 vdd.n1064 185
R16957 vdd.n2586 vdd.n1064 185
R16958 vdd.n1445 vdd.n1444 185
R16959 vdd.n1444 vdd.n1062 185
R16960 vdd.n1446 vdd.n1069 185
R16961 vdd.n2580 vdd.n1069 185
R16962 vdd.n1448 vdd.n1447 185
R16963 vdd.n1447 vdd.n1076 185
R16964 vdd.n1449 vdd.n1075 185
R16965 vdd.n2573 vdd.n1075 185
R16966 vdd.n1451 vdd.n1450 185
R16967 vdd.n1450 vdd.n1083 185
R16968 vdd.n1452 vdd.n1082 185
R16969 vdd.n2567 vdd.n1082 185
R16970 vdd.n1454 vdd.n1453 185
R16971 vdd.n1453 vdd.n1080 185
R16972 vdd.n1455 vdd.n1089 185
R16973 vdd.n2561 vdd.n1089 185
R16974 vdd.n1457 vdd.n1456 185
R16975 vdd.n1456 vdd.n1087 185
R16976 vdd.n1458 vdd.n1095 185
R16977 vdd.n2555 vdd.n1095 185
R16978 vdd.n1460 vdd.n1459 185
R16979 vdd.n1459 vdd.n1093 185
R16980 vdd.n1461 vdd.n1100 185
R16981 vdd.n2549 vdd.n1100 185
R16982 vdd.n1463 vdd.n1462 185
R16983 vdd.n1462 vdd.n1106 185
R16984 vdd.n1464 vdd.n1105 185
R16985 vdd.n2543 vdd.n1105 185
R16986 vdd.n1466 vdd.n1465 185
R16987 vdd.n1465 vdd.n1112 185
R16988 vdd.n1467 vdd.n1111 185
R16989 vdd.n2537 vdd.n1111 185
R16990 vdd.n1469 vdd.n1468 185
R16991 vdd.n1468 vdd.n1119 185
R16992 vdd.n1470 vdd.n1118 185
R16993 vdd.n2531 vdd.n1118 185
R16994 vdd.n1472 vdd.n1471 185
R16995 vdd.n1471 vdd.n1116 185
R16996 vdd.n1473 vdd.n1125 185
R16997 vdd.n2525 vdd.n1125 185
R16998 vdd.n1475 vdd.n1474 185
R16999 vdd.n1474 vdd.n1123 185
R17000 vdd.n1476 vdd.n1130 185
R17001 vdd.n2519 vdd.n1130 185
R17002 vdd.n1478 vdd.n1477 185
R17003 vdd.n1477 vdd.n1137 185
R17004 vdd.n1479 vdd.n1136 185
R17005 vdd.n2513 vdd.n1136 185
R17006 vdd.n1481 vdd.n1480 185
R17007 vdd.n1480 vdd.n1134 185
R17008 vdd.n1281 vdd.n1280 185
R17009 vdd.n1283 vdd.n1282 185
R17010 vdd.n1285 vdd.n1284 185
R17011 vdd.n1287 vdd.n1286 185
R17012 vdd.n1289 vdd.n1288 185
R17013 vdd.n1291 vdd.n1290 185
R17014 vdd.n1293 vdd.n1292 185
R17015 vdd.n1295 vdd.n1294 185
R17016 vdd.n1297 vdd.n1296 185
R17017 vdd.n1299 vdd.n1298 185
R17018 vdd.n1301 vdd.n1300 185
R17019 vdd.n1303 vdd.n1302 185
R17020 vdd.n1305 vdd.n1304 185
R17021 vdd.n1307 vdd.n1306 185
R17022 vdd.n1309 vdd.n1308 185
R17023 vdd.n1311 vdd.n1310 185
R17024 vdd.n1313 vdd.n1312 185
R17025 vdd.n1515 vdd.n1314 185
R17026 vdd.n1514 vdd.n1513 185
R17027 vdd.n1512 vdd.n1511 185
R17028 vdd.n1510 vdd.n1509 185
R17029 vdd.n1508 vdd.n1507 185
R17030 vdd.n1506 vdd.n1505 185
R17031 vdd.n1504 vdd.n1503 185
R17032 vdd.n1502 vdd.n1501 185
R17033 vdd.n1500 vdd.n1499 185
R17034 vdd.n1498 vdd.n1497 185
R17035 vdd.n1496 vdd.n1495 185
R17036 vdd.n1494 vdd.n1493 185
R17037 vdd.n1492 vdd.n1491 185
R17038 vdd.n1490 vdd.n1489 185
R17039 vdd.n1488 vdd.n1487 185
R17040 vdd.n1486 vdd.n1485 185
R17041 vdd.n1484 vdd.n1483 185
R17042 vdd.n1482 vdd.n1175 185
R17043 vdd.n2506 vdd.n1175 185
R17044 vdd.n327 vdd.n326 171.744
R17045 vdd.n326 vdd.n325 171.744
R17046 vdd.n325 vdd.n294 171.744
R17047 vdd.n318 vdd.n294 171.744
R17048 vdd.n318 vdd.n317 171.744
R17049 vdd.n317 vdd.n299 171.744
R17050 vdd.n310 vdd.n299 171.744
R17051 vdd.n310 vdd.n309 171.744
R17052 vdd.n309 vdd.n303 171.744
R17053 vdd.n268 vdd.n267 171.744
R17054 vdd.n267 vdd.n266 171.744
R17055 vdd.n266 vdd.n235 171.744
R17056 vdd.n259 vdd.n235 171.744
R17057 vdd.n259 vdd.n258 171.744
R17058 vdd.n258 vdd.n240 171.744
R17059 vdd.n251 vdd.n240 171.744
R17060 vdd.n251 vdd.n250 171.744
R17061 vdd.n250 vdd.n244 171.744
R17062 vdd.n225 vdd.n224 171.744
R17063 vdd.n224 vdd.n223 171.744
R17064 vdd.n223 vdd.n192 171.744
R17065 vdd.n216 vdd.n192 171.744
R17066 vdd.n216 vdd.n215 171.744
R17067 vdd.n215 vdd.n197 171.744
R17068 vdd.n208 vdd.n197 171.744
R17069 vdd.n208 vdd.n207 171.744
R17070 vdd.n207 vdd.n201 171.744
R17071 vdd.n166 vdd.n165 171.744
R17072 vdd.n165 vdd.n164 171.744
R17073 vdd.n164 vdd.n133 171.744
R17074 vdd.n157 vdd.n133 171.744
R17075 vdd.n157 vdd.n156 171.744
R17076 vdd.n156 vdd.n138 171.744
R17077 vdd.n149 vdd.n138 171.744
R17078 vdd.n149 vdd.n148 171.744
R17079 vdd.n148 vdd.n142 171.744
R17080 vdd.n124 vdd.n123 171.744
R17081 vdd.n123 vdd.n122 171.744
R17082 vdd.n122 vdd.n91 171.744
R17083 vdd.n115 vdd.n91 171.744
R17084 vdd.n115 vdd.n114 171.744
R17085 vdd.n114 vdd.n96 171.744
R17086 vdd.n107 vdd.n96 171.744
R17087 vdd.n107 vdd.n106 171.744
R17088 vdd.n106 vdd.n100 171.744
R17089 vdd.n65 vdd.n64 171.744
R17090 vdd.n64 vdd.n63 171.744
R17091 vdd.n63 vdd.n32 171.744
R17092 vdd.n56 vdd.n32 171.744
R17093 vdd.n56 vdd.n55 171.744
R17094 vdd.n55 vdd.n37 171.744
R17095 vdd.n48 vdd.n37 171.744
R17096 vdd.n48 vdd.n47 171.744
R17097 vdd.n47 vdd.n41 171.744
R17098 vdd.n2201 vdd.n2200 171.744
R17099 vdd.n2200 vdd.n2199 171.744
R17100 vdd.n2199 vdd.n2168 171.744
R17101 vdd.n2192 vdd.n2168 171.744
R17102 vdd.n2192 vdd.n2191 171.744
R17103 vdd.n2191 vdd.n2173 171.744
R17104 vdd.n2184 vdd.n2173 171.744
R17105 vdd.n2184 vdd.n2183 171.744
R17106 vdd.n2183 vdd.n2177 171.744
R17107 vdd.n2260 vdd.n2259 171.744
R17108 vdd.n2259 vdd.n2258 171.744
R17109 vdd.n2258 vdd.n2227 171.744
R17110 vdd.n2251 vdd.n2227 171.744
R17111 vdd.n2251 vdd.n2250 171.744
R17112 vdd.n2250 vdd.n2232 171.744
R17113 vdd.n2243 vdd.n2232 171.744
R17114 vdd.n2243 vdd.n2242 171.744
R17115 vdd.n2242 vdd.n2236 171.744
R17116 vdd.n2099 vdd.n2098 171.744
R17117 vdd.n2098 vdd.n2097 171.744
R17118 vdd.n2097 vdd.n2066 171.744
R17119 vdd.n2090 vdd.n2066 171.744
R17120 vdd.n2090 vdd.n2089 171.744
R17121 vdd.n2089 vdd.n2071 171.744
R17122 vdd.n2082 vdd.n2071 171.744
R17123 vdd.n2082 vdd.n2081 171.744
R17124 vdd.n2081 vdd.n2075 171.744
R17125 vdd.n2158 vdd.n2157 171.744
R17126 vdd.n2157 vdd.n2156 171.744
R17127 vdd.n2156 vdd.n2125 171.744
R17128 vdd.n2149 vdd.n2125 171.744
R17129 vdd.n2149 vdd.n2148 171.744
R17130 vdd.n2148 vdd.n2130 171.744
R17131 vdd.n2141 vdd.n2130 171.744
R17132 vdd.n2141 vdd.n2140 171.744
R17133 vdd.n2140 vdd.n2134 171.744
R17134 vdd.n1998 vdd.n1997 171.744
R17135 vdd.n1997 vdd.n1996 171.744
R17136 vdd.n1996 vdd.n1965 171.744
R17137 vdd.n1989 vdd.n1965 171.744
R17138 vdd.n1989 vdd.n1988 171.744
R17139 vdd.n1988 vdd.n1970 171.744
R17140 vdd.n1981 vdd.n1970 171.744
R17141 vdd.n1981 vdd.n1980 171.744
R17142 vdd.n1980 vdd.n1974 171.744
R17143 vdd.n2057 vdd.n2056 171.744
R17144 vdd.n2056 vdd.n2055 171.744
R17145 vdd.n2055 vdd.n2024 171.744
R17146 vdd.n2048 vdd.n2024 171.744
R17147 vdd.n2048 vdd.n2047 171.744
R17148 vdd.n2047 vdd.n2029 171.744
R17149 vdd.n2040 vdd.n2029 171.744
R17150 vdd.n2040 vdd.n2039 171.744
R17151 vdd.n2039 vdd.n2033 171.744
R17152 vdd.n468 vdd.n467 146.341
R17153 vdd.n474 vdd.n473 146.341
R17154 vdd.n478 vdd.n477 146.341
R17155 vdd.n484 vdd.n483 146.341
R17156 vdd.n488 vdd.n487 146.341
R17157 vdd.n494 vdd.n493 146.341
R17158 vdd.n498 vdd.n497 146.341
R17159 vdd.n504 vdd.n503 146.341
R17160 vdd.n508 vdd.n507 146.341
R17161 vdd.n514 vdd.n513 146.341
R17162 vdd.n518 vdd.n517 146.341
R17163 vdd.n524 vdd.n523 146.341
R17164 vdd.n528 vdd.n527 146.341
R17165 vdd.n534 vdd.n533 146.341
R17166 vdd.n538 vdd.n537 146.341
R17167 vdd.n544 vdd.n543 146.341
R17168 vdd.n548 vdd.n547 146.341
R17169 vdd.n554 vdd.n553 146.341
R17170 vdd.n558 vdd.n557 146.341
R17171 vdd.n564 vdd.n563 146.341
R17172 vdd.n568 vdd.n567 146.341
R17173 vdd.n574 vdd.n573 146.341
R17174 vdd.n578 vdd.n577 146.341
R17175 vdd.n584 vdd.n583 146.341
R17176 vdd.n588 vdd.n587 146.341
R17177 vdd.n594 vdd.n593 146.341
R17178 vdd.n598 vdd.n597 146.341
R17179 vdd.n604 vdd.n603 146.341
R17180 vdd.n608 vdd.n607 146.341
R17181 vdd.n614 vdd.n613 146.341
R17182 vdd.n616 vdd.n425 146.341
R17183 vdd.n3502 vdd.n685 146.341
R17184 vdd.n3502 vdd.n677 146.341
R17185 vdd.n3512 vdd.n677 146.341
R17186 vdd.n3512 vdd.n673 146.341
R17187 vdd.n3518 vdd.n673 146.341
R17188 vdd.n3518 vdd.n667 146.341
R17189 vdd.n3529 vdd.n667 146.341
R17190 vdd.n3529 vdd.n663 146.341
R17191 vdd.n3535 vdd.n663 146.341
R17192 vdd.n3535 vdd.n654 146.341
R17193 vdd.n3545 vdd.n654 146.341
R17194 vdd.n3545 vdd.n650 146.341
R17195 vdd.n3551 vdd.n650 146.341
R17196 vdd.n3551 vdd.n643 146.341
R17197 vdd.n3562 vdd.n643 146.341
R17198 vdd.n3562 vdd.n639 146.341
R17199 vdd.n3571 vdd.n639 146.341
R17200 vdd.n3571 vdd.n632 146.341
R17201 vdd.n3581 vdd.n632 146.341
R17202 vdd.n3582 vdd.n3581 146.341
R17203 vdd.n3582 vdd.n341 146.341
R17204 vdd.n342 vdd.n341 146.341
R17205 vdd.n343 vdd.n342 146.341
R17206 vdd.n3589 vdd.n343 146.341
R17207 vdd.n3589 vdd.n351 146.341
R17208 vdd.n352 vdd.n351 146.341
R17209 vdd.n353 vdd.n352 146.341
R17210 vdd.n3596 vdd.n353 146.341
R17211 vdd.n3596 vdd.n362 146.341
R17212 vdd.n363 vdd.n362 146.341
R17213 vdd.n364 vdd.n363 146.341
R17214 vdd.n3604 vdd.n364 146.341
R17215 vdd.n3604 vdd.n372 146.341
R17216 vdd.n373 vdd.n372 146.341
R17217 vdd.n374 vdd.n373 146.341
R17218 vdd.n3611 vdd.n374 146.341
R17219 vdd.n3611 vdd.n383 146.341
R17220 vdd.n384 vdd.n383 146.341
R17221 vdd.n385 vdd.n384 146.341
R17222 vdd.n3618 vdd.n385 146.341
R17223 vdd.n3618 vdd.n393 146.341
R17224 vdd.n725 vdd.n724 146.341
R17225 vdd.n728 vdd.n724 146.341
R17226 vdd.n734 vdd.n733 146.341
R17227 vdd.n3484 vdd.n3483 146.341
R17228 vdd.n3480 vdd.n3479 146.341
R17229 vdd.n3476 vdd.n3475 146.341
R17230 vdd.n3472 vdd.n3471 146.341
R17231 vdd.n3468 vdd.n3467 146.341
R17232 vdd.n3464 vdd.n3463 146.341
R17233 vdd.n3460 vdd.n3459 146.341
R17234 vdd.n3451 vdd.n3450 146.341
R17235 vdd.n3448 vdd.n3447 146.341
R17236 vdd.n3444 vdd.n3443 146.341
R17237 vdd.n3440 vdd.n3439 146.341
R17238 vdd.n3436 vdd.n3435 146.341
R17239 vdd.n3432 vdd.n3431 146.341
R17240 vdd.n3428 vdd.n3427 146.341
R17241 vdd.n3424 vdd.n3423 146.341
R17242 vdd.n3420 vdd.n3419 146.341
R17243 vdd.n3416 vdd.n3415 146.341
R17244 vdd.n3412 vdd.n3411 146.341
R17245 vdd.n3405 vdd.n3404 146.341
R17246 vdd.n3402 vdd.n3401 146.341
R17247 vdd.n3398 vdd.n3397 146.341
R17248 vdd.n3394 vdd.n3393 146.341
R17249 vdd.n3390 vdd.n3389 146.341
R17250 vdd.n3386 vdd.n3385 146.341
R17251 vdd.n3382 vdd.n3381 146.341
R17252 vdd.n3378 vdd.n3377 146.341
R17253 vdd.n3374 vdd.n3373 146.341
R17254 vdd.n3370 vdd.n3369 146.341
R17255 vdd.n3496 vdd.n691 146.341
R17256 vdd.n3504 vdd.n684 146.341
R17257 vdd.n3504 vdd.n680 146.341
R17258 vdd.n3510 vdd.n680 146.341
R17259 vdd.n3510 vdd.n672 146.341
R17260 vdd.n3521 vdd.n672 146.341
R17261 vdd.n3521 vdd.n668 146.341
R17262 vdd.n3527 vdd.n668 146.341
R17263 vdd.n3527 vdd.n661 146.341
R17264 vdd.n3537 vdd.n661 146.341
R17265 vdd.n3537 vdd.n657 146.341
R17266 vdd.n3543 vdd.n657 146.341
R17267 vdd.n3543 vdd.n649 146.341
R17268 vdd.n3554 vdd.n649 146.341
R17269 vdd.n3554 vdd.n645 146.341
R17270 vdd.n3560 vdd.n645 146.341
R17271 vdd.n3560 vdd.n638 146.341
R17272 vdd.n3573 vdd.n638 146.341
R17273 vdd.n3573 vdd.n634 146.341
R17274 vdd.n3579 vdd.n634 146.341
R17275 vdd.n3579 vdd.n338 146.341
R17276 vdd.n3668 vdd.n338 146.341
R17277 vdd.n3668 vdd.n339 146.341
R17278 vdd.n3664 vdd.n339 146.341
R17279 vdd.n3664 vdd.n345 146.341
R17280 vdd.n3660 vdd.n345 146.341
R17281 vdd.n3660 vdd.n350 146.341
R17282 vdd.n3656 vdd.n350 146.341
R17283 vdd.n3656 vdd.n354 146.341
R17284 vdd.n3652 vdd.n354 146.341
R17285 vdd.n3652 vdd.n360 146.341
R17286 vdd.n3648 vdd.n360 146.341
R17287 vdd.n3648 vdd.n365 146.341
R17288 vdd.n3644 vdd.n365 146.341
R17289 vdd.n3644 vdd.n371 146.341
R17290 vdd.n3640 vdd.n371 146.341
R17291 vdd.n3640 vdd.n376 146.341
R17292 vdd.n3636 vdd.n376 146.341
R17293 vdd.n3636 vdd.n382 146.341
R17294 vdd.n3632 vdd.n382 146.341
R17295 vdd.n3632 vdd.n387 146.341
R17296 vdd.n3628 vdd.n387 146.341
R17297 vdd.n2471 vdd.n2470 146.341
R17298 vdd.n2468 vdd.n2465 146.341
R17299 vdd.n2463 vdd.n1185 146.341
R17300 vdd.n2459 vdd.n2458 146.341
R17301 vdd.n2456 vdd.n1189 146.341
R17302 vdd.n2452 vdd.n2451 146.341
R17303 vdd.n2449 vdd.n1196 146.341
R17304 vdd.n2445 vdd.n2444 146.341
R17305 vdd.n2442 vdd.n1203 146.341
R17306 vdd.n1214 vdd.n1211 146.341
R17307 vdd.n2434 vdd.n2433 146.341
R17308 vdd.n2431 vdd.n1216 146.341
R17309 vdd.n2427 vdd.n2426 146.341
R17310 vdd.n2424 vdd.n1222 146.341
R17311 vdd.n2420 vdd.n2419 146.341
R17312 vdd.n2417 vdd.n1229 146.341
R17313 vdd.n2413 vdd.n2412 146.341
R17314 vdd.n2410 vdd.n1236 146.341
R17315 vdd.n2406 vdd.n2405 146.341
R17316 vdd.n2403 vdd.n1243 146.341
R17317 vdd.n1254 vdd.n1251 146.341
R17318 vdd.n2395 vdd.n2394 146.341
R17319 vdd.n2392 vdd.n1256 146.341
R17320 vdd.n2388 vdd.n2387 146.341
R17321 vdd.n2385 vdd.n1262 146.341
R17322 vdd.n2381 vdd.n2380 146.341
R17323 vdd.n2378 vdd.n1269 146.341
R17324 vdd.n2374 vdd.n2373 146.341
R17325 vdd.n2371 vdd.n1276 146.341
R17326 vdd.n1522 vdd.n1520 146.341
R17327 vdd.n1525 vdd.n1524 146.341
R17328 vdd.n1883 vdd.n1643 146.341
R17329 vdd.n1883 vdd.n1639 146.341
R17330 vdd.n1889 vdd.n1639 146.341
R17331 vdd.n1889 vdd.n1631 146.341
R17332 vdd.n1900 vdd.n1631 146.341
R17333 vdd.n1900 vdd.n1627 146.341
R17334 vdd.n1906 vdd.n1627 146.341
R17335 vdd.n1906 vdd.n1621 146.341
R17336 vdd.n1917 vdd.n1621 146.341
R17337 vdd.n1917 vdd.n1617 146.341
R17338 vdd.n1923 vdd.n1617 146.341
R17339 vdd.n1923 vdd.n1608 146.341
R17340 vdd.n1933 vdd.n1608 146.341
R17341 vdd.n1933 vdd.n1604 146.341
R17342 vdd.n1939 vdd.n1604 146.341
R17343 vdd.n1939 vdd.n1597 146.341
R17344 vdd.n1950 vdd.n1597 146.341
R17345 vdd.n1950 vdd.n1593 146.341
R17346 vdd.n1956 vdd.n1593 146.341
R17347 vdd.n1956 vdd.n1586 146.341
R17348 vdd.n2273 vdd.n1586 146.341
R17349 vdd.n2273 vdd.n1582 146.341
R17350 vdd.n2279 vdd.n1582 146.341
R17351 vdd.n2279 vdd.n1574 146.341
R17352 vdd.n2290 vdd.n1574 146.341
R17353 vdd.n2290 vdd.n1570 146.341
R17354 vdd.n2296 vdd.n1570 146.341
R17355 vdd.n2296 vdd.n1564 146.341
R17356 vdd.n2307 vdd.n1564 146.341
R17357 vdd.n2307 vdd.n1560 146.341
R17358 vdd.n2313 vdd.n1560 146.341
R17359 vdd.n2313 vdd.n1551 146.341
R17360 vdd.n2323 vdd.n1551 146.341
R17361 vdd.n2323 vdd.n1547 146.341
R17362 vdd.n2329 vdd.n1547 146.341
R17363 vdd.n2329 vdd.n1541 146.341
R17364 vdd.n2340 vdd.n1541 146.341
R17365 vdd.n2340 vdd.n1536 146.341
R17366 vdd.n2348 vdd.n1536 146.341
R17367 vdd.n2348 vdd.n1527 146.341
R17368 vdd.n2359 vdd.n1527 146.341
R17369 vdd.n1872 vdd.n1648 146.341
R17370 vdd.n1872 vdd.n1681 146.341
R17371 vdd.n1685 vdd.n1684 146.341
R17372 vdd.n1687 vdd.n1686 146.341
R17373 vdd.n1691 vdd.n1690 146.341
R17374 vdd.n1693 vdd.n1692 146.341
R17375 vdd.n1697 vdd.n1696 146.341
R17376 vdd.n1699 vdd.n1698 146.341
R17377 vdd.n1703 vdd.n1702 146.341
R17378 vdd.n1705 vdd.n1704 146.341
R17379 vdd.n1711 vdd.n1710 146.341
R17380 vdd.n1713 vdd.n1712 146.341
R17381 vdd.n1717 vdd.n1716 146.341
R17382 vdd.n1719 vdd.n1718 146.341
R17383 vdd.n1723 vdd.n1722 146.341
R17384 vdd.n1725 vdd.n1724 146.341
R17385 vdd.n1729 vdd.n1728 146.341
R17386 vdd.n1731 vdd.n1730 146.341
R17387 vdd.n1735 vdd.n1734 146.341
R17388 vdd.n1737 vdd.n1736 146.341
R17389 vdd.n1809 vdd.n1740 146.341
R17390 vdd.n1742 vdd.n1741 146.341
R17391 vdd.n1746 vdd.n1745 146.341
R17392 vdd.n1748 vdd.n1747 146.341
R17393 vdd.n1752 vdd.n1751 146.341
R17394 vdd.n1754 vdd.n1753 146.341
R17395 vdd.n1758 vdd.n1757 146.341
R17396 vdd.n1760 vdd.n1759 146.341
R17397 vdd.n1764 vdd.n1763 146.341
R17398 vdd.n1766 vdd.n1765 146.341
R17399 vdd.n1770 vdd.n1769 146.341
R17400 vdd.n1771 vdd.n1679 146.341
R17401 vdd.n1881 vdd.n1644 146.341
R17402 vdd.n1881 vdd.n1637 146.341
R17403 vdd.n1892 vdd.n1637 146.341
R17404 vdd.n1892 vdd.n1633 146.341
R17405 vdd.n1898 vdd.n1633 146.341
R17406 vdd.n1898 vdd.n1626 146.341
R17407 vdd.n1909 vdd.n1626 146.341
R17408 vdd.n1909 vdd.n1622 146.341
R17409 vdd.n1915 vdd.n1622 146.341
R17410 vdd.n1915 vdd.n1615 146.341
R17411 vdd.n1925 vdd.n1615 146.341
R17412 vdd.n1925 vdd.n1611 146.341
R17413 vdd.n1931 vdd.n1611 146.341
R17414 vdd.n1931 vdd.n1603 146.341
R17415 vdd.n1942 vdd.n1603 146.341
R17416 vdd.n1942 vdd.n1599 146.341
R17417 vdd.n1948 vdd.n1599 146.341
R17418 vdd.n1948 vdd.n1592 146.341
R17419 vdd.n1958 vdd.n1592 146.341
R17420 vdd.n1958 vdd.n1588 146.341
R17421 vdd.n2271 vdd.n1588 146.341
R17422 vdd.n2271 vdd.n1580 146.341
R17423 vdd.n2282 vdd.n1580 146.341
R17424 vdd.n2282 vdd.n1576 146.341
R17425 vdd.n2288 vdd.n1576 146.341
R17426 vdd.n2288 vdd.n1569 146.341
R17427 vdd.n2299 vdd.n1569 146.341
R17428 vdd.n2299 vdd.n1565 146.341
R17429 vdd.n2305 vdd.n1565 146.341
R17430 vdd.n2305 vdd.n1558 146.341
R17431 vdd.n2315 vdd.n1558 146.341
R17432 vdd.n2315 vdd.n1554 146.341
R17433 vdd.n2321 vdd.n1554 146.341
R17434 vdd.n2321 vdd.n1546 146.341
R17435 vdd.n2332 vdd.n1546 146.341
R17436 vdd.n2332 vdd.n1542 146.341
R17437 vdd.n2338 vdd.n1542 146.341
R17438 vdd.n2338 vdd.n1534 146.341
R17439 vdd.n2351 vdd.n1534 146.341
R17440 vdd.n2351 vdd.n1529 146.341
R17441 vdd.n2357 vdd.n1529 146.341
R17442 vdd.n1315 vdd.t90 127.284
R17443 vdd.n1010 vdd.t130 127.284
R17444 vdd.n1319 vdd.t127 127.284
R17445 vdd.n1001 vdd.t151 127.284
R17446 vdd.n896 vdd.t114 127.284
R17447 vdd.n896 vdd.t115 127.284
R17448 vdd.n2823 vdd.t145 127.284
R17449 vdd.n832 vdd.t106 127.284
R17450 vdd.n2820 vdd.t138 127.284
R17451 vdd.n799 vdd.t85 127.284
R17452 vdd.n1071 vdd.t141 127.284
R17453 vdd.n1071 vdd.t142 127.284
R17454 vdd.n22 vdd.n20 117.314
R17455 vdd.n17 vdd.n15 117.314
R17456 vdd.n27 vdd.n26 116.927
R17457 vdd.n24 vdd.n23 116.927
R17458 vdd.n22 vdd.n21 116.927
R17459 vdd.n17 vdd.n16 116.927
R17460 vdd.n19 vdd.n18 116.927
R17461 vdd.n27 vdd.n25 116.927
R17462 vdd.n1316 vdd.t89 111.188
R17463 vdd.n1011 vdd.t131 111.188
R17464 vdd.n1320 vdd.t126 111.188
R17465 vdd.n1002 vdd.t152 111.188
R17466 vdd.n2824 vdd.t144 111.188
R17467 vdd.n833 vdd.t107 111.188
R17468 vdd.n2821 vdd.t137 111.188
R17469 vdd.n800 vdd.t86 111.188
R17470 vdd.n3094 vdd.n960 99.5127
R17471 vdd.n3094 vdd.n951 99.5127
R17472 vdd.n3102 vdd.n951 99.5127
R17473 vdd.n3102 vdd.n949 99.5127
R17474 vdd.n3106 vdd.n949 99.5127
R17475 vdd.n3106 vdd.n939 99.5127
R17476 vdd.n3114 vdd.n939 99.5127
R17477 vdd.n3114 vdd.n937 99.5127
R17478 vdd.n3118 vdd.n937 99.5127
R17479 vdd.n3118 vdd.n928 99.5127
R17480 vdd.n3126 vdd.n928 99.5127
R17481 vdd.n3126 vdd.n926 99.5127
R17482 vdd.n3130 vdd.n926 99.5127
R17483 vdd.n3130 vdd.n917 99.5127
R17484 vdd.n3138 vdd.n917 99.5127
R17485 vdd.n3138 vdd.n915 99.5127
R17486 vdd.n3142 vdd.n915 99.5127
R17487 vdd.n3142 vdd.n904 99.5127
R17488 vdd.n3151 vdd.n904 99.5127
R17489 vdd.n3151 vdd.n902 99.5127
R17490 vdd.n3155 vdd.n902 99.5127
R17491 vdd.n3155 vdd.n892 99.5127
R17492 vdd.n3163 vdd.n892 99.5127
R17493 vdd.n3163 vdd.n890 99.5127
R17494 vdd.n3167 vdd.n890 99.5127
R17495 vdd.n3167 vdd.n880 99.5127
R17496 vdd.n3175 vdd.n880 99.5127
R17497 vdd.n3175 vdd.n878 99.5127
R17498 vdd.n3179 vdd.n878 99.5127
R17499 vdd.n3179 vdd.n867 99.5127
R17500 vdd.n3187 vdd.n867 99.5127
R17501 vdd.n3187 vdd.n865 99.5127
R17502 vdd.n3191 vdd.n865 99.5127
R17503 vdd.n3191 vdd.n856 99.5127
R17504 vdd.n3199 vdd.n856 99.5127
R17505 vdd.n3199 vdd.n854 99.5127
R17506 vdd.n3203 vdd.n854 99.5127
R17507 vdd.n3203 vdd.n842 99.5127
R17508 vdd.n3256 vdd.n842 99.5127
R17509 vdd.n3256 vdd.n840 99.5127
R17510 vdd.n3260 vdd.n840 99.5127
R17511 vdd.n3260 vdd.n808 99.5127
R17512 vdd.n3330 vdd.n808 99.5127
R17513 vdd.n3326 vdd.n809 99.5127
R17514 vdd.n3324 vdd.n3323 99.5127
R17515 vdd.n3321 vdd.n813 99.5127
R17516 vdd.n3317 vdd.n3316 99.5127
R17517 vdd.n3314 vdd.n816 99.5127
R17518 vdd.n3310 vdd.n3309 99.5127
R17519 vdd.n3307 vdd.n819 99.5127
R17520 vdd.n3303 vdd.n3302 99.5127
R17521 vdd.n3300 vdd.n3298 99.5127
R17522 vdd.n3296 vdd.n822 99.5127
R17523 vdd.n3292 vdd.n3291 99.5127
R17524 vdd.n3289 vdd.n825 99.5127
R17525 vdd.n3285 vdd.n3284 99.5127
R17526 vdd.n3282 vdd.n828 99.5127
R17527 vdd.n3278 vdd.n3277 99.5127
R17528 vdd.n3275 vdd.n831 99.5127
R17529 vdd.n3270 vdd.n3269 99.5127
R17530 vdd.n3021 vdd.n958 99.5127
R17531 vdd.n3017 vdd.n958 99.5127
R17532 vdd.n3017 vdd.n952 99.5127
R17533 vdd.n2899 vdd.n952 99.5127
R17534 vdd.n2899 vdd.n947 99.5127
R17535 vdd.n2902 vdd.n947 99.5127
R17536 vdd.n2902 vdd.n941 99.5127
R17537 vdd.n3003 vdd.n941 99.5127
R17538 vdd.n3003 vdd.n935 99.5127
R17539 vdd.n2999 vdd.n935 99.5127
R17540 vdd.n2999 vdd.n929 99.5127
R17541 vdd.n2946 vdd.n929 99.5127
R17542 vdd.n2946 vdd.n923 99.5127
R17543 vdd.n2943 vdd.n923 99.5127
R17544 vdd.n2943 vdd.n918 99.5127
R17545 vdd.n2940 vdd.n918 99.5127
R17546 vdd.n2940 vdd.n913 99.5127
R17547 vdd.n2937 vdd.n913 99.5127
R17548 vdd.n2937 vdd.n906 99.5127
R17549 vdd.n2934 vdd.n906 99.5127
R17550 vdd.n2934 vdd.n899 99.5127
R17551 vdd.n2931 vdd.n899 99.5127
R17552 vdd.n2931 vdd.n893 99.5127
R17553 vdd.n2928 vdd.n893 99.5127
R17554 vdd.n2928 vdd.n888 99.5127
R17555 vdd.n2925 vdd.n888 99.5127
R17556 vdd.n2925 vdd.n882 99.5127
R17557 vdd.n2922 vdd.n882 99.5127
R17558 vdd.n2922 vdd.n875 99.5127
R17559 vdd.n2919 vdd.n875 99.5127
R17560 vdd.n2919 vdd.n868 99.5127
R17561 vdd.n2916 vdd.n868 99.5127
R17562 vdd.n2916 vdd.n862 99.5127
R17563 vdd.n2913 vdd.n862 99.5127
R17564 vdd.n2913 vdd.n857 99.5127
R17565 vdd.n2910 vdd.n857 99.5127
R17566 vdd.n2910 vdd.n852 99.5127
R17567 vdd.n2907 vdd.n852 99.5127
R17568 vdd.n2907 vdd.n844 99.5127
R17569 vdd.n844 vdd.n837 99.5127
R17570 vdd.n3262 vdd.n837 99.5127
R17571 vdd.n3263 vdd.n3262 99.5127
R17572 vdd.n3263 vdd.n806 99.5127
R17573 vdd.n3087 vdd.n962 99.5127
R17574 vdd.n3087 vdd.n2819 99.5127
R17575 vdd.n3083 vdd.n3082 99.5127
R17576 vdd.n3079 vdd.n3078 99.5127
R17577 vdd.n3075 vdd.n3074 99.5127
R17578 vdd.n3071 vdd.n3070 99.5127
R17579 vdd.n3067 vdd.n3066 99.5127
R17580 vdd.n3063 vdd.n3062 99.5127
R17581 vdd.n3059 vdd.n3058 99.5127
R17582 vdd.n3055 vdd.n3054 99.5127
R17583 vdd.n3051 vdd.n3050 99.5127
R17584 vdd.n3047 vdd.n3046 99.5127
R17585 vdd.n3043 vdd.n3042 99.5127
R17586 vdd.n3039 vdd.n3038 99.5127
R17587 vdd.n3035 vdd.n3034 99.5127
R17588 vdd.n3031 vdd.n3030 99.5127
R17589 vdd.n3026 vdd.n3025 99.5127
R17590 vdd.n2783 vdd.n999 99.5127
R17591 vdd.n2779 vdd.n2778 99.5127
R17592 vdd.n2775 vdd.n2774 99.5127
R17593 vdd.n2771 vdd.n2770 99.5127
R17594 vdd.n2767 vdd.n2766 99.5127
R17595 vdd.n2763 vdd.n2762 99.5127
R17596 vdd.n2759 vdd.n2758 99.5127
R17597 vdd.n2755 vdd.n2754 99.5127
R17598 vdd.n2751 vdd.n2750 99.5127
R17599 vdd.n2747 vdd.n2746 99.5127
R17600 vdd.n2743 vdd.n2742 99.5127
R17601 vdd.n2739 vdd.n2738 99.5127
R17602 vdd.n2735 vdd.n2734 99.5127
R17603 vdd.n2731 vdd.n2730 99.5127
R17604 vdd.n2727 vdd.n2726 99.5127
R17605 vdd.n2723 vdd.n2722 99.5127
R17606 vdd.n2718 vdd.n2717 99.5127
R17607 vdd.n1355 vdd.n1135 99.5127
R17608 vdd.n1358 vdd.n1135 99.5127
R17609 vdd.n1358 vdd.n1129 99.5127
R17610 vdd.n1361 vdd.n1129 99.5127
R17611 vdd.n1361 vdd.n1124 99.5127
R17612 vdd.n1364 vdd.n1124 99.5127
R17613 vdd.n1364 vdd.n1117 99.5127
R17614 vdd.n1367 vdd.n1117 99.5127
R17615 vdd.n1367 vdd.n1110 99.5127
R17616 vdd.n1370 vdd.n1110 99.5127
R17617 vdd.n1370 vdd.n1104 99.5127
R17618 vdd.n1373 vdd.n1104 99.5127
R17619 vdd.n1373 vdd.n1099 99.5127
R17620 vdd.n1376 vdd.n1099 99.5127
R17621 vdd.n1376 vdd.n1094 99.5127
R17622 vdd.n1379 vdd.n1094 99.5127
R17623 vdd.n1379 vdd.n1088 99.5127
R17624 vdd.n1382 vdd.n1088 99.5127
R17625 vdd.n1382 vdd.n1081 99.5127
R17626 vdd.n1385 vdd.n1081 99.5127
R17627 vdd.n1385 vdd.n1074 99.5127
R17628 vdd.n1388 vdd.n1074 99.5127
R17629 vdd.n1388 vdd.n1068 99.5127
R17630 vdd.n1391 vdd.n1068 99.5127
R17631 vdd.n1391 vdd.n1063 99.5127
R17632 vdd.n1394 vdd.n1063 99.5127
R17633 vdd.n1394 vdd.n1057 99.5127
R17634 vdd.n1436 vdd.n1057 99.5127
R17635 vdd.n1436 vdd.n1050 99.5127
R17636 vdd.n1432 vdd.n1050 99.5127
R17637 vdd.n1432 vdd.n1044 99.5127
R17638 vdd.n1429 vdd.n1044 99.5127
R17639 vdd.n1429 vdd.n1039 99.5127
R17640 vdd.n1426 vdd.n1039 99.5127
R17641 vdd.n1426 vdd.n1034 99.5127
R17642 vdd.n1406 vdd.n1034 99.5127
R17643 vdd.n1406 vdd.n1029 99.5127
R17644 vdd.n1403 vdd.n1029 99.5127
R17645 vdd.n1403 vdd.n1022 99.5127
R17646 vdd.n1400 vdd.n1022 99.5127
R17647 vdd.n1400 vdd.n1015 99.5127
R17648 vdd.n1015 vdd.n1004 99.5127
R17649 vdd.n2713 vdd.n1004 99.5127
R17650 vdd.n2505 vdd.n1140 99.5127
R17651 vdd.n2505 vdd.n1176 99.5127
R17652 vdd.n2501 vdd.n2500 99.5127
R17653 vdd.n2497 vdd.n2496 99.5127
R17654 vdd.n2493 vdd.n2492 99.5127
R17655 vdd.n2489 vdd.n2488 99.5127
R17656 vdd.n2485 vdd.n2484 99.5127
R17657 vdd.n2481 vdd.n2480 99.5127
R17658 vdd.n2477 vdd.n2476 99.5127
R17659 vdd.n1322 vdd.n1321 99.5127
R17660 vdd.n1326 vdd.n1325 99.5127
R17661 vdd.n1330 vdd.n1329 99.5127
R17662 vdd.n1334 vdd.n1333 99.5127
R17663 vdd.n1338 vdd.n1337 99.5127
R17664 vdd.n1342 vdd.n1341 99.5127
R17665 vdd.n1346 vdd.n1345 99.5127
R17666 vdd.n1351 vdd.n1350 99.5127
R17667 vdd.n2512 vdd.n1138 99.5127
R17668 vdd.n2512 vdd.n1128 99.5127
R17669 vdd.n2520 vdd.n1128 99.5127
R17670 vdd.n2520 vdd.n1126 99.5127
R17671 vdd.n2524 vdd.n1126 99.5127
R17672 vdd.n2524 vdd.n1115 99.5127
R17673 vdd.n2532 vdd.n1115 99.5127
R17674 vdd.n2532 vdd.n1113 99.5127
R17675 vdd.n2536 vdd.n1113 99.5127
R17676 vdd.n2536 vdd.n1103 99.5127
R17677 vdd.n2544 vdd.n1103 99.5127
R17678 vdd.n2544 vdd.n1101 99.5127
R17679 vdd.n2548 vdd.n1101 99.5127
R17680 vdd.n2548 vdd.n1092 99.5127
R17681 vdd.n2556 vdd.n1092 99.5127
R17682 vdd.n2556 vdd.n1090 99.5127
R17683 vdd.n2560 vdd.n1090 99.5127
R17684 vdd.n2560 vdd.n1079 99.5127
R17685 vdd.n2568 vdd.n1079 99.5127
R17686 vdd.n2568 vdd.n1077 99.5127
R17687 vdd.n2572 vdd.n1077 99.5127
R17688 vdd.n2572 vdd.n1067 99.5127
R17689 vdd.n2581 vdd.n1067 99.5127
R17690 vdd.n2581 vdd.n1065 99.5127
R17691 vdd.n2585 vdd.n1065 99.5127
R17692 vdd.n2585 vdd.n1055 99.5127
R17693 vdd.n2593 vdd.n1055 99.5127
R17694 vdd.n2593 vdd.n1053 99.5127
R17695 vdd.n2597 vdd.n1053 99.5127
R17696 vdd.n2597 vdd.n1043 99.5127
R17697 vdd.n2605 vdd.n1043 99.5127
R17698 vdd.n2605 vdd.n1041 99.5127
R17699 vdd.n2609 vdd.n1041 99.5127
R17700 vdd.n2609 vdd.n1033 99.5127
R17701 vdd.n2617 vdd.n1033 99.5127
R17702 vdd.n2617 vdd.n1031 99.5127
R17703 vdd.n2621 vdd.n1031 99.5127
R17704 vdd.n2621 vdd.n1020 99.5127
R17705 vdd.n2631 vdd.n1020 99.5127
R17706 vdd.n2631 vdd.n1017 99.5127
R17707 vdd.n2636 vdd.n1017 99.5127
R17708 vdd.n2636 vdd.n1018 99.5127
R17709 vdd.n1018 vdd.n998 99.5127
R17710 vdd.n3246 vdd.n3245 99.5127
R17711 vdd.n3243 vdd.n3209 99.5127
R17712 vdd.n3239 vdd.n3238 99.5127
R17713 vdd.n3236 vdd.n3212 99.5127
R17714 vdd.n3232 vdd.n3231 99.5127
R17715 vdd.n3229 vdd.n3215 99.5127
R17716 vdd.n3225 vdd.n3224 99.5127
R17717 vdd.n3222 vdd.n3219 99.5127
R17718 vdd.n3363 vdd.n787 99.5127
R17719 vdd.n3361 vdd.n3360 99.5127
R17720 vdd.n3358 vdd.n789 99.5127
R17721 vdd.n3354 vdd.n3353 99.5127
R17722 vdd.n3351 vdd.n792 99.5127
R17723 vdd.n3347 vdd.n3346 99.5127
R17724 vdd.n3344 vdd.n795 99.5127
R17725 vdd.n3340 vdd.n3339 99.5127
R17726 vdd.n3337 vdd.n798 99.5127
R17727 vdd.n2895 vdd.n959 99.5127
R17728 vdd.n3015 vdd.n959 99.5127
R17729 vdd.n3015 vdd.n953 99.5127
R17730 vdd.n3011 vdd.n953 99.5127
R17731 vdd.n3011 vdd.n948 99.5127
R17732 vdd.n3008 vdd.n948 99.5127
R17733 vdd.n3008 vdd.n942 99.5127
R17734 vdd.n3005 vdd.n942 99.5127
R17735 vdd.n3005 vdd.n936 99.5127
R17736 vdd.n2997 vdd.n936 99.5127
R17737 vdd.n2997 vdd.n930 99.5127
R17738 vdd.n2993 vdd.n930 99.5127
R17739 vdd.n2993 vdd.n924 99.5127
R17740 vdd.n2990 vdd.n924 99.5127
R17741 vdd.n2990 vdd.n919 99.5127
R17742 vdd.n2987 vdd.n919 99.5127
R17743 vdd.n2987 vdd.n914 99.5127
R17744 vdd.n2984 vdd.n914 99.5127
R17745 vdd.n2984 vdd.n907 99.5127
R17746 vdd.n2981 vdd.n907 99.5127
R17747 vdd.n2981 vdd.n900 99.5127
R17748 vdd.n2978 vdd.n900 99.5127
R17749 vdd.n2978 vdd.n894 99.5127
R17750 vdd.n2975 vdd.n894 99.5127
R17751 vdd.n2975 vdd.n889 99.5127
R17752 vdd.n2972 vdd.n889 99.5127
R17753 vdd.n2972 vdd.n883 99.5127
R17754 vdd.n2969 vdd.n883 99.5127
R17755 vdd.n2969 vdd.n876 99.5127
R17756 vdd.n2966 vdd.n876 99.5127
R17757 vdd.n2966 vdd.n869 99.5127
R17758 vdd.n2963 vdd.n869 99.5127
R17759 vdd.n2963 vdd.n863 99.5127
R17760 vdd.n2960 vdd.n863 99.5127
R17761 vdd.n2960 vdd.n858 99.5127
R17762 vdd.n2957 vdd.n858 99.5127
R17763 vdd.n2957 vdd.n853 99.5127
R17764 vdd.n2954 vdd.n853 99.5127
R17765 vdd.n2954 vdd.n845 99.5127
R17766 vdd.n2951 vdd.n845 99.5127
R17767 vdd.n2951 vdd.n838 99.5127
R17768 vdd.n838 vdd.n804 99.5127
R17769 vdd.n3332 vdd.n804 99.5127
R17770 vdd.n2830 vdd.n2829 99.5127
R17771 vdd.n2834 vdd.n2833 99.5127
R17772 vdd.n2838 vdd.n2837 99.5127
R17773 vdd.n2842 vdd.n2841 99.5127
R17774 vdd.n2846 vdd.n2845 99.5127
R17775 vdd.n2850 vdd.n2849 99.5127
R17776 vdd.n2854 vdd.n2853 99.5127
R17777 vdd.n2858 vdd.n2857 99.5127
R17778 vdd.n2862 vdd.n2861 99.5127
R17779 vdd.n2866 vdd.n2865 99.5127
R17780 vdd.n2870 vdd.n2869 99.5127
R17781 vdd.n2874 vdd.n2873 99.5127
R17782 vdd.n2878 vdd.n2877 99.5127
R17783 vdd.n2882 vdd.n2881 99.5127
R17784 vdd.n2886 vdd.n2885 99.5127
R17785 vdd.n2890 vdd.n2889 99.5127
R17786 vdd.n2892 vdd.n2818 99.5127
R17787 vdd.n3096 vdd.n956 99.5127
R17788 vdd.n3096 vdd.n954 99.5127
R17789 vdd.n3100 vdd.n954 99.5127
R17790 vdd.n3100 vdd.n945 99.5127
R17791 vdd.n3108 vdd.n945 99.5127
R17792 vdd.n3108 vdd.n943 99.5127
R17793 vdd.n3112 vdd.n943 99.5127
R17794 vdd.n3112 vdd.n934 99.5127
R17795 vdd.n3120 vdd.n934 99.5127
R17796 vdd.n3120 vdd.n932 99.5127
R17797 vdd.n3124 vdd.n932 99.5127
R17798 vdd.n3124 vdd.n922 99.5127
R17799 vdd.n3132 vdd.n922 99.5127
R17800 vdd.n3132 vdd.n920 99.5127
R17801 vdd.n3136 vdd.n920 99.5127
R17802 vdd.n3136 vdd.n911 99.5127
R17803 vdd.n3144 vdd.n911 99.5127
R17804 vdd.n3144 vdd.n909 99.5127
R17805 vdd.n3149 vdd.n909 99.5127
R17806 vdd.n3149 vdd.n898 99.5127
R17807 vdd.n3157 vdd.n898 99.5127
R17808 vdd.n3157 vdd.n895 99.5127
R17809 vdd.n3161 vdd.n895 99.5127
R17810 vdd.n3161 vdd.n886 99.5127
R17811 vdd.n3169 vdd.n886 99.5127
R17812 vdd.n3169 vdd.n884 99.5127
R17813 vdd.n3173 vdd.n884 99.5127
R17814 vdd.n3173 vdd.n873 99.5127
R17815 vdd.n3181 vdd.n873 99.5127
R17816 vdd.n3181 vdd.n871 99.5127
R17817 vdd.n3185 vdd.n871 99.5127
R17818 vdd.n3185 vdd.n861 99.5127
R17819 vdd.n3193 vdd.n861 99.5127
R17820 vdd.n3193 vdd.n859 99.5127
R17821 vdd.n3197 vdd.n859 99.5127
R17822 vdd.n3197 vdd.n850 99.5127
R17823 vdd.n3205 vdd.n850 99.5127
R17824 vdd.n3205 vdd.n847 99.5127
R17825 vdd.n3254 vdd.n847 99.5127
R17826 vdd.n3254 vdd.n848 99.5127
R17827 vdd.n848 vdd.n839 99.5127
R17828 vdd.n3249 vdd.n839 99.5127
R17829 vdd.n3249 vdd.n807 99.5127
R17830 vdd.n2707 vdd.n2706 99.5127
R17831 vdd.n2703 vdd.n2702 99.5127
R17832 vdd.n2699 vdd.n2698 99.5127
R17833 vdd.n2695 vdd.n2694 99.5127
R17834 vdd.n2691 vdd.n2690 99.5127
R17835 vdd.n2687 vdd.n2686 99.5127
R17836 vdd.n2683 vdd.n2682 99.5127
R17837 vdd.n2679 vdd.n2678 99.5127
R17838 vdd.n2675 vdd.n2674 99.5127
R17839 vdd.n2671 vdd.n2670 99.5127
R17840 vdd.n2667 vdd.n2666 99.5127
R17841 vdd.n2663 vdd.n2662 99.5127
R17842 vdd.n2659 vdd.n2658 99.5127
R17843 vdd.n2655 vdd.n2654 99.5127
R17844 vdd.n2651 vdd.n2650 99.5127
R17845 vdd.n2647 vdd.n2646 99.5127
R17846 vdd.n2643 vdd.n980 99.5127
R17847 vdd.n1480 vdd.n1136 99.5127
R17848 vdd.n1477 vdd.n1136 99.5127
R17849 vdd.n1477 vdd.n1130 99.5127
R17850 vdd.n1474 vdd.n1130 99.5127
R17851 vdd.n1474 vdd.n1125 99.5127
R17852 vdd.n1471 vdd.n1125 99.5127
R17853 vdd.n1471 vdd.n1118 99.5127
R17854 vdd.n1468 vdd.n1118 99.5127
R17855 vdd.n1468 vdd.n1111 99.5127
R17856 vdd.n1465 vdd.n1111 99.5127
R17857 vdd.n1465 vdd.n1105 99.5127
R17858 vdd.n1462 vdd.n1105 99.5127
R17859 vdd.n1462 vdd.n1100 99.5127
R17860 vdd.n1459 vdd.n1100 99.5127
R17861 vdd.n1459 vdd.n1095 99.5127
R17862 vdd.n1456 vdd.n1095 99.5127
R17863 vdd.n1456 vdd.n1089 99.5127
R17864 vdd.n1453 vdd.n1089 99.5127
R17865 vdd.n1453 vdd.n1082 99.5127
R17866 vdd.n1450 vdd.n1082 99.5127
R17867 vdd.n1450 vdd.n1075 99.5127
R17868 vdd.n1447 vdd.n1075 99.5127
R17869 vdd.n1447 vdd.n1069 99.5127
R17870 vdd.n1444 vdd.n1069 99.5127
R17871 vdd.n1444 vdd.n1064 99.5127
R17872 vdd.n1441 vdd.n1064 99.5127
R17873 vdd.n1441 vdd.n1058 99.5127
R17874 vdd.n1438 vdd.n1058 99.5127
R17875 vdd.n1438 vdd.n1051 99.5127
R17876 vdd.n1409 vdd.n1051 99.5127
R17877 vdd.n1409 vdd.n1045 99.5127
R17878 vdd.n1412 vdd.n1045 99.5127
R17879 vdd.n1412 vdd.n1040 99.5127
R17880 vdd.n1424 vdd.n1040 99.5127
R17881 vdd.n1424 vdd.n1035 99.5127
R17882 vdd.n1420 vdd.n1035 99.5127
R17883 vdd.n1420 vdd.n1030 99.5127
R17884 vdd.n1417 vdd.n1030 99.5127
R17885 vdd.n1417 vdd.n1023 99.5127
R17886 vdd.n1023 vdd.n1014 99.5127
R17887 vdd.n2638 vdd.n1014 99.5127
R17888 vdd.n2639 vdd.n2638 99.5127
R17889 vdd.n2639 vdd.n1006 99.5127
R17890 vdd.n1284 vdd.n1283 99.5127
R17891 vdd.n1288 vdd.n1287 99.5127
R17892 vdd.n1292 vdd.n1291 99.5127
R17893 vdd.n1296 vdd.n1295 99.5127
R17894 vdd.n1300 vdd.n1299 99.5127
R17895 vdd.n1304 vdd.n1303 99.5127
R17896 vdd.n1308 vdd.n1307 99.5127
R17897 vdd.n1312 vdd.n1311 99.5127
R17898 vdd.n1513 vdd.n1314 99.5127
R17899 vdd.n1511 vdd.n1510 99.5127
R17900 vdd.n1507 vdd.n1506 99.5127
R17901 vdd.n1503 vdd.n1502 99.5127
R17902 vdd.n1499 vdd.n1498 99.5127
R17903 vdd.n1495 vdd.n1494 99.5127
R17904 vdd.n1491 vdd.n1490 99.5127
R17905 vdd.n1487 vdd.n1486 99.5127
R17906 vdd.n1483 vdd.n1175 99.5127
R17907 vdd.n2514 vdd.n1133 99.5127
R17908 vdd.n2514 vdd.n1131 99.5127
R17909 vdd.n2518 vdd.n1131 99.5127
R17910 vdd.n2518 vdd.n1122 99.5127
R17911 vdd.n2526 vdd.n1122 99.5127
R17912 vdd.n2526 vdd.n1120 99.5127
R17913 vdd.n2530 vdd.n1120 99.5127
R17914 vdd.n2530 vdd.n1109 99.5127
R17915 vdd.n2538 vdd.n1109 99.5127
R17916 vdd.n2538 vdd.n1107 99.5127
R17917 vdd.n2542 vdd.n1107 99.5127
R17918 vdd.n2542 vdd.n1098 99.5127
R17919 vdd.n2550 vdd.n1098 99.5127
R17920 vdd.n2550 vdd.n1096 99.5127
R17921 vdd.n2554 vdd.n1096 99.5127
R17922 vdd.n2554 vdd.n1086 99.5127
R17923 vdd.n2562 vdd.n1086 99.5127
R17924 vdd.n2562 vdd.n1084 99.5127
R17925 vdd.n2566 vdd.n1084 99.5127
R17926 vdd.n2566 vdd.n1073 99.5127
R17927 vdd.n2574 vdd.n1073 99.5127
R17928 vdd.n2574 vdd.n1070 99.5127
R17929 vdd.n2579 vdd.n1070 99.5127
R17930 vdd.n2579 vdd.n1061 99.5127
R17931 vdd.n2587 vdd.n1061 99.5127
R17932 vdd.n2587 vdd.n1059 99.5127
R17933 vdd.n2591 vdd.n1059 99.5127
R17934 vdd.n2591 vdd.n1049 99.5127
R17935 vdd.n2599 vdd.n1049 99.5127
R17936 vdd.n2599 vdd.n1047 99.5127
R17937 vdd.n2603 vdd.n1047 99.5127
R17938 vdd.n2603 vdd.n1038 99.5127
R17939 vdd.n2611 vdd.n1038 99.5127
R17940 vdd.n2611 vdd.n1036 99.5127
R17941 vdd.n2615 vdd.n1036 99.5127
R17942 vdd.n2615 vdd.n1027 99.5127
R17943 vdd.n2623 vdd.n1027 99.5127
R17944 vdd.n2623 vdd.n1024 99.5127
R17945 vdd.n2629 vdd.n1024 99.5127
R17946 vdd.n2629 vdd.n1025 99.5127
R17947 vdd.n1025 vdd.n1016 99.5127
R17948 vdd.n1016 vdd.n1007 99.5127
R17949 vdd.n2711 vdd.n1007 99.5127
R17950 vdd.n9 vdd.n7 98.9633
R17951 vdd.n2 vdd.n0 98.9633
R17952 vdd.n9 vdd.n8 98.6055
R17953 vdd.n11 vdd.n10 98.6055
R17954 vdd.n13 vdd.n12 98.6055
R17955 vdd.n6 vdd.n5 98.6055
R17956 vdd.n4 vdd.n3 98.6055
R17957 vdd.n2 vdd.n1 98.6055
R17958 vdd.t210 vdd.n303 85.8723
R17959 vdd.t65 vdd.n244 85.8723
R17960 vdd.t185 vdd.n201 85.8723
R17961 vdd.t81 vdd.n142 85.8723
R17962 vdd.t202 vdd.n100 85.8723
R17963 vdd.t32 vdd.n41 85.8723
R17964 vdd.t211 vdd.n2177 85.8723
R17965 vdd.t38 vdd.n2236 85.8723
R17966 vdd.t165 vdd.n2075 85.8723
R17967 vdd.t60 vdd.n2134 85.8723
R17968 vdd.t48 vdd.n1974 85.8723
R17969 vdd.t225 vdd.n2033 85.8723
R17970 vdd.n897 vdd.n896 78.546
R17971 vdd.n2577 vdd.n1071 78.546
R17972 vdd.n290 vdd.n289 75.1835
R17973 vdd.n288 vdd.n287 75.1835
R17974 vdd.n286 vdd.n285 75.1835
R17975 vdd.n284 vdd.n283 75.1835
R17976 vdd.n282 vdd.n281 75.1835
R17977 vdd.n280 vdd.n279 75.1835
R17978 vdd.n278 vdd.n277 75.1835
R17979 vdd.n276 vdd.n275 75.1835
R17980 vdd.n274 vdd.n273 75.1835
R17981 vdd.n188 vdd.n187 75.1835
R17982 vdd.n186 vdd.n185 75.1835
R17983 vdd.n184 vdd.n183 75.1835
R17984 vdd.n182 vdd.n181 75.1835
R17985 vdd.n180 vdd.n179 75.1835
R17986 vdd.n178 vdd.n177 75.1835
R17987 vdd.n176 vdd.n175 75.1835
R17988 vdd.n174 vdd.n173 75.1835
R17989 vdd.n172 vdd.n171 75.1835
R17990 vdd.n87 vdd.n86 75.1835
R17991 vdd.n85 vdd.n84 75.1835
R17992 vdd.n83 vdd.n82 75.1835
R17993 vdd.n81 vdd.n80 75.1835
R17994 vdd.n79 vdd.n78 75.1835
R17995 vdd.n77 vdd.n76 75.1835
R17996 vdd.n75 vdd.n74 75.1835
R17997 vdd.n73 vdd.n72 75.1835
R17998 vdd.n71 vdd.n70 75.1835
R17999 vdd.n2207 vdd.n2206 75.1835
R18000 vdd.n2209 vdd.n2208 75.1835
R18001 vdd.n2211 vdd.n2210 75.1835
R18002 vdd.n2213 vdd.n2212 75.1835
R18003 vdd.n2215 vdd.n2214 75.1835
R18004 vdd.n2217 vdd.n2216 75.1835
R18005 vdd.n2219 vdd.n2218 75.1835
R18006 vdd.n2221 vdd.n2220 75.1835
R18007 vdd.n2223 vdd.n2222 75.1835
R18008 vdd.n2105 vdd.n2104 75.1835
R18009 vdd.n2107 vdd.n2106 75.1835
R18010 vdd.n2109 vdd.n2108 75.1835
R18011 vdd.n2111 vdd.n2110 75.1835
R18012 vdd.n2113 vdd.n2112 75.1835
R18013 vdd.n2115 vdd.n2114 75.1835
R18014 vdd.n2117 vdd.n2116 75.1835
R18015 vdd.n2119 vdd.n2118 75.1835
R18016 vdd.n2121 vdd.n2120 75.1835
R18017 vdd.n2004 vdd.n2003 75.1835
R18018 vdd.n2006 vdd.n2005 75.1835
R18019 vdd.n2008 vdd.n2007 75.1835
R18020 vdd.n2010 vdd.n2009 75.1835
R18021 vdd.n2012 vdd.n2011 75.1835
R18022 vdd.n2014 vdd.n2013 75.1835
R18023 vdd.n2016 vdd.n2015 75.1835
R18024 vdd.n2018 vdd.n2017 75.1835
R18025 vdd.n2020 vdd.n2019 75.1835
R18026 vdd.n3088 vdd.n2801 72.8958
R18027 vdd.n3088 vdd.n2802 72.8958
R18028 vdd.n3088 vdd.n2803 72.8958
R18029 vdd.n3088 vdd.n2804 72.8958
R18030 vdd.n3088 vdd.n2805 72.8958
R18031 vdd.n3088 vdd.n2806 72.8958
R18032 vdd.n3088 vdd.n2807 72.8958
R18033 vdd.n3088 vdd.n2808 72.8958
R18034 vdd.n3088 vdd.n2809 72.8958
R18035 vdd.n3088 vdd.n2810 72.8958
R18036 vdd.n3088 vdd.n2811 72.8958
R18037 vdd.n3088 vdd.n2812 72.8958
R18038 vdd.n3088 vdd.n2813 72.8958
R18039 vdd.n3088 vdd.n2814 72.8958
R18040 vdd.n3088 vdd.n2815 72.8958
R18041 vdd.n3088 vdd.n2816 72.8958
R18042 vdd.n3088 vdd.n2817 72.8958
R18043 vdd.n803 vdd.n692 72.8958
R18044 vdd.n3338 vdd.n692 72.8958
R18045 vdd.n797 vdd.n692 72.8958
R18046 vdd.n3345 vdd.n692 72.8958
R18047 vdd.n794 vdd.n692 72.8958
R18048 vdd.n3352 vdd.n692 72.8958
R18049 vdd.n791 vdd.n692 72.8958
R18050 vdd.n3359 vdd.n692 72.8958
R18051 vdd.n3362 vdd.n692 72.8958
R18052 vdd.n3218 vdd.n692 72.8958
R18053 vdd.n3223 vdd.n692 72.8958
R18054 vdd.n3217 vdd.n692 72.8958
R18055 vdd.n3230 vdd.n692 72.8958
R18056 vdd.n3214 vdd.n692 72.8958
R18057 vdd.n3237 vdd.n692 72.8958
R18058 vdd.n3211 vdd.n692 72.8958
R18059 vdd.n3244 vdd.n692 72.8958
R18060 vdd.n2507 vdd.n2506 72.8958
R18061 vdd.n2506 vdd.n1142 72.8958
R18062 vdd.n2506 vdd.n1143 72.8958
R18063 vdd.n2506 vdd.n1144 72.8958
R18064 vdd.n2506 vdd.n1145 72.8958
R18065 vdd.n2506 vdd.n1146 72.8958
R18066 vdd.n2506 vdd.n1147 72.8958
R18067 vdd.n2506 vdd.n1148 72.8958
R18068 vdd.n2506 vdd.n1149 72.8958
R18069 vdd.n2506 vdd.n1150 72.8958
R18070 vdd.n2506 vdd.n1151 72.8958
R18071 vdd.n2506 vdd.n1152 72.8958
R18072 vdd.n2506 vdd.n1153 72.8958
R18073 vdd.n2506 vdd.n1154 72.8958
R18074 vdd.n2506 vdd.n1155 72.8958
R18075 vdd.n2506 vdd.n1156 72.8958
R18076 vdd.n2506 vdd.n1157 72.8958
R18077 vdd.n2784 vdd.n981 72.8958
R18078 vdd.n2784 vdd.n982 72.8958
R18079 vdd.n2784 vdd.n983 72.8958
R18080 vdd.n2784 vdd.n984 72.8958
R18081 vdd.n2784 vdd.n985 72.8958
R18082 vdd.n2784 vdd.n986 72.8958
R18083 vdd.n2784 vdd.n987 72.8958
R18084 vdd.n2784 vdd.n988 72.8958
R18085 vdd.n2784 vdd.n989 72.8958
R18086 vdd.n2784 vdd.n990 72.8958
R18087 vdd.n2784 vdd.n991 72.8958
R18088 vdd.n2784 vdd.n992 72.8958
R18089 vdd.n2784 vdd.n993 72.8958
R18090 vdd.n2784 vdd.n994 72.8958
R18091 vdd.n2784 vdd.n995 72.8958
R18092 vdd.n2784 vdd.n996 72.8958
R18093 vdd.n2784 vdd.n997 72.8958
R18094 vdd.n3089 vdd.n3088 72.8958
R18095 vdd.n3088 vdd.n2785 72.8958
R18096 vdd.n3088 vdd.n2786 72.8958
R18097 vdd.n3088 vdd.n2787 72.8958
R18098 vdd.n3088 vdd.n2788 72.8958
R18099 vdd.n3088 vdd.n2789 72.8958
R18100 vdd.n3088 vdd.n2790 72.8958
R18101 vdd.n3088 vdd.n2791 72.8958
R18102 vdd.n3088 vdd.n2792 72.8958
R18103 vdd.n3088 vdd.n2793 72.8958
R18104 vdd.n3088 vdd.n2794 72.8958
R18105 vdd.n3088 vdd.n2795 72.8958
R18106 vdd.n3088 vdd.n2796 72.8958
R18107 vdd.n3088 vdd.n2797 72.8958
R18108 vdd.n3088 vdd.n2798 72.8958
R18109 vdd.n3088 vdd.n2799 72.8958
R18110 vdd.n3088 vdd.n2800 72.8958
R18111 vdd.n3268 vdd.n692 72.8958
R18112 vdd.n835 vdd.n692 72.8958
R18113 vdd.n3276 vdd.n692 72.8958
R18114 vdd.n830 vdd.n692 72.8958
R18115 vdd.n3283 vdd.n692 72.8958
R18116 vdd.n827 vdd.n692 72.8958
R18117 vdd.n3290 vdd.n692 72.8958
R18118 vdd.n824 vdd.n692 72.8958
R18119 vdd.n3297 vdd.n692 72.8958
R18120 vdd.n3301 vdd.n692 72.8958
R18121 vdd.n821 vdd.n692 72.8958
R18122 vdd.n3308 vdd.n692 72.8958
R18123 vdd.n818 vdd.n692 72.8958
R18124 vdd.n3315 vdd.n692 72.8958
R18125 vdd.n815 vdd.n692 72.8958
R18126 vdd.n3322 vdd.n692 72.8958
R18127 vdd.n3325 vdd.n692 72.8958
R18128 vdd.n2784 vdd.n979 72.8958
R18129 vdd.n2784 vdd.n978 72.8958
R18130 vdd.n2784 vdd.n977 72.8958
R18131 vdd.n2784 vdd.n976 72.8958
R18132 vdd.n2784 vdd.n975 72.8958
R18133 vdd.n2784 vdd.n974 72.8958
R18134 vdd.n2784 vdd.n973 72.8958
R18135 vdd.n2784 vdd.n972 72.8958
R18136 vdd.n2784 vdd.n971 72.8958
R18137 vdd.n2784 vdd.n970 72.8958
R18138 vdd.n2784 vdd.n969 72.8958
R18139 vdd.n2784 vdd.n968 72.8958
R18140 vdd.n2784 vdd.n967 72.8958
R18141 vdd.n2784 vdd.n966 72.8958
R18142 vdd.n2784 vdd.n965 72.8958
R18143 vdd.n2784 vdd.n964 72.8958
R18144 vdd.n2784 vdd.n963 72.8958
R18145 vdd.n2506 vdd.n1158 72.8958
R18146 vdd.n2506 vdd.n1159 72.8958
R18147 vdd.n2506 vdd.n1160 72.8958
R18148 vdd.n2506 vdd.n1161 72.8958
R18149 vdd.n2506 vdd.n1162 72.8958
R18150 vdd.n2506 vdd.n1163 72.8958
R18151 vdd.n2506 vdd.n1164 72.8958
R18152 vdd.n2506 vdd.n1165 72.8958
R18153 vdd.n2506 vdd.n1166 72.8958
R18154 vdd.n2506 vdd.n1167 72.8958
R18155 vdd.n2506 vdd.n1168 72.8958
R18156 vdd.n2506 vdd.n1169 72.8958
R18157 vdd.n2506 vdd.n1170 72.8958
R18158 vdd.n2506 vdd.n1171 72.8958
R18159 vdd.n2506 vdd.n1172 72.8958
R18160 vdd.n2506 vdd.n1173 72.8958
R18161 vdd.n2506 vdd.n1174 72.8958
R18162 vdd.n1874 vdd.n1873 66.2847
R18163 vdd.n1873 vdd.n1649 66.2847
R18164 vdd.n1873 vdd.n1650 66.2847
R18165 vdd.n1873 vdd.n1651 66.2847
R18166 vdd.n1873 vdd.n1652 66.2847
R18167 vdd.n1873 vdd.n1653 66.2847
R18168 vdd.n1873 vdd.n1654 66.2847
R18169 vdd.n1873 vdd.n1655 66.2847
R18170 vdd.n1873 vdd.n1656 66.2847
R18171 vdd.n1873 vdd.n1657 66.2847
R18172 vdd.n1873 vdd.n1658 66.2847
R18173 vdd.n1873 vdd.n1659 66.2847
R18174 vdd.n1873 vdd.n1660 66.2847
R18175 vdd.n1873 vdd.n1661 66.2847
R18176 vdd.n1873 vdd.n1662 66.2847
R18177 vdd.n1873 vdd.n1663 66.2847
R18178 vdd.n1873 vdd.n1664 66.2847
R18179 vdd.n1873 vdd.n1665 66.2847
R18180 vdd.n1873 vdd.n1666 66.2847
R18181 vdd.n1873 vdd.n1667 66.2847
R18182 vdd.n1873 vdd.n1668 66.2847
R18183 vdd.n1873 vdd.n1669 66.2847
R18184 vdd.n1873 vdd.n1670 66.2847
R18185 vdd.n1873 vdd.n1671 66.2847
R18186 vdd.n1873 vdd.n1672 66.2847
R18187 vdd.n1873 vdd.n1673 66.2847
R18188 vdd.n1873 vdd.n1674 66.2847
R18189 vdd.n1873 vdd.n1675 66.2847
R18190 vdd.n1873 vdd.n1676 66.2847
R18191 vdd.n1873 vdd.n1677 66.2847
R18192 vdd.n1873 vdd.n1678 66.2847
R18193 vdd.n1526 vdd.n1141 66.2847
R18194 vdd.n1523 vdd.n1141 66.2847
R18195 vdd.n1519 vdd.n1141 66.2847
R18196 vdd.n2372 vdd.n1141 66.2847
R18197 vdd.n1275 vdd.n1141 66.2847
R18198 vdd.n2379 vdd.n1141 66.2847
R18199 vdd.n1268 vdd.n1141 66.2847
R18200 vdd.n2386 vdd.n1141 66.2847
R18201 vdd.n1261 vdd.n1141 66.2847
R18202 vdd.n2393 vdd.n1141 66.2847
R18203 vdd.n1255 vdd.n1141 66.2847
R18204 vdd.n1250 vdd.n1141 66.2847
R18205 vdd.n2404 vdd.n1141 66.2847
R18206 vdd.n1242 vdd.n1141 66.2847
R18207 vdd.n2411 vdd.n1141 66.2847
R18208 vdd.n1235 vdd.n1141 66.2847
R18209 vdd.n2418 vdd.n1141 66.2847
R18210 vdd.n1228 vdd.n1141 66.2847
R18211 vdd.n2425 vdd.n1141 66.2847
R18212 vdd.n1221 vdd.n1141 66.2847
R18213 vdd.n2432 vdd.n1141 66.2847
R18214 vdd.n1215 vdd.n1141 66.2847
R18215 vdd.n1210 vdd.n1141 66.2847
R18216 vdd.n2443 vdd.n1141 66.2847
R18217 vdd.n1202 vdd.n1141 66.2847
R18218 vdd.n2450 vdd.n1141 66.2847
R18219 vdd.n1195 vdd.n1141 66.2847
R18220 vdd.n2457 vdd.n1141 66.2847
R18221 vdd.n1188 vdd.n1141 66.2847
R18222 vdd.n2464 vdd.n1141 66.2847
R18223 vdd.n2469 vdd.n1141 66.2847
R18224 vdd.n1184 vdd.n1141 66.2847
R18225 vdd.n3495 vdd.n3494 66.2847
R18226 vdd.n3495 vdd.n693 66.2847
R18227 vdd.n3495 vdd.n694 66.2847
R18228 vdd.n3495 vdd.n695 66.2847
R18229 vdd.n3495 vdd.n696 66.2847
R18230 vdd.n3495 vdd.n697 66.2847
R18231 vdd.n3495 vdd.n698 66.2847
R18232 vdd.n3495 vdd.n699 66.2847
R18233 vdd.n3495 vdd.n700 66.2847
R18234 vdd.n3495 vdd.n701 66.2847
R18235 vdd.n3495 vdd.n702 66.2847
R18236 vdd.n3495 vdd.n703 66.2847
R18237 vdd.n3495 vdd.n704 66.2847
R18238 vdd.n3495 vdd.n705 66.2847
R18239 vdd.n3495 vdd.n706 66.2847
R18240 vdd.n3495 vdd.n707 66.2847
R18241 vdd.n3495 vdd.n708 66.2847
R18242 vdd.n3495 vdd.n709 66.2847
R18243 vdd.n3495 vdd.n710 66.2847
R18244 vdd.n3495 vdd.n711 66.2847
R18245 vdd.n3495 vdd.n712 66.2847
R18246 vdd.n3495 vdd.n713 66.2847
R18247 vdd.n3495 vdd.n714 66.2847
R18248 vdd.n3495 vdd.n715 66.2847
R18249 vdd.n3495 vdd.n716 66.2847
R18250 vdd.n3495 vdd.n717 66.2847
R18251 vdd.n3495 vdd.n718 66.2847
R18252 vdd.n3495 vdd.n719 66.2847
R18253 vdd.n3495 vdd.n720 66.2847
R18254 vdd.n3495 vdd.n721 66.2847
R18255 vdd.n3495 vdd.n722 66.2847
R18256 vdd.n3626 vdd.n3625 66.2847
R18257 vdd.n3626 vdd.n424 66.2847
R18258 vdd.n3626 vdd.n423 66.2847
R18259 vdd.n3626 vdd.n422 66.2847
R18260 vdd.n3626 vdd.n421 66.2847
R18261 vdd.n3626 vdd.n420 66.2847
R18262 vdd.n3626 vdd.n419 66.2847
R18263 vdd.n3626 vdd.n418 66.2847
R18264 vdd.n3626 vdd.n417 66.2847
R18265 vdd.n3626 vdd.n416 66.2847
R18266 vdd.n3626 vdd.n415 66.2847
R18267 vdd.n3626 vdd.n414 66.2847
R18268 vdd.n3626 vdd.n413 66.2847
R18269 vdd.n3626 vdd.n412 66.2847
R18270 vdd.n3626 vdd.n411 66.2847
R18271 vdd.n3626 vdd.n410 66.2847
R18272 vdd.n3626 vdd.n409 66.2847
R18273 vdd.n3626 vdd.n408 66.2847
R18274 vdd.n3626 vdd.n407 66.2847
R18275 vdd.n3626 vdd.n406 66.2847
R18276 vdd.n3626 vdd.n405 66.2847
R18277 vdd.n3626 vdd.n404 66.2847
R18278 vdd.n3626 vdd.n403 66.2847
R18279 vdd.n3626 vdd.n402 66.2847
R18280 vdd.n3626 vdd.n401 66.2847
R18281 vdd.n3626 vdd.n400 66.2847
R18282 vdd.n3626 vdd.n399 66.2847
R18283 vdd.n3626 vdd.n398 66.2847
R18284 vdd.n3626 vdd.n397 66.2847
R18285 vdd.n3626 vdd.n396 66.2847
R18286 vdd.n3626 vdd.n395 66.2847
R18287 vdd.n3626 vdd.n394 66.2847
R18288 vdd.n467 vdd.n394 52.4337
R18289 vdd.n473 vdd.n395 52.4337
R18290 vdd.n477 vdd.n396 52.4337
R18291 vdd.n483 vdd.n397 52.4337
R18292 vdd.n487 vdd.n398 52.4337
R18293 vdd.n493 vdd.n399 52.4337
R18294 vdd.n497 vdd.n400 52.4337
R18295 vdd.n503 vdd.n401 52.4337
R18296 vdd.n507 vdd.n402 52.4337
R18297 vdd.n513 vdd.n403 52.4337
R18298 vdd.n517 vdd.n404 52.4337
R18299 vdd.n523 vdd.n405 52.4337
R18300 vdd.n527 vdd.n406 52.4337
R18301 vdd.n533 vdd.n407 52.4337
R18302 vdd.n537 vdd.n408 52.4337
R18303 vdd.n543 vdd.n409 52.4337
R18304 vdd.n547 vdd.n410 52.4337
R18305 vdd.n553 vdd.n411 52.4337
R18306 vdd.n557 vdd.n412 52.4337
R18307 vdd.n563 vdd.n413 52.4337
R18308 vdd.n567 vdd.n414 52.4337
R18309 vdd.n573 vdd.n415 52.4337
R18310 vdd.n577 vdd.n416 52.4337
R18311 vdd.n583 vdd.n417 52.4337
R18312 vdd.n587 vdd.n418 52.4337
R18313 vdd.n593 vdd.n419 52.4337
R18314 vdd.n597 vdd.n420 52.4337
R18315 vdd.n603 vdd.n421 52.4337
R18316 vdd.n607 vdd.n422 52.4337
R18317 vdd.n613 vdd.n423 52.4337
R18318 vdd.n616 vdd.n424 52.4337
R18319 vdd.n3625 vdd.n3624 52.4337
R18320 vdd.n3494 vdd.n3493 52.4337
R18321 vdd.n728 vdd.n693 52.4337
R18322 vdd.n734 vdd.n694 52.4337
R18323 vdd.n3483 vdd.n695 52.4337
R18324 vdd.n3479 vdd.n696 52.4337
R18325 vdd.n3475 vdd.n697 52.4337
R18326 vdd.n3471 vdd.n698 52.4337
R18327 vdd.n3467 vdd.n699 52.4337
R18328 vdd.n3463 vdd.n700 52.4337
R18329 vdd.n3459 vdd.n701 52.4337
R18330 vdd.n3451 vdd.n702 52.4337
R18331 vdd.n3447 vdd.n703 52.4337
R18332 vdd.n3443 vdd.n704 52.4337
R18333 vdd.n3439 vdd.n705 52.4337
R18334 vdd.n3435 vdd.n706 52.4337
R18335 vdd.n3431 vdd.n707 52.4337
R18336 vdd.n3427 vdd.n708 52.4337
R18337 vdd.n3423 vdd.n709 52.4337
R18338 vdd.n3419 vdd.n710 52.4337
R18339 vdd.n3415 vdd.n711 52.4337
R18340 vdd.n3411 vdd.n712 52.4337
R18341 vdd.n3405 vdd.n713 52.4337
R18342 vdd.n3401 vdd.n714 52.4337
R18343 vdd.n3397 vdd.n715 52.4337
R18344 vdd.n3393 vdd.n716 52.4337
R18345 vdd.n3389 vdd.n717 52.4337
R18346 vdd.n3385 vdd.n718 52.4337
R18347 vdd.n3381 vdd.n719 52.4337
R18348 vdd.n3377 vdd.n720 52.4337
R18349 vdd.n3373 vdd.n721 52.4337
R18350 vdd.n3369 vdd.n722 52.4337
R18351 vdd.n2471 vdd.n1184 52.4337
R18352 vdd.n2469 vdd.n2468 52.4337
R18353 vdd.n2464 vdd.n2463 52.4337
R18354 vdd.n2459 vdd.n1188 52.4337
R18355 vdd.n2457 vdd.n2456 52.4337
R18356 vdd.n2452 vdd.n1195 52.4337
R18357 vdd.n2450 vdd.n2449 52.4337
R18358 vdd.n2445 vdd.n1202 52.4337
R18359 vdd.n2443 vdd.n2442 52.4337
R18360 vdd.n1211 vdd.n1210 52.4337
R18361 vdd.n2434 vdd.n1215 52.4337
R18362 vdd.n2432 vdd.n2431 52.4337
R18363 vdd.n2427 vdd.n1221 52.4337
R18364 vdd.n2425 vdd.n2424 52.4337
R18365 vdd.n2420 vdd.n1228 52.4337
R18366 vdd.n2418 vdd.n2417 52.4337
R18367 vdd.n2413 vdd.n1235 52.4337
R18368 vdd.n2411 vdd.n2410 52.4337
R18369 vdd.n2406 vdd.n1242 52.4337
R18370 vdd.n2404 vdd.n2403 52.4337
R18371 vdd.n1251 vdd.n1250 52.4337
R18372 vdd.n2395 vdd.n1255 52.4337
R18373 vdd.n2393 vdd.n2392 52.4337
R18374 vdd.n2388 vdd.n1261 52.4337
R18375 vdd.n2386 vdd.n2385 52.4337
R18376 vdd.n2381 vdd.n1268 52.4337
R18377 vdd.n2379 vdd.n2378 52.4337
R18378 vdd.n2374 vdd.n1275 52.4337
R18379 vdd.n2372 vdd.n2371 52.4337
R18380 vdd.n1520 vdd.n1519 52.4337
R18381 vdd.n1524 vdd.n1523 52.4337
R18382 vdd.n2360 vdd.n1526 52.4337
R18383 vdd.n1875 vdd.n1874 52.4337
R18384 vdd.n1681 vdd.n1649 52.4337
R18385 vdd.n1685 vdd.n1650 52.4337
R18386 vdd.n1687 vdd.n1651 52.4337
R18387 vdd.n1691 vdd.n1652 52.4337
R18388 vdd.n1693 vdd.n1653 52.4337
R18389 vdd.n1697 vdd.n1654 52.4337
R18390 vdd.n1699 vdd.n1655 52.4337
R18391 vdd.n1703 vdd.n1656 52.4337
R18392 vdd.n1705 vdd.n1657 52.4337
R18393 vdd.n1711 vdd.n1658 52.4337
R18394 vdd.n1713 vdd.n1659 52.4337
R18395 vdd.n1717 vdd.n1660 52.4337
R18396 vdd.n1719 vdd.n1661 52.4337
R18397 vdd.n1723 vdd.n1662 52.4337
R18398 vdd.n1725 vdd.n1663 52.4337
R18399 vdd.n1729 vdd.n1664 52.4337
R18400 vdd.n1731 vdd.n1665 52.4337
R18401 vdd.n1735 vdd.n1666 52.4337
R18402 vdd.n1737 vdd.n1667 52.4337
R18403 vdd.n1809 vdd.n1668 52.4337
R18404 vdd.n1742 vdd.n1669 52.4337
R18405 vdd.n1746 vdd.n1670 52.4337
R18406 vdd.n1748 vdd.n1671 52.4337
R18407 vdd.n1752 vdd.n1672 52.4337
R18408 vdd.n1754 vdd.n1673 52.4337
R18409 vdd.n1758 vdd.n1674 52.4337
R18410 vdd.n1760 vdd.n1675 52.4337
R18411 vdd.n1764 vdd.n1676 52.4337
R18412 vdd.n1766 vdd.n1677 52.4337
R18413 vdd.n1770 vdd.n1678 52.4337
R18414 vdd.n1874 vdd.n1648 52.4337
R18415 vdd.n1684 vdd.n1649 52.4337
R18416 vdd.n1686 vdd.n1650 52.4337
R18417 vdd.n1690 vdd.n1651 52.4337
R18418 vdd.n1692 vdd.n1652 52.4337
R18419 vdd.n1696 vdd.n1653 52.4337
R18420 vdd.n1698 vdd.n1654 52.4337
R18421 vdd.n1702 vdd.n1655 52.4337
R18422 vdd.n1704 vdd.n1656 52.4337
R18423 vdd.n1710 vdd.n1657 52.4337
R18424 vdd.n1712 vdd.n1658 52.4337
R18425 vdd.n1716 vdd.n1659 52.4337
R18426 vdd.n1718 vdd.n1660 52.4337
R18427 vdd.n1722 vdd.n1661 52.4337
R18428 vdd.n1724 vdd.n1662 52.4337
R18429 vdd.n1728 vdd.n1663 52.4337
R18430 vdd.n1730 vdd.n1664 52.4337
R18431 vdd.n1734 vdd.n1665 52.4337
R18432 vdd.n1736 vdd.n1666 52.4337
R18433 vdd.n1740 vdd.n1667 52.4337
R18434 vdd.n1741 vdd.n1668 52.4337
R18435 vdd.n1745 vdd.n1669 52.4337
R18436 vdd.n1747 vdd.n1670 52.4337
R18437 vdd.n1751 vdd.n1671 52.4337
R18438 vdd.n1753 vdd.n1672 52.4337
R18439 vdd.n1757 vdd.n1673 52.4337
R18440 vdd.n1759 vdd.n1674 52.4337
R18441 vdd.n1763 vdd.n1675 52.4337
R18442 vdd.n1765 vdd.n1676 52.4337
R18443 vdd.n1769 vdd.n1677 52.4337
R18444 vdd.n1771 vdd.n1678 52.4337
R18445 vdd.n1526 vdd.n1525 52.4337
R18446 vdd.n1523 vdd.n1522 52.4337
R18447 vdd.n1519 vdd.n1276 52.4337
R18448 vdd.n2373 vdd.n2372 52.4337
R18449 vdd.n1275 vdd.n1269 52.4337
R18450 vdd.n2380 vdd.n2379 52.4337
R18451 vdd.n1268 vdd.n1262 52.4337
R18452 vdd.n2387 vdd.n2386 52.4337
R18453 vdd.n1261 vdd.n1256 52.4337
R18454 vdd.n2394 vdd.n2393 52.4337
R18455 vdd.n1255 vdd.n1254 52.4337
R18456 vdd.n1250 vdd.n1243 52.4337
R18457 vdd.n2405 vdd.n2404 52.4337
R18458 vdd.n1242 vdd.n1236 52.4337
R18459 vdd.n2412 vdd.n2411 52.4337
R18460 vdd.n1235 vdd.n1229 52.4337
R18461 vdd.n2419 vdd.n2418 52.4337
R18462 vdd.n1228 vdd.n1222 52.4337
R18463 vdd.n2426 vdd.n2425 52.4337
R18464 vdd.n1221 vdd.n1216 52.4337
R18465 vdd.n2433 vdd.n2432 52.4337
R18466 vdd.n1215 vdd.n1214 52.4337
R18467 vdd.n1210 vdd.n1203 52.4337
R18468 vdd.n2444 vdd.n2443 52.4337
R18469 vdd.n1202 vdd.n1196 52.4337
R18470 vdd.n2451 vdd.n2450 52.4337
R18471 vdd.n1195 vdd.n1189 52.4337
R18472 vdd.n2458 vdd.n2457 52.4337
R18473 vdd.n1188 vdd.n1185 52.4337
R18474 vdd.n2465 vdd.n2464 52.4337
R18475 vdd.n2470 vdd.n2469 52.4337
R18476 vdd.n1530 vdd.n1184 52.4337
R18477 vdd.n3494 vdd.n725 52.4337
R18478 vdd.n733 vdd.n693 52.4337
R18479 vdd.n3484 vdd.n694 52.4337
R18480 vdd.n3480 vdd.n695 52.4337
R18481 vdd.n3476 vdd.n696 52.4337
R18482 vdd.n3472 vdd.n697 52.4337
R18483 vdd.n3468 vdd.n698 52.4337
R18484 vdd.n3464 vdd.n699 52.4337
R18485 vdd.n3460 vdd.n700 52.4337
R18486 vdd.n3450 vdd.n701 52.4337
R18487 vdd.n3448 vdd.n702 52.4337
R18488 vdd.n3444 vdd.n703 52.4337
R18489 vdd.n3440 vdd.n704 52.4337
R18490 vdd.n3436 vdd.n705 52.4337
R18491 vdd.n3432 vdd.n706 52.4337
R18492 vdd.n3428 vdd.n707 52.4337
R18493 vdd.n3424 vdd.n708 52.4337
R18494 vdd.n3420 vdd.n709 52.4337
R18495 vdd.n3416 vdd.n710 52.4337
R18496 vdd.n3412 vdd.n711 52.4337
R18497 vdd.n3404 vdd.n712 52.4337
R18498 vdd.n3402 vdd.n713 52.4337
R18499 vdd.n3398 vdd.n714 52.4337
R18500 vdd.n3394 vdd.n715 52.4337
R18501 vdd.n3390 vdd.n716 52.4337
R18502 vdd.n3386 vdd.n717 52.4337
R18503 vdd.n3382 vdd.n718 52.4337
R18504 vdd.n3378 vdd.n719 52.4337
R18505 vdd.n3374 vdd.n720 52.4337
R18506 vdd.n3370 vdd.n721 52.4337
R18507 vdd.n722 vdd.n691 52.4337
R18508 vdd.n3625 vdd.n425 52.4337
R18509 vdd.n614 vdd.n424 52.4337
R18510 vdd.n608 vdd.n423 52.4337
R18511 vdd.n604 vdd.n422 52.4337
R18512 vdd.n598 vdd.n421 52.4337
R18513 vdd.n594 vdd.n420 52.4337
R18514 vdd.n588 vdd.n419 52.4337
R18515 vdd.n584 vdd.n418 52.4337
R18516 vdd.n578 vdd.n417 52.4337
R18517 vdd.n574 vdd.n416 52.4337
R18518 vdd.n568 vdd.n415 52.4337
R18519 vdd.n564 vdd.n414 52.4337
R18520 vdd.n558 vdd.n413 52.4337
R18521 vdd.n554 vdd.n412 52.4337
R18522 vdd.n548 vdd.n411 52.4337
R18523 vdd.n544 vdd.n410 52.4337
R18524 vdd.n538 vdd.n409 52.4337
R18525 vdd.n534 vdd.n408 52.4337
R18526 vdd.n528 vdd.n407 52.4337
R18527 vdd.n524 vdd.n406 52.4337
R18528 vdd.n518 vdd.n405 52.4337
R18529 vdd.n514 vdd.n404 52.4337
R18530 vdd.n508 vdd.n403 52.4337
R18531 vdd.n504 vdd.n402 52.4337
R18532 vdd.n498 vdd.n401 52.4337
R18533 vdd.n494 vdd.n400 52.4337
R18534 vdd.n488 vdd.n399 52.4337
R18535 vdd.n484 vdd.n398 52.4337
R18536 vdd.n478 vdd.n397 52.4337
R18537 vdd.n474 vdd.n396 52.4337
R18538 vdd.n468 vdd.n395 52.4337
R18539 vdd.n394 vdd.n392 52.4337
R18540 vdd.t240 vdd.t264 51.4683
R18541 vdd.n274 vdd.n272 42.0461
R18542 vdd.n172 vdd.n170 42.0461
R18543 vdd.n71 vdd.n69 42.0461
R18544 vdd.n2207 vdd.n2205 42.0461
R18545 vdd.n2105 vdd.n2103 42.0461
R18546 vdd.n2004 vdd.n2002 42.0461
R18547 vdd.n332 vdd.n331 41.6884
R18548 vdd.n230 vdd.n229 41.6884
R18549 vdd.n129 vdd.n128 41.6884
R18550 vdd.n2265 vdd.n2264 41.6884
R18551 vdd.n2163 vdd.n2162 41.6884
R18552 vdd.n2062 vdd.n2061 41.6884
R18553 vdd.n1774 vdd.n1773 41.1157
R18554 vdd.n1812 vdd.n1811 41.1157
R18555 vdd.n1708 vdd.n1707 41.1157
R18556 vdd.n428 vdd.n427 41.1157
R18557 vdd.n566 vdd.n441 41.1157
R18558 vdd.n454 vdd.n453 41.1157
R18559 vdd.n3325 vdd.n3324 39.2114
R18560 vdd.n3322 vdd.n3321 39.2114
R18561 vdd.n3317 vdd.n815 39.2114
R18562 vdd.n3315 vdd.n3314 39.2114
R18563 vdd.n3310 vdd.n818 39.2114
R18564 vdd.n3308 vdd.n3307 39.2114
R18565 vdd.n3303 vdd.n821 39.2114
R18566 vdd.n3301 vdd.n3300 39.2114
R18567 vdd.n3297 vdd.n3296 39.2114
R18568 vdd.n3292 vdd.n824 39.2114
R18569 vdd.n3290 vdd.n3289 39.2114
R18570 vdd.n3285 vdd.n827 39.2114
R18571 vdd.n3283 vdd.n3282 39.2114
R18572 vdd.n3278 vdd.n830 39.2114
R18573 vdd.n3276 vdd.n3275 39.2114
R18574 vdd.n3270 vdd.n835 39.2114
R18575 vdd.n3268 vdd.n3267 39.2114
R18576 vdd.n3090 vdd.n3089 39.2114
R18577 vdd.n2819 vdd.n2785 39.2114
R18578 vdd.n3082 vdd.n2786 39.2114
R18579 vdd.n3078 vdd.n2787 39.2114
R18580 vdd.n3074 vdd.n2788 39.2114
R18581 vdd.n3070 vdd.n2789 39.2114
R18582 vdd.n3066 vdd.n2790 39.2114
R18583 vdd.n3062 vdd.n2791 39.2114
R18584 vdd.n3058 vdd.n2792 39.2114
R18585 vdd.n3054 vdd.n2793 39.2114
R18586 vdd.n3050 vdd.n2794 39.2114
R18587 vdd.n3046 vdd.n2795 39.2114
R18588 vdd.n3042 vdd.n2796 39.2114
R18589 vdd.n3038 vdd.n2797 39.2114
R18590 vdd.n3034 vdd.n2798 39.2114
R18591 vdd.n3030 vdd.n2799 39.2114
R18592 vdd.n3025 vdd.n2800 39.2114
R18593 vdd.n2779 vdd.n997 39.2114
R18594 vdd.n2775 vdd.n996 39.2114
R18595 vdd.n2771 vdd.n995 39.2114
R18596 vdd.n2767 vdd.n994 39.2114
R18597 vdd.n2763 vdd.n993 39.2114
R18598 vdd.n2759 vdd.n992 39.2114
R18599 vdd.n2755 vdd.n991 39.2114
R18600 vdd.n2751 vdd.n990 39.2114
R18601 vdd.n2747 vdd.n989 39.2114
R18602 vdd.n2743 vdd.n988 39.2114
R18603 vdd.n2739 vdd.n987 39.2114
R18604 vdd.n2735 vdd.n986 39.2114
R18605 vdd.n2731 vdd.n985 39.2114
R18606 vdd.n2727 vdd.n984 39.2114
R18607 vdd.n2723 vdd.n983 39.2114
R18608 vdd.n2718 vdd.n982 39.2114
R18609 vdd.n2714 vdd.n981 39.2114
R18610 vdd.n2508 vdd.n2507 39.2114
R18611 vdd.n1176 vdd.n1142 39.2114
R18612 vdd.n2500 vdd.n1143 39.2114
R18613 vdd.n2496 vdd.n1144 39.2114
R18614 vdd.n2492 vdd.n1145 39.2114
R18615 vdd.n2488 vdd.n1146 39.2114
R18616 vdd.n2484 vdd.n1147 39.2114
R18617 vdd.n2480 vdd.n1148 39.2114
R18618 vdd.n2476 vdd.n1149 39.2114
R18619 vdd.n1322 vdd.n1150 39.2114
R18620 vdd.n1326 vdd.n1151 39.2114
R18621 vdd.n1330 vdd.n1152 39.2114
R18622 vdd.n1334 vdd.n1153 39.2114
R18623 vdd.n1338 vdd.n1154 39.2114
R18624 vdd.n1342 vdd.n1155 39.2114
R18625 vdd.n1346 vdd.n1156 39.2114
R18626 vdd.n1351 vdd.n1157 39.2114
R18627 vdd.n3244 vdd.n3243 39.2114
R18628 vdd.n3239 vdd.n3211 39.2114
R18629 vdd.n3237 vdd.n3236 39.2114
R18630 vdd.n3232 vdd.n3214 39.2114
R18631 vdd.n3230 vdd.n3229 39.2114
R18632 vdd.n3225 vdd.n3217 39.2114
R18633 vdd.n3223 vdd.n3222 39.2114
R18634 vdd.n3218 vdd.n787 39.2114
R18635 vdd.n3362 vdd.n3361 39.2114
R18636 vdd.n3359 vdd.n3358 39.2114
R18637 vdd.n3354 vdd.n791 39.2114
R18638 vdd.n3352 vdd.n3351 39.2114
R18639 vdd.n3347 vdd.n794 39.2114
R18640 vdd.n3345 vdd.n3344 39.2114
R18641 vdd.n3340 vdd.n797 39.2114
R18642 vdd.n3338 vdd.n3337 39.2114
R18643 vdd.n3333 vdd.n803 39.2114
R18644 vdd.n2826 vdd.n2801 39.2114
R18645 vdd.n2830 vdd.n2802 39.2114
R18646 vdd.n2834 vdd.n2803 39.2114
R18647 vdd.n2838 vdd.n2804 39.2114
R18648 vdd.n2842 vdd.n2805 39.2114
R18649 vdd.n2846 vdd.n2806 39.2114
R18650 vdd.n2850 vdd.n2807 39.2114
R18651 vdd.n2854 vdd.n2808 39.2114
R18652 vdd.n2858 vdd.n2809 39.2114
R18653 vdd.n2862 vdd.n2810 39.2114
R18654 vdd.n2866 vdd.n2811 39.2114
R18655 vdd.n2870 vdd.n2812 39.2114
R18656 vdd.n2874 vdd.n2813 39.2114
R18657 vdd.n2878 vdd.n2814 39.2114
R18658 vdd.n2882 vdd.n2815 39.2114
R18659 vdd.n2886 vdd.n2816 39.2114
R18660 vdd.n2890 vdd.n2817 39.2114
R18661 vdd.n2829 vdd.n2801 39.2114
R18662 vdd.n2833 vdd.n2802 39.2114
R18663 vdd.n2837 vdd.n2803 39.2114
R18664 vdd.n2841 vdd.n2804 39.2114
R18665 vdd.n2845 vdd.n2805 39.2114
R18666 vdd.n2849 vdd.n2806 39.2114
R18667 vdd.n2853 vdd.n2807 39.2114
R18668 vdd.n2857 vdd.n2808 39.2114
R18669 vdd.n2861 vdd.n2809 39.2114
R18670 vdd.n2865 vdd.n2810 39.2114
R18671 vdd.n2869 vdd.n2811 39.2114
R18672 vdd.n2873 vdd.n2812 39.2114
R18673 vdd.n2877 vdd.n2813 39.2114
R18674 vdd.n2881 vdd.n2814 39.2114
R18675 vdd.n2885 vdd.n2815 39.2114
R18676 vdd.n2889 vdd.n2816 39.2114
R18677 vdd.n2892 vdd.n2817 39.2114
R18678 vdd.n803 vdd.n798 39.2114
R18679 vdd.n3339 vdd.n3338 39.2114
R18680 vdd.n797 vdd.n795 39.2114
R18681 vdd.n3346 vdd.n3345 39.2114
R18682 vdd.n794 vdd.n792 39.2114
R18683 vdd.n3353 vdd.n3352 39.2114
R18684 vdd.n791 vdd.n789 39.2114
R18685 vdd.n3360 vdd.n3359 39.2114
R18686 vdd.n3363 vdd.n3362 39.2114
R18687 vdd.n3219 vdd.n3218 39.2114
R18688 vdd.n3224 vdd.n3223 39.2114
R18689 vdd.n3217 vdd.n3215 39.2114
R18690 vdd.n3231 vdd.n3230 39.2114
R18691 vdd.n3214 vdd.n3212 39.2114
R18692 vdd.n3238 vdd.n3237 39.2114
R18693 vdd.n3211 vdd.n3209 39.2114
R18694 vdd.n3245 vdd.n3244 39.2114
R18695 vdd.n2507 vdd.n1140 39.2114
R18696 vdd.n2501 vdd.n1142 39.2114
R18697 vdd.n2497 vdd.n1143 39.2114
R18698 vdd.n2493 vdd.n1144 39.2114
R18699 vdd.n2489 vdd.n1145 39.2114
R18700 vdd.n2485 vdd.n1146 39.2114
R18701 vdd.n2481 vdd.n1147 39.2114
R18702 vdd.n2477 vdd.n1148 39.2114
R18703 vdd.n1321 vdd.n1149 39.2114
R18704 vdd.n1325 vdd.n1150 39.2114
R18705 vdd.n1329 vdd.n1151 39.2114
R18706 vdd.n1333 vdd.n1152 39.2114
R18707 vdd.n1337 vdd.n1153 39.2114
R18708 vdd.n1341 vdd.n1154 39.2114
R18709 vdd.n1345 vdd.n1155 39.2114
R18710 vdd.n1350 vdd.n1156 39.2114
R18711 vdd.n1354 vdd.n1157 39.2114
R18712 vdd.n2717 vdd.n981 39.2114
R18713 vdd.n2722 vdd.n982 39.2114
R18714 vdd.n2726 vdd.n983 39.2114
R18715 vdd.n2730 vdd.n984 39.2114
R18716 vdd.n2734 vdd.n985 39.2114
R18717 vdd.n2738 vdd.n986 39.2114
R18718 vdd.n2742 vdd.n987 39.2114
R18719 vdd.n2746 vdd.n988 39.2114
R18720 vdd.n2750 vdd.n989 39.2114
R18721 vdd.n2754 vdd.n990 39.2114
R18722 vdd.n2758 vdd.n991 39.2114
R18723 vdd.n2762 vdd.n992 39.2114
R18724 vdd.n2766 vdd.n993 39.2114
R18725 vdd.n2770 vdd.n994 39.2114
R18726 vdd.n2774 vdd.n995 39.2114
R18727 vdd.n2778 vdd.n996 39.2114
R18728 vdd.n999 vdd.n997 39.2114
R18729 vdd.n3089 vdd.n962 39.2114
R18730 vdd.n3083 vdd.n2785 39.2114
R18731 vdd.n3079 vdd.n2786 39.2114
R18732 vdd.n3075 vdd.n2787 39.2114
R18733 vdd.n3071 vdd.n2788 39.2114
R18734 vdd.n3067 vdd.n2789 39.2114
R18735 vdd.n3063 vdd.n2790 39.2114
R18736 vdd.n3059 vdd.n2791 39.2114
R18737 vdd.n3055 vdd.n2792 39.2114
R18738 vdd.n3051 vdd.n2793 39.2114
R18739 vdd.n3047 vdd.n2794 39.2114
R18740 vdd.n3043 vdd.n2795 39.2114
R18741 vdd.n3039 vdd.n2796 39.2114
R18742 vdd.n3035 vdd.n2797 39.2114
R18743 vdd.n3031 vdd.n2798 39.2114
R18744 vdd.n3026 vdd.n2799 39.2114
R18745 vdd.n3022 vdd.n2800 39.2114
R18746 vdd.n3269 vdd.n3268 39.2114
R18747 vdd.n835 vdd.n831 39.2114
R18748 vdd.n3277 vdd.n3276 39.2114
R18749 vdd.n830 vdd.n828 39.2114
R18750 vdd.n3284 vdd.n3283 39.2114
R18751 vdd.n827 vdd.n825 39.2114
R18752 vdd.n3291 vdd.n3290 39.2114
R18753 vdd.n824 vdd.n822 39.2114
R18754 vdd.n3298 vdd.n3297 39.2114
R18755 vdd.n3302 vdd.n3301 39.2114
R18756 vdd.n821 vdd.n819 39.2114
R18757 vdd.n3309 vdd.n3308 39.2114
R18758 vdd.n818 vdd.n816 39.2114
R18759 vdd.n3316 vdd.n3315 39.2114
R18760 vdd.n815 vdd.n813 39.2114
R18761 vdd.n3323 vdd.n3322 39.2114
R18762 vdd.n3326 vdd.n3325 39.2114
R18763 vdd.n1008 vdd.n963 39.2114
R18764 vdd.n2706 vdd.n964 39.2114
R18765 vdd.n2702 vdd.n965 39.2114
R18766 vdd.n2698 vdd.n966 39.2114
R18767 vdd.n2694 vdd.n967 39.2114
R18768 vdd.n2690 vdd.n968 39.2114
R18769 vdd.n2686 vdd.n969 39.2114
R18770 vdd.n2682 vdd.n970 39.2114
R18771 vdd.n2678 vdd.n971 39.2114
R18772 vdd.n2674 vdd.n972 39.2114
R18773 vdd.n2670 vdd.n973 39.2114
R18774 vdd.n2666 vdd.n974 39.2114
R18775 vdd.n2662 vdd.n975 39.2114
R18776 vdd.n2658 vdd.n976 39.2114
R18777 vdd.n2654 vdd.n977 39.2114
R18778 vdd.n2650 vdd.n978 39.2114
R18779 vdd.n2646 vdd.n979 39.2114
R18780 vdd.n1280 vdd.n1158 39.2114
R18781 vdd.n1284 vdd.n1159 39.2114
R18782 vdd.n1288 vdd.n1160 39.2114
R18783 vdd.n1292 vdd.n1161 39.2114
R18784 vdd.n1296 vdd.n1162 39.2114
R18785 vdd.n1300 vdd.n1163 39.2114
R18786 vdd.n1304 vdd.n1164 39.2114
R18787 vdd.n1308 vdd.n1165 39.2114
R18788 vdd.n1312 vdd.n1166 39.2114
R18789 vdd.n1513 vdd.n1167 39.2114
R18790 vdd.n1510 vdd.n1168 39.2114
R18791 vdd.n1506 vdd.n1169 39.2114
R18792 vdd.n1502 vdd.n1170 39.2114
R18793 vdd.n1498 vdd.n1171 39.2114
R18794 vdd.n1494 vdd.n1172 39.2114
R18795 vdd.n1490 vdd.n1173 39.2114
R18796 vdd.n1486 vdd.n1174 39.2114
R18797 vdd.n2643 vdd.n979 39.2114
R18798 vdd.n2647 vdd.n978 39.2114
R18799 vdd.n2651 vdd.n977 39.2114
R18800 vdd.n2655 vdd.n976 39.2114
R18801 vdd.n2659 vdd.n975 39.2114
R18802 vdd.n2663 vdd.n974 39.2114
R18803 vdd.n2667 vdd.n973 39.2114
R18804 vdd.n2671 vdd.n972 39.2114
R18805 vdd.n2675 vdd.n971 39.2114
R18806 vdd.n2679 vdd.n970 39.2114
R18807 vdd.n2683 vdd.n969 39.2114
R18808 vdd.n2687 vdd.n968 39.2114
R18809 vdd.n2691 vdd.n967 39.2114
R18810 vdd.n2695 vdd.n966 39.2114
R18811 vdd.n2699 vdd.n965 39.2114
R18812 vdd.n2703 vdd.n964 39.2114
R18813 vdd.n2707 vdd.n963 39.2114
R18814 vdd.n1283 vdd.n1158 39.2114
R18815 vdd.n1287 vdd.n1159 39.2114
R18816 vdd.n1291 vdd.n1160 39.2114
R18817 vdd.n1295 vdd.n1161 39.2114
R18818 vdd.n1299 vdd.n1162 39.2114
R18819 vdd.n1303 vdd.n1163 39.2114
R18820 vdd.n1307 vdd.n1164 39.2114
R18821 vdd.n1311 vdd.n1165 39.2114
R18822 vdd.n1314 vdd.n1166 39.2114
R18823 vdd.n1511 vdd.n1167 39.2114
R18824 vdd.n1507 vdd.n1168 39.2114
R18825 vdd.n1503 vdd.n1169 39.2114
R18826 vdd.n1499 vdd.n1170 39.2114
R18827 vdd.n1495 vdd.n1171 39.2114
R18828 vdd.n1491 vdd.n1172 39.2114
R18829 vdd.n1487 vdd.n1173 39.2114
R18830 vdd.n1483 vdd.n1174 39.2114
R18831 vdd.n2364 vdd.n2363 37.2369
R18832 vdd.n2400 vdd.n1249 37.2369
R18833 vdd.n2439 vdd.n1209 37.2369
R18834 vdd.n3410 vdd.n769 37.2369
R18835 vdd.n3458 vdd.n3457 37.2369
R18836 vdd.n690 vdd.n689 37.2369
R18837 vdd.n1317 vdd.n1316 30.449
R18838 vdd.n1012 vdd.n1011 30.449
R18839 vdd.n1348 vdd.n1320 30.449
R18840 vdd.n2720 vdd.n1002 30.449
R18841 vdd.n2825 vdd.n2824 30.449
R18842 vdd.n3272 vdd.n833 30.449
R18843 vdd.n3028 vdd.n2821 30.449
R18844 vdd.n801 vdd.n800 30.449
R18845 vdd.n2510 vdd.n2509 29.8151
R18846 vdd.n2782 vdd.n1000 29.8151
R18847 vdd.n2715 vdd.n1003 29.8151
R18848 vdd.n1356 vdd.n1353 29.8151
R18849 vdd.n3023 vdd.n3020 29.8151
R18850 vdd.n3266 vdd.n3265 29.8151
R18851 vdd.n3092 vdd.n3091 29.8151
R18852 vdd.n3329 vdd.n3328 29.8151
R18853 vdd.n3248 vdd.n3247 29.8151
R18854 vdd.n3334 vdd.n802 29.8151
R18855 vdd.n2896 vdd.n2894 29.8151
R18856 vdd.n2827 vdd.n955 29.8151
R18857 vdd.n1281 vdd.n1132 29.8151
R18858 vdd.n2710 vdd.n2709 29.8151
R18859 vdd.n2642 vdd.n2641 29.8151
R18860 vdd.n1482 vdd.n1481 29.8151
R18861 vdd.n1873 vdd.n1680 22.2201
R18862 vdd.n2358 vdd.n1141 22.2201
R18863 vdd.n3495 vdd.n723 22.2201
R18864 vdd.n3627 vdd.n3626 22.2201
R18865 vdd.n1884 vdd.n1642 19.3944
R18866 vdd.n1884 vdd.n1640 19.3944
R18867 vdd.n1888 vdd.n1640 19.3944
R18868 vdd.n1888 vdd.n1630 19.3944
R18869 vdd.n1901 vdd.n1630 19.3944
R18870 vdd.n1901 vdd.n1628 19.3944
R18871 vdd.n1905 vdd.n1628 19.3944
R18872 vdd.n1905 vdd.n1620 19.3944
R18873 vdd.n1918 vdd.n1620 19.3944
R18874 vdd.n1918 vdd.n1618 19.3944
R18875 vdd.n1922 vdd.n1618 19.3944
R18876 vdd.n1922 vdd.n1607 19.3944
R18877 vdd.n1934 vdd.n1607 19.3944
R18878 vdd.n1934 vdd.n1605 19.3944
R18879 vdd.n1938 vdd.n1605 19.3944
R18880 vdd.n1938 vdd.n1596 19.3944
R18881 vdd.n1951 vdd.n1596 19.3944
R18882 vdd.n1951 vdd.n1594 19.3944
R18883 vdd.n1955 vdd.n1594 19.3944
R18884 vdd.n1955 vdd.n1585 19.3944
R18885 vdd.n2274 vdd.n1585 19.3944
R18886 vdd.n2274 vdd.n1583 19.3944
R18887 vdd.n2278 vdd.n1583 19.3944
R18888 vdd.n2278 vdd.n1573 19.3944
R18889 vdd.n2291 vdd.n1573 19.3944
R18890 vdd.n2291 vdd.n1571 19.3944
R18891 vdd.n2295 vdd.n1571 19.3944
R18892 vdd.n2295 vdd.n1563 19.3944
R18893 vdd.n2308 vdd.n1563 19.3944
R18894 vdd.n2308 vdd.n1561 19.3944
R18895 vdd.n2312 vdd.n1561 19.3944
R18896 vdd.n2312 vdd.n1550 19.3944
R18897 vdd.n2324 vdd.n1550 19.3944
R18898 vdd.n2324 vdd.n1548 19.3944
R18899 vdd.n2328 vdd.n1548 19.3944
R18900 vdd.n2328 vdd.n1540 19.3944
R18901 vdd.n2341 vdd.n1540 19.3944
R18902 vdd.n2341 vdd.n1537 19.3944
R18903 vdd.n2347 vdd.n1537 19.3944
R18904 vdd.n2347 vdd.n1538 19.3944
R18905 vdd.n1538 vdd.n1528 19.3944
R18906 vdd.n1808 vdd.n1743 19.3944
R18907 vdd.n1804 vdd.n1743 19.3944
R18908 vdd.n1804 vdd.n1803 19.3944
R18909 vdd.n1803 vdd.n1802 19.3944
R18910 vdd.n1802 vdd.n1749 19.3944
R18911 vdd.n1798 vdd.n1749 19.3944
R18912 vdd.n1798 vdd.n1797 19.3944
R18913 vdd.n1797 vdd.n1796 19.3944
R18914 vdd.n1796 vdd.n1755 19.3944
R18915 vdd.n1792 vdd.n1755 19.3944
R18916 vdd.n1792 vdd.n1791 19.3944
R18917 vdd.n1791 vdd.n1790 19.3944
R18918 vdd.n1790 vdd.n1761 19.3944
R18919 vdd.n1786 vdd.n1761 19.3944
R18920 vdd.n1786 vdd.n1785 19.3944
R18921 vdd.n1785 vdd.n1784 19.3944
R18922 vdd.n1784 vdd.n1767 19.3944
R18923 vdd.n1780 vdd.n1767 19.3944
R18924 vdd.n1780 vdd.n1779 19.3944
R18925 vdd.n1779 vdd.n1778 19.3944
R18926 vdd.n1843 vdd.n1842 19.3944
R18927 vdd.n1842 vdd.n1841 19.3944
R18928 vdd.n1841 vdd.n1714 19.3944
R18929 vdd.n1837 vdd.n1714 19.3944
R18930 vdd.n1837 vdd.n1836 19.3944
R18931 vdd.n1836 vdd.n1835 19.3944
R18932 vdd.n1835 vdd.n1720 19.3944
R18933 vdd.n1831 vdd.n1720 19.3944
R18934 vdd.n1831 vdd.n1830 19.3944
R18935 vdd.n1830 vdd.n1829 19.3944
R18936 vdd.n1829 vdd.n1726 19.3944
R18937 vdd.n1825 vdd.n1726 19.3944
R18938 vdd.n1825 vdd.n1824 19.3944
R18939 vdd.n1824 vdd.n1823 19.3944
R18940 vdd.n1823 vdd.n1732 19.3944
R18941 vdd.n1819 vdd.n1732 19.3944
R18942 vdd.n1819 vdd.n1818 19.3944
R18943 vdd.n1818 vdd.n1817 19.3944
R18944 vdd.n1817 vdd.n1738 19.3944
R18945 vdd.n1813 vdd.n1738 19.3944
R18946 vdd.n1876 vdd.n1647 19.3944
R18947 vdd.n1871 vdd.n1647 19.3944
R18948 vdd.n1871 vdd.n1682 19.3944
R18949 vdd.n1867 vdd.n1682 19.3944
R18950 vdd.n1867 vdd.n1866 19.3944
R18951 vdd.n1866 vdd.n1865 19.3944
R18952 vdd.n1865 vdd.n1688 19.3944
R18953 vdd.n1861 vdd.n1688 19.3944
R18954 vdd.n1861 vdd.n1860 19.3944
R18955 vdd.n1860 vdd.n1859 19.3944
R18956 vdd.n1859 vdd.n1694 19.3944
R18957 vdd.n1855 vdd.n1694 19.3944
R18958 vdd.n1855 vdd.n1854 19.3944
R18959 vdd.n1854 vdd.n1853 19.3944
R18960 vdd.n1853 vdd.n1700 19.3944
R18961 vdd.n1849 vdd.n1700 19.3944
R18962 vdd.n1849 vdd.n1848 19.3944
R18963 vdd.n1848 vdd.n1847 19.3944
R18964 vdd.n2396 vdd.n1247 19.3944
R18965 vdd.n2396 vdd.n1253 19.3944
R18966 vdd.n2391 vdd.n1253 19.3944
R18967 vdd.n2391 vdd.n2390 19.3944
R18968 vdd.n2390 vdd.n2389 19.3944
R18969 vdd.n2389 vdd.n1260 19.3944
R18970 vdd.n2384 vdd.n1260 19.3944
R18971 vdd.n2384 vdd.n2383 19.3944
R18972 vdd.n2383 vdd.n2382 19.3944
R18973 vdd.n2382 vdd.n1267 19.3944
R18974 vdd.n2377 vdd.n1267 19.3944
R18975 vdd.n2377 vdd.n2376 19.3944
R18976 vdd.n2376 vdd.n2375 19.3944
R18977 vdd.n2375 vdd.n1274 19.3944
R18978 vdd.n2370 vdd.n1274 19.3944
R18979 vdd.n2370 vdd.n2369 19.3944
R18980 vdd.n1521 vdd.n1279 19.3944
R18981 vdd.n2365 vdd.n1518 19.3944
R18982 vdd.n2435 vdd.n1207 19.3944
R18983 vdd.n2435 vdd.n1213 19.3944
R18984 vdd.n2430 vdd.n1213 19.3944
R18985 vdd.n2430 vdd.n2429 19.3944
R18986 vdd.n2429 vdd.n2428 19.3944
R18987 vdd.n2428 vdd.n1220 19.3944
R18988 vdd.n2423 vdd.n1220 19.3944
R18989 vdd.n2423 vdd.n2422 19.3944
R18990 vdd.n2422 vdd.n2421 19.3944
R18991 vdd.n2421 vdd.n1227 19.3944
R18992 vdd.n2416 vdd.n1227 19.3944
R18993 vdd.n2416 vdd.n2415 19.3944
R18994 vdd.n2415 vdd.n2414 19.3944
R18995 vdd.n2414 vdd.n1234 19.3944
R18996 vdd.n2409 vdd.n1234 19.3944
R18997 vdd.n2409 vdd.n2408 19.3944
R18998 vdd.n2408 vdd.n2407 19.3944
R18999 vdd.n2407 vdd.n1241 19.3944
R19000 vdd.n2402 vdd.n1241 19.3944
R19001 vdd.n2402 vdd.n2401 19.3944
R19002 vdd.n2472 vdd.n1182 19.3944
R19003 vdd.n2472 vdd.n1183 19.3944
R19004 vdd.n2467 vdd.n2466 19.3944
R19005 vdd.n2462 vdd.n2461 19.3944
R19006 vdd.n2461 vdd.n2460 19.3944
R19007 vdd.n2460 vdd.n1187 19.3944
R19008 vdd.n2455 vdd.n1187 19.3944
R19009 vdd.n2455 vdd.n2454 19.3944
R19010 vdd.n2454 vdd.n2453 19.3944
R19011 vdd.n2453 vdd.n1194 19.3944
R19012 vdd.n2448 vdd.n1194 19.3944
R19013 vdd.n2448 vdd.n2447 19.3944
R19014 vdd.n2447 vdd.n2446 19.3944
R19015 vdd.n2446 vdd.n1201 19.3944
R19016 vdd.n2441 vdd.n1201 19.3944
R19017 vdd.n2441 vdd.n2440 19.3944
R19018 vdd.n1880 vdd.n1645 19.3944
R19019 vdd.n1880 vdd.n1636 19.3944
R19020 vdd.n1893 vdd.n1636 19.3944
R19021 vdd.n1893 vdd.n1634 19.3944
R19022 vdd.n1897 vdd.n1634 19.3944
R19023 vdd.n1897 vdd.n1625 19.3944
R19024 vdd.n1910 vdd.n1625 19.3944
R19025 vdd.n1910 vdd.n1623 19.3944
R19026 vdd.n1914 vdd.n1623 19.3944
R19027 vdd.n1914 vdd.n1614 19.3944
R19028 vdd.n1926 vdd.n1614 19.3944
R19029 vdd.n1926 vdd.n1612 19.3944
R19030 vdd.n1930 vdd.n1612 19.3944
R19031 vdd.n1930 vdd.n1602 19.3944
R19032 vdd.n1943 vdd.n1602 19.3944
R19033 vdd.n1943 vdd.n1600 19.3944
R19034 vdd.n1947 vdd.n1600 19.3944
R19035 vdd.n1947 vdd.n1591 19.3944
R19036 vdd.n1959 vdd.n1591 19.3944
R19037 vdd.n1959 vdd.n1589 19.3944
R19038 vdd.n2270 vdd.n1589 19.3944
R19039 vdd.n2270 vdd.n1579 19.3944
R19040 vdd.n2283 vdd.n1579 19.3944
R19041 vdd.n2283 vdd.n1577 19.3944
R19042 vdd.n2287 vdd.n1577 19.3944
R19043 vdd.n2287 vdd.n1568 19.3944
R19044 vdd.n2300 vdd.n1568 19.3944
R19045 vdd.n2300 vdd.n1566 19.3944
R19046 vdd.n2304 vdd.n1566 19.3944
R19047 vdd.n2304 vdd.n1557 19.3944
R19048 vdd.n2316 vdd.n1557 19.3944
R19049 vdd.n2316 vdd.n1555 19.3944
R19050 vdd.n2320 vdd.n1555 19.3944
R19051 vdd.n2320 vdd.n1545 19.3944
R19052 vdd.n2333 vdd.n1545 19.3944
R19053 vdd.n2333 vdd.n1543 19.3944
R19054 vdd.n2337 vdd.n1543 19.3944
R19055 vdd.n2337 vdd.n1533 19.3944
R19056 vdd.n2352 vdd.n1533 19.3944
R19057 vdd.n2352 vdd.n1531 19.3944
R19058 vdd.n2356 vdd.n1531 19.3944
R19059 vdd.n3501 vdd.n686 19.3944
R19060 vdd.n3501 vdd.n676 19.3944
R19061 vdd.n3513 vdd.n676 19.3944
R19062 vdd.n3513 vdd.n674 19.3944
R19063 vdd.n3517 vdd.n674 19.3944
R19064 vdd.n3517 vdd.n666 19.3944
R19065 vdd.n3530 vdd.n666 19.3944
R19066 vdd.n3530 vdd.n664 19.3944
R19067 vdd.n3534 vdd.n664 19.3944
R19068 vdd.n3534 vdd.n653 19.3944
R19069 vdd.n3546 vdd.n653 19.3944
R19070 vdd.n3546 vdd.n651 19.3944
R19071 vdd.n3550 vdd.n651 19.3944
R19072 vdd.n3550 vdd.n642 19.3944
R19073 vdd.n3563 vdd.n642 19.3944
R19074 vdd.n3563 vdd.n640 19.3944
R19075 vdd.n3570 vdd.n640 19.3944
R19076 vdd.n3570 vdd.n3569 19.3944
R19077 vdd.n3569 vdd.n631 19.3944
R19078 vdd.n3583 vdd.n631 19.3944
R19079 vdd.n3584 vdd.n3583 19.3944
R19080 vdd.n3584 vdd.n629 19.3944
R19081 vdd.n3588 vdd.n629 19.3944
R19082 vdd.n3590 vdd.n3588 19.3944
R19083 vdd.n3591 vdd.n3590 19.3944
R19084 vdd.n3591 vdd.n627 19.3944
R19085 vdd.n3595 vdd.n627 19.3944
R19086 vdd.n3597 vdd.n3595 19.3944
R19087 vdd.n3598 vdd.n3597 19.3944
R19088 vdd.n3598 vdd.n625 19.3944
R19089 vdd.n3602 vdd.n625 19.3944
R19090 vdd.n3605 vdd.n3602 19.3944
R19091 vdd.n3606 vdd.n3605 19.3944
R19092 vdd.n3606 vdd.n623 19.3944
R19093 vdd.n3610 vdd.n623 19.3944
R19094 vdd.n3612 vdd.n3610 19.3944
R19095 vdd.n3613 vdd.n3612 19.3944
R19096 vdd.n3613 vdd.n621 19.3944
R19097 vdd.n3617 vdd.n621 19.3944
R19098 vdd.n3619 vdd.n3617 19.3944
R19099 vdd.n3620 vdd.n3619 19.3944
R19100 vdd.n569 vdd.n438 19.3944
R19101 vdd.n575 vdd.n438 19.3944
R19102 vdd.n576 vdd.n575 19.3944
R19103 vdd.n579 vdd.n576 19.3944
R19104 vdd.n579 vdd.n436 19.3944
R19105 vdd.n585 vdd.n436 19.3944
R19106 vdd.n586 vdd.n585 19.3944
R19107 vdd.n589 vdd.n586 19.3944
R19108 vdd.n589 vdd.n434 19.3944
R19109 vdd.n595 vdd.n434 19.3944
R19110 vdd.n596 vdd.n595 19.3944
R19111 vdd.n599 vdd.n596 19.3944
R19112 vdd.n599 vdd.n432 19.3944
R19113 vdd.n605 vdd.n432 19.3944
R19114 vdd.n606 vdd.n605 19.3944
R19115 vdd.n609 vdd.n606 19.3944
R19116 vdd.n609 vdd.n430 19.3944
R19117 vdd.n615 vdd.n430 19.3944
R19118 vdd.n617 vdd.n615 19.3944
R19119 vdd.n618 vdd.n617 19.3944
R19120 vdd.n516 vdd.n515 19.3944
R19121 vdd.n519 vdd.n516 19.3944
R19122 vdd.n519 vdd.n450 19.3944
R19123 vdd.n525 vdd.n450 19.3944
R19124 vdd.n526 vdd.n525 19.3944
R19125 vdd.n529 vdd.n526 19.3944
R19126 vdd.n529 vdd.n448 19.3944
R19127 vdd.n535 vdd.n448 19.3944
R19128 vdd.n536 vdd.n535 19.3944
R19129 vdd.n539 vdd.n536 19.3944
R19130 vdd.n539 vdd.n446 19.3944
R19131 vdd.n545 vdd.n446 19.3944
R19132 vdd.n546 vdd.n545 19.3944
R19133 vdd.n549 vdd.n546 19.3944
R19134 vdd.n549 vdd.n444 19.3944
R19135 vdd.n555 vdd.n444 19.3944
R19136 vdd.n556 vdd.n555 19.3944
R19137 vdd.n559 vdd.n556 19.3944
R19138 vdd.n559 vdd.n442 19.3944
R19139 vdd.n565 vdd.n442 19.3944
R19140 vdd.n466 vdd.n465 19.3944
R19141 vdd.n469 vdd.n466 19.3944
R19142 vdd.n469 vdd.n462 19.3944
R19143 vdd.n475 vdd.n462 19.3944
R19144 vdd.n476 vdd.n475 19.3944
R19145 vdd.n479 vdd.n476 19.3944
R19146 vdd.n479 vdd.n460 19.3944
R19147 vdd.n485 vdd.n460 19.3944
R19148 vdd.n486 vdd.n485 19.3944
R19149 vdd.n489 vdd.n486 19.3944
R19150 vdd.n489 vdd.n458 19.3944
R19151 vdd.n495 vdd.n458 19.3944
R19152 vdd.n496 vdd.n495 19.3944
R19153 vdd.n499 vdd.n496 19.3944
R19154 vdd.n499 vdd.n456 19.3944
R19155 vdd.n505 vdd.n456 19.3944
R19156 vdd.n506 vdd.n505 19.3944
R19157 vdd.n509 vdd.n506 19.3944
R19158 vdd.n3505 vdd.n683 19.3944
R19159 vdd.n3505 vdd.n681 19.3944
R19160 vdd.n3509 vdd.n681 19.3944
R19161 vdd.n3509 vdd.n671 19.3944
R19162 vdd.n3522 vdd.n671 19.3944
R19163 vdd.n3522 vdd.n669 19.3944
R19164 vdd.n3526 vdd.n669 19.3944
R19165 vdd.n3526 vdd.n660 19.3944
R19166 vdd.n3538 vdd.n660 19.3944
R19167 vdd.n3538 vdd.n658 19.3944
R19168 vdd.n3542 vdd.n658 19.3944
R19169 vdd.n3542 vdd.n648 19.3944
R19170 vdd.n3555 vdd.n648 19.3944
R19171 vdd.n3555 vdd.n646 19.3944
R19172 vdd.n3559 vdd.n646 19.3944
R19173 vdd.n3559 vdd.n637 19.3944
R19174 vdd.n3574 vdd.n637 19.3944
R19175 vdd.n3574 vdd.n635 19.3944
R19176 vdd.n3578 vdd.n635 19.3944
R19177 vdd.n3578 vdd.n336 19.3944
R19178 vdd.n3669 vdd.n336 19.3944
R19179 vdd.n3669 vdd.n337 19.3944
R19180 vdd.n3663 vdd.n337 19.3944
R19181 vdd.n3663 vdd.n3662 19.3944
R19182 vdd.n3662 vdd.n3661 19.3944
R19183 vdd.n3661 vdd.n349 19.3944
R19184 vdd.n3655 vdd.n349 19.3944
R19185 vdd.n3655 vdd.n3654 19.3944
R19186 vdd.n3654 vdd.n3653 19.3944
R19187 vdd.n3653 vdd.n359 19.3944
R19188 vdd.n3647 vdd.n359 19.3944
R19189 vdd.n3647 vdd.n3646 19.3944
R19190 vdd.n3646 vdd.n3645 19.3944
R19191 vdd.n3645 vdd.n370 19.3944
R19192 vdd.n3639 vdd.n370 19.3944
R19193 vdd.n3639 vdd.n3638 19.3944
R19194 vdd.n3638 vdd.n3637 19.3944
R19195 vdd.n3637 vdd.n381 19.3944
R19196 vdd.n3631 vdd.n381 19.3944
R19197 vdd.n3631 vdd.n3630 19.3944
R19198 vdd.n3630 vdd.n3629 19.3944
R19199 vdd.n3452 vdd.n747 19.3944
R19200 vdd.n3452 vdd.n3449 19.3944
R19201 vdd.n3449 vdd.n3446 19.3944
R19202 vdd.n3446 vdd.n3445 19.3944
R19203 vdd.n3445 vdd.n3442 19.3944
R19204 vdd.n3442 vdd.n3441 19.3944
R19205 vdd.n3441 vdd.n3438 19.3944
R19206 vdd.n3438 vdd.n3437 19.3944
R19207 vdd.n3437 vdd.n3434 19.3944
R19208 vdd.n3434 vdd.n3433 19.3944
R19209 vdd.n3433 vdd.n3430 19.3944
R19210 vdd.n3430 vdd.n3429 19.3944
R19211 vdd.n3429 vdd.n3426 19.3944
R19212 vdd.n3426 vdd.n3425 19.3944
R19213 vdd.n3425 vdd.n3422 19.3944
R19214 vdd.n3422 vdd.n3421 19.3944
R19215 vdd.n3421 vdd.n3418 19.3944
R19216 vdd.n3418 vdd.n3417 19.3944
R19217 vdd.n3417 vdd.n3414 19.3944
R19218 vdd.n3414 vdd.n3413 19.3944
R19219 vdd.n3492 vdd.n3491 19.3944
R19220 vdd.n3491 vdd.n3490 19.3944
R19221 vdd.n732 vdd.n729 19.3944
R19222 vdd.n3486 vdd.n3485 19.3944
R19223 vdd.n3485 vdd.n3482 19.3944
R19224 vdd.n3482 vdd.n3481 19.3944
R19225 vdd.n3481 vdd.n3478 19.3944
R19226 vdd.n3478 vdd.n3477 19.3944
R19227 vdd.n3477 vdd.n3474 19.3944
R19228 vdd.n3474 vdd.n3473 19.3944
R19229 vdd.n3473 vdd.n3470 19.3944
R19230 vdd.n3470 vdd.n3469 19.3944
R19231 vdd.n3469 vdd.n3466 19.3944
R19232 vdd.n3466 vdd.n3465 19.3944
R19233 vdd.n3465 vdd.n3462 19.3944
R19234 vdd.n3462 vdd.n3461 19.3944
R19235 vdd.n3406 vdd.n767 19.3944
R19236 vdd.n3406 vdd.n3403 19.3944
R19237 vdd.n3403 vdd.n3400 19.3944
R19238 vdd.n3400 vdd.n3399 19.3944
R19239 vdd.n3399 vdd.n3396 19.3944
R19240 vdd.n3396 vdd.n3395 19.3944
R19241 vdd.n3395 vdd.n3392 19.3944
R19242 vdd.n3392 vdd.n3391 19.3944
R19243 vdd.n3391 vdd.n3388 19.3944
R19244 vdd.n3388 vdd.n3387 19.3944
R19245 vdd.n3387 vdd.n3384 19.3944
R19246 vdd.n3384 vdd.n3383 19.3944
R19247 vdd.n3383 vdd.n3380 19.3944
R19248 vdd.n3380 vdd.n3379 19.3944
R19249 vdd.n3379 vdd.n3376 19.3944
R19250 vdd.n3376 vdd.n3375 19.3944
R19251 vdd.n3372 vdd.n3371 19.3944
R19252 vdd.n3368 vdd.n3367 19.3944
R19253 vdd.n1812 vdd.n1808 19.0066
R19254 vdd.n2400 vdd.n1247 19.0066
R19255 vdd.n569 vdd.n566 19.0066
R19256 vdd.n3410 vdd.n767 19.0066
R19257 vdd.n1316 vdd.n1315 16.0975
R19258 vdd.n1011 vdd.n1010 16.0975
R19259 vdd.n1773 vdd.n1772 16.0975
R19260 vdd.n1811 vdd.n1810 16.0975
R19261 vdd.n1707 vdd.n1706 16.0975
R19262 vdd.n2363 vdd.n2362 16.0975
R19263 vdd.n1249 vdd.n1248 16.0975
R19264 vdd.n1209 vdd.n1208 16.0975
R19265 vdd.n1320 vdd.n1319 16.0975
R19266 vdd.n1002 vdd.n1001 16.0975
R19267 vdd.n2824 vdd.n2823 16.0975
R19268 vdd.n427 vdd.n426 16.0975
R19269 vdd.n441 vdd.n440 16.0975
R19270 vdd.n453 vdd.n452 16.0975
R19271 vdd.n769 vdd.n768 16.0975
R19272 vdd.n3457 vdd.n3456 16.0975
R19273 vdd.n833 vdd.n832 16.0975
R19274 vdd.n2821 vdd.n2820 16.0975
R19275 vdd.n689 vdd.n688 16.0975
R19276 vdd.n800 vdd.n799 16.0975
R19277 vdd.t264 vdd.n2784 15.4182
R19278 vdd.n3088 vdd.t240 15.4182
R19279 vdd.n28 vdd.n27 14.7303
R19280 vdd.n328 vdd.n293 13.1884
R19281 vdd.n269 vdd.n234 13.1884
R19282 vdd.n226 vdd.n191 13.1884
R19283 vdd.n167 vdd.n132 13.1884
R19284 vdd.n125 vdd.n90 13.1884
R19285 vdd.n66 vdd.n31 13.1884
R19286 vdd.n2202 vdd.n2167 13.1884
R19287 vdd.n2261 vdd.n2226 13.1884
R19288 vdd.n2100 vdd.n2065 13.1884
R19289 vdd.n2159 vdd.n2124 13.1884
R19290 vdd.n1999 vdd.n1964 13.1884
R19291 vdd.n2058 vdd.n2023 13.1884
R19292 vdd.n2506 vdd.n1134 13.1509
R19293 vdd.n3331 vdd.n692 13.1509
R19294 vdd.n1843 vdd.n1708 12.9944
R19295 vdd.n1847 vdd.n1708 12.9944
R19296 vdd.n2439 vdd.n1207 12.9944
R19297 vdd.n2440 vdd.n2439 12.9944
R19298 vdd.n515 vdd.n454 12.9944
R19299 vdd.n509 vdd.n454 12.9944
R19300 vdd.n3458 vdd.n747 12.9944
R19301 vdd.n3461 vdd.n3458 12.9944
R19302 vdd.n329 vdd.n291 12.8005
R19303 vdd.n324 vdd.n295 12.8005
R19304 vdd.n270 vdd.n232 12.8005
R19305 vdd.n265 vdd.n236 12.8005
R19306 vdd.n227 vdd.n189 12.8005
R19307 vdd.n222 vdd.n193 12.8005
R19308 vdd.n168 vdd.n130 12.8005
R19309 vdd.n163 vdd.n134 12.8005
R19310 vdd.n126 vdd.n88 12.8005
R19311 vdd.n121 vdd.n92 12.8005
R19312 vdd.n67 vdd.n29 12.8005
R19313 vdd.n62 vdd.n33 12.8005
R19314 vdd.n2203 vdd.n2165 12.8005
R19315 vdd.n2198 vdd.n2169 12.8005
R19316 vdd.n2262 vdd.n2224 12.8005
R19317 vdd.n2257 vdd.n2228 12.8005
R19318 vdd.n2101 vdd.n2063 12.8005
R19319 vdd.n2096 vdd.n2067 12.8005
R19320 vdd.n2160 vdd.n2122 12.8005
R19321 vdd.n2155 vdd.n2126 12.8005
R19322 vdd.n2000 vdd.n1962 12.8005
R19323 vdd.n1995 vdd.n1966 12.8005
R19324 vdd.n2059 vdd.n2021 12.8005
R19325 vdd.n2054 vdd.n2025 12.8005
R19326 vdd.n323 vdd.n296 12.0247
R19327 vdd.n264 vdd.n237 12.0247
R19328 vdd.n221 vdd.n194 12.0247
R19329 vdd.n162 vdd.n135 12.0247
R19330 vdd.n120 vdd.n93 12.0247
R19331 vdd.n61 vdd.n34 12.0247
R19332 vdd.n2197 vdd.n2170 12.0247
R19333 vdd.n2256 vdd.n2229 12.0247
R19334 vdd.n2095 vdd.n2068 12.0247
R19335 vdd.n2154 vdd.n2127 12.0247
R19336 vdd.n1994 vdd.n1967 12.0247
R19337 vdd.n2053 vdd.n2026 12.0247
R19338 vdd.n1882 vdd.n1638 11.337
R19339 vdd.n1891 vdd.n1638 11.337
R19340 vdd.n1891 vdd.n1890 11.337
R19341 vdd.n1899 vdd.n1632 11.337
R19342 vdd.n1908 vdd.n1907 11.337
R19343 vdd.n1924 vdd.n1616 11.337
R19344 vdd.n1932 vdd.n1609 11.337
R19345 vdd.n1941 vdd.n1940 11.337
R19346 vdd.n1949 vdd.n1598 11.337
R19347 vdd.n2272 vdd.n1587 11.337
R19348 vdd.n2281 vdd.n1581 11.337
R19349 vdd.n2289 vdd.n1575 11.337
R19350 vdd.n2298 vdd.n2297 11.337
R19351 vdd.n2314 vdd.n1559 11.337
R19352 vdd.n2322 vdd.n1552 11.337
R19353 vdd.n2331 vdd.n2330 11.337
R19354 vdd.n2339 vdd.n1535 11.337
R19355 vdd.n2350 vdd.n1535 11.337
R19356 vdd.n2350 vdd.n2349 11.337
R19357 vdd.n3503 vdd.n678 11.337
R19358 vdd.n3511 vdd.n678 11.337
R19359 vdd.n3511 vdd.n679 11.337
R19360 vdd.n3520 vdd.n3519 11.337
R19361 vdd.n3536 vdd.n662 11.337
R19362 vdd.n3544 vdd.n655 11.337
R19363 vdd.n3553 vdd.n3552 11.337
R19364 vdd.n3561 vdd.n644 11.337
R19365 vdd.n3580 vdd.n633 11.337
R19366 vdd.n3667 vdd.n340 11.337
R19367 vdd.n3665 vdd.n344 11.337
R19368 vdd.n3659 vdd.n3658 11.337
R19369 vdd.n3651 vdd.n361 11.337
R19370 vdd.n3650 vdd.n3649 11.337
R19371 vdd.n3643 vdd.n3642 11.337
R19372 vdd.n3641 vdd.n375 11.337
R19373 vdd.n3635 vdd.n3634 11.337
R19374 vdd.n3634 vdd.n3633 11.337
R19375 vdd.n3633 vdd.n386 11.337
R19376 vdd.n320 vdd.n319 11.249
R19377 vdd.n261 vdd.n260 11.249
R19378 vdd.n218 vdd.n217 11.249
R19379 vdd.n159 vdd.n158 11.249
R19380 vdd.n117 vdd.n116 11.249
R19381 vdd.n58 vdd.n57 11.249
R19382 vdd.n2194 vdd.n2193 11.249
R19383 vdd.n2253 vdd.n2252 11.249
R19384 vdd.n2092 vdd.n2091 11.249
R19385 vdd.n2151 vdd.n2150 11.249
R19386 vdd.n1991 vdd.n1990 11.249
R19387 vdd.n2050 vdd.n2049 11.249
R19388 vdd.n1680 vdd.t147 11.2237
R19389 vdd.n3627 vdd.t96 11.2237
R19390 vdd.t193 vdd.n1553 10.7702
R19391 vdd.n3528 vdd.t62 10.7702
R19392 vdd.n305 vdd.n304 10.7238
R19393 vdd.n246 vdd.n245 10.7238
R19394 vdd.n203 vdd.n202 10.7238
R19395 vdd.n144 vdd.n143 10.7238
R19396 vdd.n102 vdd.n101 10.7238
R19397 vdd.n43 vdd.n42 10.7238
R19398 vdd.n2179 vdd.n2178 10.7238
R19399 vdd.n2238 vdd.n2237 10.7238
R19400 vdd.n2077 vdd.n2076 10.7238
R19401 vdd.n2136 vdd.n2135 10.7238
R19402 vdd.n1976 vdd.n1975 10.7238
R19403 vdd.n2035 vdd.n2034 10.7238
R19404 vdd.n2511 vdd.n2510 10.6151
R19405 vdd.n2511 vdd.n1127 10.6151
R19406 vdd.n2521 vdd.n1127 10.6151
R19407 vdd.n2522 vdd.n2521 10.6151
R19408 vdd.n2523 vdd.n2522 10.6151
R19409 vdd.n2523 vdd.n1114 10.6151
R19410 vdd.n2533 vdd.n1114 10.6151
R19411 vdd.n2534 vdd.n2533 10.6151
R19412 vdd.n2535 vdd.n2534 10.6151
R19413 vdd.n2535 vdd.n1102 10.6151
R19414 vdd.n2545 vdd.n1102 10.6151
R19415 vdd.n2546 vdd.n2545 10.6151
R19416 vdd.n2547 vdd.n2546 10.6151
R19417 vdd.n2547 vdd.n1091 10.6151
R19418 vdd.n2557 vdd.n1091 10.6151
R19419 vdd.n2558 vdd.n2557 10.6151
R19420 vdd.n2559 vdd.n2558 10.6151
R19421 vdd.n2559 vdd.n1078 10.6151
R19422 vdd.n2569 vdd.n1078 10.6151
R19423 vdd.n2570 vdd.n2569 10.6151
R19424 vdd.n2571 vdd.n2570 10.6151
R19425 vdd.n2571 vdd.n1066 10.6151
R19426 vdd.n2582 vdd.n1066 10.6151
R19427 vdd.n2583 vdd.n2582 10.6151
R19428 vdd.n2584 vdd.n2583 10.6151
R19429 vdd.n2584 vdd.n1054 10.6151
R19430 vdd.n2594 vdd.n1054 10.6151
R19431 vdd.n2595 vdd.n2594 10.6151
R19432 vdd.n2596 vdd.n2595 10.6151
R19433 vdd.n2596 vdd.n1042 10.6151
R19434 vdd.n2606 vdd.n1042 10.6151
R19435 vdd.n2607 vdd.n2606 10.6151
R19436 vdd.n2608 vdd.n2607 10.6151
R19437 vdd.n2608 vdd.n1032 10.6151
R19438 vdd.n2618 vdd.n1032 10.6151
R19439 vdd.n2619 vdd.n2618 10.6151
R19440 vdd.n2620 vdd.n2619 10.6151
R19441 vdd.n2620 vdd.n1019 10.6151
R19442 vdd.n2632 vdd.n1019 10.6151
R19443 vdd.n2633 vdd.n2632 10.6151
R19444 vdd.n2635 vdd.n2633 10.6151
R19445 vdd.n2635 vdd.n2634 10.6151
R19446 vdd.n2634 vdd.n1000 10.6151
R19447 vdd.n2782 vdd.n2781 10.6151
R19448 vdd.n2781 vdd.n2780 10.6151
R19449 vdd.n2780 vdd.n2777 10.6151
R19450 vdd.n2777 vdd.n2776 10.6151
R19451 vdd.n2776 vdd.n2773 10.6151
R19452 vdd.n2773 vdd.n2772 10.6151
R19453 vdd.n2772 vdd.n2769 10.6151
R19454 vdd.n2769 vdd.n2768 10.6151
R19455 vdd.n2768 vdd.n2765 10.6151
R19456 vdd.n2765 vdd.n2764 10.6151
R19457 vdd.n2764 vdd.n2761 10.6151
R19458 vdd.n2761 vdd.n2760 10.6151
R19459 vdd.n2760 vdd.n2757 10.6151
R19460 vdd.n2757 vdd.n2756 10.6151
R19461 vdd.n2756 vdd.n2753 10.6151
R19462 vdd.n2753 vdd.n2752 10.6151
R19463 vdd.n2752 vdd.n2749 10.6151
R19464 vdd.n2749 vdd.n2748 10.6151
R19465 vdd.n2748 vdd.n2745 10.6151
R19466 vdd.n2745 vdd.n2744 10.6151
R19467 vdd.n2744 vdd.n2741 10.6151
R19468 vdd.n2741 vdd.n2740 10.6151
R19469 vdd.n2740 vdd.n2737 10.6151
R19470 vdd.n2737 vdd.n2736 10.6151
R19471 vdd.n2736 vdd.n2733 10.6151
R19472 vdd.n2733 vdd.n2732 10.6151
R19473 vdd.n2732 vdd.n2729 10.6151
R19474 vdd.n2729 vdd.n2728 10.6151
R19475 vdd.n2728 vdd.n2725 10.6151
R19476 vdd.n2725 vdd.n2724 10.6151
R19477 vdd.n2724 vdd.n2721 10.6151
R19478 vdd.n2719 vdd.n2716 10.6151
R19479 vdd.n2716 vdd.n2715 10.6151
R19480 vdd.n1357 vdd.n1356 10.6151
R19481 vdd.n1359 vdd.n1357 10.6151
R19482 vdd.n1360 vdd.n1359 10.6151
R19483 vdd.n1362 vdd.n1360 10.6151
R19484 vdd.n1363 vdd.n1362 10.6151
R19485 vdd.n1365 vdd.n1363 10.6151
R19486 vdd.n1366 vdd.n1365 10.6151
R19487 vdd.n1368 vdd.n1366 10.6151
R19488 vdd.n1369 vdd.n1368 10.6151
R19489 vdd.n1371 vdd.n1369 10.6151
R19490 vdd.n1372 vdd.n1371 10.6151
R19491 vdd.n1374 vdd.n1372 10.6151
R19492 vdd.n1375 vdd.n1374 10.6151
R19493 vdd.n1377 vdd.n1375 10.6151
R19494 vdd.n1378 vdd.n1377 10.6151
R19495 vdd.n1380 vdd.n1378 10.6151
R19496 vdd.n1381 vdd.n1380 10.6151
R19497 vdd.n1383 vdd.n1381 10.6151
R19498 vdd.n1384 vdd.n1383 10.6151
R19499 vdd.n1386 vdd.n1384 10.6151
R19500 vdd.n1387 vdd.n1386 10.6151
R19501 vdd.n1389 vdd.n1387 10.6151
R19502 vdd.n1390 vdd.n1389 10.6151
R19503 vdd.n1392 vdd.n1390 10.6151
R19504 vdd.n1393 vdd.n1392 10.6151
R19505 vdd.n1395 vdd.n1393 10.6151
R19506 vdd.n1396 vdd.n1395 10.6151
R19507 vdd.n1435 vdd.n1396 10.6151
R19508 vdd.n1435 vdd.n1434 10.6151
R19509 vdd.n1434 vdd.n1433 10.6151
R19510 vdd.n1433 vdd.n1431 10.6151
R19511 vdd.n1431 vdd.n1430 10.6151
R19512 vdd.n1430 vdd.n1428 10.6151
R19513 vdd.n1428 vdd.n1427 10.6151
R19514 vdd.n1427 vdd.n1408 10.6151
R19515 vdd.n1408 vdd.n1407 10.6151
R19516 vdd.n1407 vdd.n1405 10.6151
R19517 vdd.n1405 vdd.n1404 10.6151
R19518 vdd.n1404 vdd.n1402 10.6151
R19519 vdd.n1402 vdd.n1401 10.6151
R19520 vdd.n1401 vdd.n1398 10.6151
R19521 vdd.n1398 vdd.n1397 10.6151
R19522 vdd.n1397 vdd.n1003 10.6151
R19523 vdd.n2509 vdd.n1139 10.6151
R19524 vdd.n2504 vdd.n1139 10.6151
R19525 vdd.n2504 vdd.n2503 10.6151
R19526 vdd.n2503 vdd.n2502 10.6151
R19527 vdd.n2502 vdd.n2499 10.6151
R19528 vdd.n2499 vdd.n2498 10.6151
R19529 vdd.n2498 vdd.n2495 10.6151
R19530 vdd.n2495 vdd.n2494 10.6151
R19531 vdd.n2494 vdd.n2491 10.6151
R19532 vdd.n2491 vdd.n2490 10.6151
R19533 vdd.n2490 vdd.n2487 10.6151
R19534 vdd.n2487 vdd.n2486 10.6151
R19535 vdd.n2486 vdd.n2483 10.6151
R19536 vdd.n2483 vdd.n2482 10.6151
R19537 vdd.n2482 vdd.n2479 10.6151
R19538 vdd.n2479 vdd.n2478 10.6151
R19539 vdd.n2478 vdd.n2475 10.6151
R19540 vdd.n2475 vdd.n1177 10.6151
R19541 vdd.n1323 vdd.n1177 10.6151
R19542 vdd.n1324 vdd.n1323 10.6151
R19543 vdd.n1327 vdd.n1324 10.6151
R19544 vdd.n1328 vdd.n1327 10.6151
R19545 vdd.n1331 vdd.n1328 10.6151
R19546 vdd.n1332 vdd.n1331 10.6151
R19547 vdd.n1335 vdd.n1332 10.6151
R19548 vdd.n1336 vdd.n1335 10.6151
R19549 vdd.n1339 vdd.n1336 10.6151
R19550 vdd.n1340 vdd.n1339 10.6151
R19551 vdd.n1343 vdd.n1340 10.6151
R19552 vdd.n1344 vdd.n1343 10.6151
R19553 vdd.n1347 vdd.n1344 10.6151
R19554 vdd.n1352 vdd.n1349 10.6151
R19555 vdd.n1353 vdd.n1352 10.6151
R19556 vdd.n3020 vdd.n3019 10.6151
R19557 vdd.n3019 vdd.n3018 10.6151
R19558 vdd.n3018 vdd.n2822 10.6151
R19559 vdd.n2900 vdd.n2822 10.6151
R19560 vdd.n2901 vdd.n2900 10.6151
R19561 vdd.n2903 vdd.n2901 10.6151
R19562 vdd.n2904 vdd.n2903 10.6151
R19563 vdd.n3002 vdd.n2904 10.6151
R19564 vdd.n3002 vdd.n3001 10.6151
R19565 vdd.n3001 vdd.n3000 10.6151
R19566 vdd.n3000 vdd.n2948 10.6151
R19567 vdd.n2948 vdd.n2947 10.6151
R19568 vdd.n2947 vdd.n2945 10.6151
R19569 vdd.n2945 vdd.n2944 10.6151
R19570 vdd.n2944 vdd.n2942 10.6151
R19571 vdd.n2942 vdd.n2941 10.6151
R19572 vdd.n2941 vdd.n2939 10.6151
R19573 vdd.n2939 vdd.n2938 10.6151
R19574 vdd.n2938 vdd.n2936 10.6151
R19575 vdd.n2936 vdd.n2935 10.6151
R19576 vdd.n2935 vdd.n2933 10.6151
R19577 vdd.n2933 vdd.n2932 10.6151
R19578 vdd.n2932 vdd.n2930 10.6151
R19579 vdd.n2930 vdd.n2929 10.6151
R19580 vdd.n2929 vdd.n2927 10.6151
R19581 vdd.n2927 vdd.n2926 10.6151
R19582 vdd.n2926 vdd.n2924 10.6151
R19583 vdd.n2924 vdd.n2923 10.6151
R19584 vdd.n2923 vdd.n2921 10.6151
R19585 vdd.n2921 vdd.n2920 10.6151
R19586 vdd.n2920 vdd.n2918 10.6151
R19587 vdd.n2918 vdd.n2917 10.6151
R19588 vdd.n2917 vdd.n2915 10.6151
R19589 vdd.n2915 vdd.n2914 10.6151
R19590 vdd.n2914 vdd.n2912 10.6151
R19591 vdd.n2912 vdd.n2911 10.6151
R19592 vdd.n2911 vdd.n2909 10.6151
R19593 vdd.n2909 vdd.n2908 10.6151
R19594 vdd.n2908 vdd.n2906 10.6151
R19595 vdd.n2906 vdd.n2905 10.6151
R19596 vdd.n2905 vdd.n836 10.6151
R19597 vdd.n3264 vdd.n836 10.6151
R19598 vdd.n3265 vdd.n3264 10.6151
R19599 vdd.n3091 vdd.n961 10.6151
R19600 vdd.n3086 vdd.n961 10.6151
R19601 vdd.n3086 vdd.n3085 10.6151
R19602 vdd.n3085 vdd.n3084 10.6151
R19603 vdd.n3084 vdd.n3081 10.6151
R19604 vdd.n3081 vdd.n3080 10.6151
R19605 vdd.n3080 vdd.n3077 10.6151
R19606 vdd.n3077 vdd.n3076 10.6151
R19607 vdd.n3076 vdd.n3073 10.6151
R19608 vdd.n3073 vdd.n3072 10.6151
R19609 vdd.n3072 vdd.n3069 10.6151
R19610 vdd.n3069 vdd.n3068 10.6151
R19611 vdd.n3068 vdd.n3065 10.6151
R19612 vdd.n3065 vdd.n3064 10.6151
R19613 vdd.n3064 vdd.n3061 10.6151
R19614 vdd.n3061 vdd.n3060 10.6151
R19615 vdd.n3060 vdd.n3057 10.6151
R19616 vdd.n3057 vdd.n3056 10.6151
R19617 vdd.n3056 vdd.n3053 10.6151
R19618 vdd.n3053 vdd.n3052 10.6151
R19619 vdd.n3052 vdd.n3049 10.6151
R19620 vdd.n3049 vdd.n3048 10.6151
R19621 vdd.n3048 vdd.n3045 10.6151
R19622 vdd.n3045 vdd.n3044 10.6151
R19623 vdd.n3044 vdd.n3041 10.6151
R19624 vdd.n3041 vdd.n3040 10.6151
R19625 vdd.n3040 vdd.n3037 10.6151
R19626 vdd.n3037 vdd.n3036 10.6151
R19627 vdd.n3036 vdd.n3033 10.6151
R19628 vdd.n3033 vdd.n3032 10.6151
R19629 vdd.n3032 vdd.n3029 10.6151
R19630 vdd.n3027 vdd.n3024 10.6151
R19631 vdd.n3024 vdd.n3023 10.6151
R19632 vdd.n3093 vdd.n3092 10.6151
R19633 vdd.n3093 vdd.n950 10.6151
R19634 vdd.n3103 vdd.n950 10.6151
R19635 vdd.n3104 vdd.n3103 10.6151
R19636 vdd.n3105 vdd.n3104 10.6151
R19637 vdd.n3105 vdd.n938 10.6151
R19638 vdd.n3115 vdd.n938 10.6151
R19639 vdd.n3116 vdd.n3115 10.6151
R19640 vdd.n3117 vdd.n3116 10.6151
R19641 vdd.n3117 vdd.n927 10.6151
R19642 vdd.n3127 vdd.n927 10.6151
R19643 vdd.n3128 vdd.n3127 10.6151
R19644 vdd.n3129 vdd.n3128 10.6151
R19645 vdd.n3129 vdd.n916 10.6151
R19646 vdd.n3139 vdd.n916 10.6151
R19647 vdd.n3140 vdd.n3139 10.6151
R19648 vdd.n3141 vdd.n3140 10.6151
R19649 vdd.n3141 vdd.n903 10.6151
R19650 vdd.n3152 vdd.n903 10.6151
R19651 vdd.n3153 vdd.n3152 10.6151
R19652 vdd.n3154 vdd.n3153 10.6151
R19653 vdd.n3154 vdd.n891 10.6151
R19654 vdd.n3164 vdd.n891 10.6151
R19655 vdd.n3165 vdd.n3164 10.6151
R19656 vdd.n3166 vdd.n3165 10.6151
R19657 vdd.n3166 vdd.n879 10.6151
R19658 vdd.n3176 vdd.n879 10.6151
R19659 vdd.n3177 vdd.n3176 10.6151
R19660 vdd.n3178 vdd.n3177 10.6151
R19661 vdd.n3178 vdd.n866 10.6151
R19662 vdd.n3188 vdd.n866 10.6151
R19663 vdd.n3189 vdd.n3188 10.6151
R19664 vdd.n3190 vdd.n3189 10.6151
R19665 vdd.n3190 vdd.n855 10.6151
R19666 vdd.n3200 vdd.n855 10.6151
R19667 vdd.n3201 vdd.n3200 10.6151
R19668 vdd.n3202 vdd.n3201 10.6151
R19669 vdd.n3202 vdd.n841 10.6151
R19670 vdd.n3257 vdd.n841 10.6151
R19671 vdd.n3258 vdd.n3257 10.6151
R19672 vdd.n3259 vdd.n3258 10.6151
R19673 vdd.n3259 vdd.n810 10.6151
R19674 vdd.n3329 vdd.n810 10.6151
R19675 vdd.n3328 vdd.n3327 10.6151
R19676 vdd.n3327 vdd.n811 10.6151
R19677 vdd.n812 vdd.n811 10.6151
R19678 vdd.n3320 vdd.n812 10.6151
R19679 vdd.n3320 vdd.n3319 10.6151
R19680 vdd.n3319 vdd.n3318 10.6151
R19681 vdd.n3318 vdd.n814 10.6151
R19682 vdd.n3313 vdd.n814 10.6151
R19683 vdd.n3313 vdd.n3312 10.6151
R19684 vdd.n3312 vdd.n3311 10.6151
R19685 vdd.n3311 vdd.n817 10.6151
R19686 vdd.n3306 vdd.n817 10.6151
R19687 vdd.n3306 vdd.n3305 10.6151
R19688 vdd.n3305 vdd.n3304 10.6151
R19689 vdd.n3304 vdd.n820 10.6151
R19690 vdd.n3299 vdd.n820 10.6151
R19691 vdd.n3299 vdd.n731 10.6151
R19692 vdd.n3295 vdd.n731 10.6151
R19693 vdd.n3295 vdd.n3294 10.6151
R19694 vdd.n3294 vdd.n3293 10.6151
R19695 vdd.n3293 vdd.n823 10.6151
R19696 vdd.n3288 vdd.n823 10.6151
R19697 vdd.n3288 vdd.n3287 10.6151
R19698 vdd.n3287 vdd.n3286 10.6151
R19699 vdd.n3286 vdd.n826 10.6151
R19700 vdd.n3281 vdd.n826 10.6151
R19701 vdd.n3281 vdd.n3280 10.6151
R19702 vdd.n3280 vdd.n3279 10.6151
R19703 vdd.n3279 vdd.n829 10.6151
R19704 vdd.n3274 vdd.n829 10.6151
R19705 vdd.n3274 vdd.n3273 10.6151
R19706 vdd.n3271 vdd.n834 10.6151
R19707 vdd.n3266 vdd.n834 10.6151
R19708 vdd.n3247 vdd.n3208 10.6151
R19709 vdd.n3242 vdd.n3208 10.6151
R19710 vdd.n3242 vdd.n3241 10.6151
R19711 vdd.n3241 vdd.n3240 10.6151
R19712 vdd.n3240 vdd.n3210 10.6151
R19713 vdd.n3235 vdd.n3210 10.6151
R19714 vdd.n3235 vdd.n3234 10.6151
R19715 vdd.n3234 vdd.n3233 10.6151
R19716 vdd.n3233 vdd.n3213 10.6151
R19717 vdd.n3228 vdd.n3213 10.6151
R19718 vdd.n3228 vdd.n3227 10.6151
R19719 vdd.n3227 vdd.n3226 10.6151
R19720 vdd.n3226 vdd.n3216 10.6151
R19721 vdd.n3221 vdd.n3216 10.6151
R19722 vdd.n3221 vdd.n3220 10.6151
R19723 vdd.n3220 vdd.n785 10.6151
R19724 vdd.n3364 vdd.n785 10.6151
R19725 vdd.n3364 vdd.n786 10.6151
R19726 vdd.n788 vdd.n786 10.6151
R19727 vdd.n3357 vdd.n788 10.6151
R19728 vdd.n3357 vdd.n3356 10.6151
R19729 vdd.n3356 vdd.n3355 10.6151
R19730 vdd.n3355 vdd.n790 10.6151
R19731 vdd.n3350 vdd.n790 10.6151
R19732 vdd.n3350 vdd.n3349 10.6151
R19733 vdd.n3349 vdd.n3348 10.6151
R19734 vdd.n3348 vdd.n793 10.6151
R19735 vdd.n3343 vdd.n793 10.6151
R19736 vdd.n3343 vdd.n3342 10.6151
R19737 vdd.n3342 vdd.n3341 10.6151
R19738 vdd.n3341 vdd.n796 10.6151
R19739 vdd.n3336 vdd.n3335 10.6151
R19740 vdd.n3335 vdd.n3334 10.6151
R19741 vdd.n2897 vdd.n2896 10.6151
R19742 vdd.n3014 vdd.n2897 10.6151
R19743 vdd.n3014 vdd.n3013 10.6151
R19744 vdd.n3013 vdd.n3012 10.6151
R19745 vdd.n3012 vdd.n3010 10.6151
R19746 vdd.n3010 vdd.n3009 10.6151
R19747 vdd.n3009 vdd.n3007 10.6151
R19748 vdd.n3007 vdd.n3006 10.6151
R19749 vdd.n3006 vdd.n2898 10.6151
R19750 vdd.n2996 vdd.n2898 10.6151
R19751 vdd.n2996 vdd.n2995 10.6151
R19752 vdd.n2995 vdd.n2994 10.6151
R19753 vdd.n2994 vdd.n2992 10.6151
R19754 vdd.n2992 vdd.n2991 10.6151
R19755 vdd.n2991 vdd.n2989 10.6151
R19756 vdd.n2989 vdd.n2988 10.6151
R19757 vdd.n2988 vdd.n2986 10.6151
R19758 vdd.n2986 vdd.n2985 10.6151
R19759 vdd.n2985 vdd.n2983 10.6151
R19760 vdd.n2983 vdd.n2982 10.6151
R19761 vdd.n2982 vdd.n2980 10.6151
R19762 vdd.n2980 vdd.n2979 10.6151
R19763 vdd.n2979 vdd.n2977 10.6151
R19764 vdd.n2977 vdd.n2976 10.6151
R19765 vdd.n2976 vdd.n2974 10.6151
R19766 vdd.n2974 vdd.n2973 10.6151
R19767 vdd.n2973 vdd.n2971 10.6151
R19768 vdd.n2971 vdd.n2970 10.6151
R19769 vdd.n2970 vdd.n2968 10.6151
R19770 vdd.n2968 vdd.n2967 10.6151
R19771 vdd.n2967 vdd.n2965 10.6151
R19772 vdd.n2965 vdd.n2964 10.6151
R19773 vdd.n2964 vdd.n2962 10.6151
R19774 vdd.n2962 vdd.n2961 10.6151
R19775 vdd.n2961 vdd.n2959 10.6151
R19776 vdd.n2959 vdd.n2958 10.6151
R19777 vdd.n2958 vdd.n2956 10.6151
R19778 vdd.n2956 vdd.n2955 10.6151
R19779 vdd.n2955 vdd.n2953 10.6151
R19780 vdd.n2953 vdd.n2952 10.6151
R19781 vdd.n2952 vdd.n2950 10.6151
R19782 vdd.n2950 vdd.n2949 10.6151
R19783 vdd.n2949 vdd.n802 10.6151
R19784 vdd.n2828 vdd.n2827 10.6151
R19785 vdd.n2831 vdd.n2828 10.6151
R19786 vdd.n2832 vdd.n2831 10.6151
R19787 vdd.n2835 vdd.n2832 10.6151
R19788 vdd.n2836 vdd.n2835 10.6151
R19789 vdd.n2839 vdd.n2836 10.6151
R19790 vdd.n2840 vdd.n2839 10.6151
R19791 vdd.n2843 vdd.n2840 10.6151
R19792 vdd.n2844 vdd.n2843 10.6151
R19793 vdd.n2847 vdd.n2844 10.6151
R19794 vdd.n2848 vdd.n2847 10.6151
R19795 vdd.n2851 vdd.n2848 10.6151
R19796 vdd.n2852 vdd.n2851 10.6151
R19797 vdd.n2855 vdd.n2852 10.6151
R19798 vdd.n2856 vdd.n2855 10.6151
R19799 vdd.n2859 vdd.n2856 10.6151
R19800 vdd.n2860 vdd.n2859 10.6151
R19801 vdd.n2863 vdd.n2860 10.6151
R19802 vdd.n2864 vdd.n2863 10.6151
R19803 vdd.n2867 vdd.n2864 10.6151
R19804 vdd.n2868 vdd.n2867 10.6151
R19805 vdd.n2871 vdd.n2868 10.6151
R19806 vdd.n2872 vdd.n2871 10.6151
R19807 vdd.n2875 vdd.n2872 10.6151
R19808 vdd.n2876 vdd.n2875 10.6151
R19809 vdd.n2879 vdd.n2876 10.6151
R19810 vdd.n2880 vdd.n2879 10.6151
R19811 vdd.n2883 vdd.n2880 10.6151
R19812 vdd.n2884 vdd.n2883 10.6151
R19813 vdd.n2887 vdd.n2884 10.6151
R19814 vdd.n2888 vdd.n2887 10.6151
R19815 vdd.n2893 vdd.n2891 10.6151
R19816 vdd.n2894 vdd.n2893 10.6151
R19817 vdd.n3097 vdd.n955 10.6151
R19818 vdd.n3098 vdd.n3097 10.6151
R19819 vdd.n3099 vdd.n3098 10.6151
R19820 vdd.n3099 vdd.n944 10.6151
R19821 vdd.n3109 vdd.n944 10.6151
R19822 vdd.n3110 vdd.n3109 10.6151
R19823 vdd.n3111 vdd.n3110 10.6151
R19824 vdd.n3111 vdd.n933 10.6151
R19825 vdd.n3121 vdd.n933 10.6151
R19826 vdd.n3122 vdd.n3121 10.6151
R19827 vdd.n3123 vdd.n3122 10.6151
R19828 vdd.n3123 vdd.n921 10.6151
R19829 vdd.n3133 vdd.n921 10.6151
R19830 vdd.n3134 vdd.n3133 10.6151
R19831 vdd.n3135 vdd.n3134 10.6151
R19832 vdd.n3135 vdd.n910 10.6151
R19833 vdd.n3145 vdd.n910 10.6151
R19834 vdd.n3146 vdd.n3145 10.6151
R19835 vdd.n3148 vdd.n3146 10.6151
R19836 vdd.n3148 vdd.n3147 10.6151
R19837 vdd.n3159 vdd.n3158 10.6151
R19838 vdd.n3160 vdd.n3159 10.6151
R19839 vdd.n3160 vdd.n885 10.6151
R19840 vdd.n3170 vdd.n885 10.6151
R19841 vdd.n3171 vdd.n3170 10.6151
R19842 vdd.n3172 vdd.n3171 10.6151
R19843 vdd.n3172 vdd.n872 10.6151
R19844 vdd.n3182 vdd.n872 10.6151
R19845 vdd.n3183 vdd.n3182 10.6151
R19846 vdd.n3184 vdd.n3183 10.6151
R19847 vdd.n3184 vdd.n860 10.6151
R19848 vdd.n3194 vdd.n860 10.6151
R19849 vdd.n3195 vdd.n3194 10.6151
R19850 vdd.n3196 vdd.n3195 10.6151
R19851 vdd.n3196 vdd.n849 10.6151
R19852 vdd.n3206 vdd.n849 10.6151
R19853 vdd.n3207 vdd.n3206 10.6151
R19854 vdd.n3253 vdd.n3207 10.6151
R19855 vdd.n3253 vdd.n3252 10.6151
R19856 vdd.n3252 vdd.n3251 10.6151
R19857 vdd.n3251 vdd.n3250 10.6151
R19858 vdd.n3250 vdd.n3248 10.6151
R19859 vdd.n2515 vdd.n1132 10.6151
R19860 vdd.n2516 vdd.n2515 10.6151
R19861 vdd.n2517 vdd.n2516 10.6151
R19862 vdd.n2517 vdd.n1121 10.6151
R19863 vdd.n2527 vdd.n1121 10.6151
R19864 vdd.n2528 vdd.n2527 10.6151
R19865 vdd.n2529 vdd.n2528 10.6151
R19866 vdd.n2529 vdd.n1108 10.6151
R19867 vdd.n2539 vdd.n1108 10.6151
R19868 vdd.n2540 vdd.n2539 10.6151
R19869 vdd.n2541 vdd.n2540 10.6151
R19870 vdd.n2541 vdd.n1097 10.6151
R19871 vdd.n2551 vdd.n1097 10.6151
R19872 vdd.n2552 vdd.n2551 10.6151
R19873 vdd.n2553 vdd.n2552 10.6151
R19874 vdd.n2553 vdd.n1085 10.6151
R19875 vdd.n2563 vdd.n1085 10.6151
R19876 vdd.n2564 vdd.n2563 10.6151
R19877 vdd.n2565 vdd.n2564 10.6151
R19878 vdd.n2565 vdd.n1072 10.6151
R19879 vdd.n2575 vdd.n1072 10.6151
R19880 vdd.n2576 vdd.n2575 10.6151
R19881 vdd.n2578 vdd.n1060 10.6151
R19882 vdd.n2588 vdd.n1060 10.6151
R19883 vdd.n2589 vdd.n2588 10.6151
R19884 vdd.n2590 vdd.n2589 10.6151
R19885 vdd.n2590 vdd.n1048 10.6151
R19886 vdd.n2600 vdd.n1048 10.6151
R19887 vdd.n2601 vdd.n2600 10.6151
R19888 vdd.n2602 vdd.n2601 10.6151
R19889 vdd.n2602 vdd.n1037 10.6151
R19890 vdd.n2612 vdd.n1037 10.6151
R19891 vdd.n2613 vdd.n2612 10.6151
R19892 vdd.n2614 vdd.n2613 10.6151
R19893 vdd.n2614 vdd.n1026 10.6151
R19894 vdd.n2624 vdd.n1026 10.6151
R19895 vdd.n2625 vdd.n2624 10.6151
R19896 vdd.n2628 vdd.n2625 10.6151
R19897 vdd.n2628 vdd.n2627 10.6151
R19898 vdd.n2627 vdd.n2626 10.6151
R19899 vdd.n2626 vdd.n1009 10.6151
R19900 vdd.n2710 vdd.n1009 10.6151
R19901 vdd.n2709 vdd.n2708 10.6151
R19902 vdd.n2708 vdd.n2705 10.6151
R19903 vdd.n2705 vdd.n2704 10.6151
R19904 vdd.n2704 vdd.n2701 10.6151
R19905 vdd.n2701 vdd.n2700 10.6151
R19906 vdd.n2700 vdd.n2697 10.6151
R19907 vdd.n2697 vdd.n2696 10.6151
R19908 vdd.n2696 vdd.n2693 10.6151
R19909 vdd.n2693 vdd.n2692 10.6151
R19910 vdd.n2692 vdd.n2689 10.6151
R19911 vdd.n2689 vdd.n2688 10.6151
R19912 vdd.n2688 vdd.n2685 10.6151
R19913 vdd.n2685 vdd.n2684 10.6151
R19914 vdd.n2684 vdd.n2681 10.6151
R19915 vdd.n2681 vdd.n2680 10.6151
R19916 vdd.n2680 vdd.n2677 10.6151
R19917 vdd.n2677 vdd.n2676 10.6151
R19918 vdd.n2676 vdd.n2673 10.6151
R19919 vdd.n2673 vdd.n2672 10.6151
R19920 vdd.n2672 vdd.n2669 10.6151
R19921 vdd.n2669 vdd.n2668 10.6151
R19922 vdd.n2668 vdd.n2665 10.6151
R19923 vdd.n2665 vdd.n2664 10.6151
R19924 vdd.n2664 vdd.n2661 10.6151
R19925 vdd.n2661 vdd.n2660 10.6151
R19926 vdd.n2660 vdd.n2657 10.6151
R19927 vdd.n2657 vdd.n2656 10.6151
R19928 vdd.n2656 vdd.n2653 10.6151
R19929 vdd.n2653 vdd.n2652 10.6151
R19930 vdd.n2652 vdd.n2649 10.6151
R19931 vdd.n2649 vdd.n2648 10.6151
R19932 vdd.n2645 vdd.n2644 10.6151
R19933 vdd.n2644 vdd.n2642 10.6151
R19934 vdd.n1481 vdd.n1479 10.6151
R19935 vdd.n1479 vdd.n1478 10.6151
R19936 vdd.n1478 vdd.n1476 10.6151
R19937 vdd.n1476 vdd.n1475 10.6151
R19938 vdd.n1475 vdd.n1473 10.6151
R19939 vdd.n1473 vdd.n1472 10.6151
R19940 vdd.n1472 vdd.n1470 10.6151
R19941 vdd.n1470 vdd.n1469 10.6151
R19942 vdd.n1469 vdd.n1467 10.6151
R19943 vdd.n1467 vdd.n1466 10.6151
R19944 vdd.n1466 vdd.n1464 10.6151
R19945 vdd.n1464 vdd.n1463 10.6151
R19946 vdd.n1463 vdd.n1461 10.6151
R19947 vdd.n1461 vdd.n1460 10.6151
R19948 vdd.n1460 vdd.n1458 10.6151
R19949 vdd.n1458 vdd.n1457 10.6151
R19950 vdd.n1457 vdd.n1455 10.6151
R19951 vdd.n1455 vdd.n1454 10.6151
R19952 vdd.n1454 vdd.n1452 10.6151
R19953 vdd.n1452 vdd.n1451 10.6151
R19954 vdd.n1451 vdd.n1449 10.6151
R19955 vdd.n1449 vdd.n1448 10.6151
R19956 vdd.n1448 vdd.n1446 10.6151
R19957 vdd.n1446 vdd.n1445 10.6151
R19958 vdd.n1445 vdd.n1443 10.6151
R19959 vdd.n1443 vdd.n1442 10.6151
R19960 vdd.n1442 vdd.n1440 10.6151
R19961 vdd.n1440 vdd.n1439 10.6151
R19962 vdd.n1439 vdd.n1318 10.6151
R19963 vdd.n1410 vdd.n1318 10.6151
R19964 vdd.n1411 vdd.n1410 10.6151
R19965 vdd.n1413 vdd.n1411 10.6151
R19966 vdd.n1414 vdd.n1413 10.6151
R19967 vdd.n1423 vdd.n1414 10.6151
R19968 vdd.n1423 vdd.n1422 10.6151
R19969 vdd.n1422 vdd.n1421 10.6151
R19970 vdd.n1421 vdd.n1419 10.6151
R19971 vdd.n1419 vdd.n1418 10.6151
R19972 vdd.n1418 vdd.n1416 10.6151
R19973 vdd.n1416 vdd.n1415 10.6151
R19974 vdd.n1415 vdd.n1013 10.6151
R19975 vdd.n2640 vdd.n1013 10.6151
R19976 vdd.n2641 vdd.n2640 10.6151
R19977 vdd.n1282 vdd.n1281 10.6151
R19978 vdd.n1285 vdd.n1282 10.6151
R19979 vdd.n1286 vdd.n1285 10.6151
R19980 vdd.n1289 vdd.n1286 10.6151
R19981 vdd.n1290 vdd.n1289 10.6151
R19982 vdd.n1293 vdd.n1290 10.6151
R19983 vdd.n1294 vdd.n1293 10.6151
R19984 vdd.n1297 vdd.n1294 10.6151
R19985 vdd.n1298 vdd.n1297 10.6151
R19986 vdd.n1301 vdd.n1298 10.6151
R19987 vdd.n1302 vdd.n1301 10.6151
R19988 vdd.n1305 vdd.n1302 10.6151
R19989 vdd.n1306 vdd.n1305 10.6151
R19990 vdd.n1309 vdd.n1306 10.6151
R19991 vdd.n1310 vdd.n1309 10.6151
R19992 vdd.n1313 vdd.n1310 10.6151
R19993 vdd.n1515 vdd.n1313 10.6151
R19994 vdd.n1515 vdd.n1514 10.6151
R19995 vdd.n1514 vdd.n1512 10.6151
R19996 vdd.n1512 vdd.n1509 10.6151
R19997 vdd.n1509 vdd.n1508 10.6151
R19998 vdd.n1508 vdd.n1505 10.6151
R19999 vdd.n1505 vdd.n1504 10.6151
R20000 vdd.n1504 vdd.n1501 10.6151
R20001 vdd.n1501 vdd.n1500 10.6151
R20002 vdd.n1500 vdd.n1497 10.6151
R20003 vdd.n1497 vdd.n1496 10.6151
R20004 vdd.n1496 vdd.n1493 10.6151
R20005 vdd.n1493 vdd.n1492 10.6151
R20006 vdd.n1492 vdd.n1489 10.6151
R20007 vdd.n1489 vdd.n1488 10.6151
R20008 vdd.n1485 vdd.n1484 10.6151
R20009 vdd.n1484 vdd.n1482 10.6151
R20010 vdd.n2306 vdd.t43 10.5435
R20011 vdd.n656 vdd.t24 10.5435
R20012 vdd.n316 vdd.n298 10.4732
R20013 vdd.n257 vdd.n239 10.4732
R20014 vdd.n214 vdd.n196 10.4732
R20015 vdd.n155 vdd.n137 10.4732
R20016 vdd.n113 vdd.n95 10.4732
R20017 vdd.n54 vdd.n36 10.4732
R20018 vdd.n2190 vdd.n2172 10.4732
R20019 vdd.n2249 vdd.n2231 10.4732
R20020 vdd.n2088 vdd.n2070 10.4732
R20021 vdd.n2147 vdd.n2129 10.4732
R20022 vdd.n1987 vdd.n1969 10.4732
R20023 vdd.n2046 vdd.n2028 10.4732
R20024 vdd.t207 vdd.n2280 10.3167
R20025 vdd.n3572 vdd.t159 10.3167
R20026 vdd.n1957 vdd.t179 10.09
R20027 vdd.n3666 vdd.t39 10.09
R20028 vdd.n2475 vdd.n2474 9.98956
R20029 vdd.n3488 vdd.n731 9.98956
R20030 vdd.n3365 vdd.n3364 9.98956
R20031 vdd.n2367 vdd.n1515 9.98956
R20032 vdd.t163 vdd.n1610 9.86327
R20033 vdd.n3657 vdd.t66 9.86327
R20034 vdd.n2712 vdd.t284 9.7499
R20035 vdd.t269 vdd.n957 9.7499
R20036 vdd.n315 vdd.n300 9.69747
R20037 vdd.n256 vdd.n241 9.69747
R20038 vdd.n213 vdd.n198 9.69747
R20039 vdd.n154 vdd.n139 9.69747
R20040 vdd.n112 vdd.n97 9.69747
R20041 vdd.n53 vdd.n38 9.69747
R20042 vdd.n2189 vdd.n2174 9.69747
R20043 vdd.n2248 vdd.n2233 9.69747
R20044 vdd.n2087 vdd.n2072 9.69747
R20045 vdd.n2146 vdd.n2131 9.69747
R20046 vdd.n1986 vdd.n1971 9.69747
R20047 vdd.n2045 vdd.n2030 9.69747
R20048 vdd.n1916 vdd.t58 9.63654
R20049 vdd.n3603 vdd.t0 9.63654
R20050 vdd.n331 vdd.n330 9.45567
R20051 vdd.n272 vdd.n271 9.45567
R20052 vdd.n229 vdd.n228 9.45567
R20053 vdd.n170 vdd.n169 9.45567
R20054 vdd.n128 vdd.n127 9.45567
R20055 vdd.n69 vdd.n68 9.45567
R20056 vdd.n2205 vdd.n2204 9.45567
R20057 vdd.n2264 vdd.n2263 9.45567
R20058 vdd.n2103 vdd.n2102 9.45567
R20059 vdd.n2162 vdd.n2161 9.45567
R20060 vdd.n2002 vdd.n2001 9.45567
R20061 vdd.n2061 vdd.n2060 9.45567
R20062 vdd.n1890 vdd.t37 9.40981
R20063 vdd.n3635 vdd.t184 9.40981
R20064 vdd.n2437 vdd.n1207 9.3005
R20065 vdd.n2436 vdd.n2435 9.3005
R20066 vdd.n1213 vdd.n1212 9.3005
R20067 vdd.n2430 vdd.n1217 9.3005
R20068 vdd.n2429 vdd.n1218 9.3005
R20069 vdd.n2428 vdd.n1219 9.3005
R20070 vdd.n1223 vdd.n1220 9.3005
R20071 vdd.n2423 vdd.n1224 9.3005
R20072 vdd.n2422 vdd.n1225 9.3005
R20073 vdd.n2421 vdd.n1226 9.3005
R20074 vdd.n1230 vdd.n1227 9.3005
R20075 vdd.n2416 vdd.n1231 9.3005
R20076 vdd.n2415 vdd.n1232 9.3005
R20077 vdd.n2414 vdd.n1233 9.3005
R20078 vdd.n1237 vdd.n1234 9.3005
R20079 vdd.n2409 vdd.n1238 9.3005
R20080 vdd.n2408 vdd.n1239 9.3005
R20081 vdd.n2407 vdd.n1240 9.3005
R20082 vdd.n1244 vdd.n1241 9.3005
R20083 vdd.n2402 vdd.n1245 9.3005
R20084 vdd.n2401 vdd.n1246 9.3005
R20085 vdd.n2400 vdd.n2399 9.3005
R20086 vdd.n2398 vdd.n1247 9.3005
R20087 vdd.n2397 vdd.n2396 9.3005
R20088 vdd.n1253 vdd.n1252 9.3005
R20089 vdd.n2391 vdd.n1257 9.3005
R20090 vdd.n2390 vdd.n1258 9.3005
R20091 vdd.n2389 vdd.n1259 9.3005
R20092 vdd.n1263 vdd.n1260 9.3005
R20093 vdd.n2384 vdd.n1264 9.3005
R20094 vdd.n2383 vdd.n1265 9.3005
R20095 vdd.n2382 vdd.n1266 9.3005
R20096 vdd.n1270 vdd.n1267 9.3005
R20097 vdd.n2377 vdd.n1271 9.3005
R20098 vdd.n2376 vdd.n1272 9.3005
R20099 vdd.n2375 vdd.n1273 9.3005
R20100 vdd.n1277 vdd.n1274 9.3005
R20101 vdd.n2370 vdd.n1278 9.3005
R20102 vdd.n2439 vdd.n2438 9.3005
R20103 vdd.n2461 vdd.n1178 9.3005
R20104 vdd.n2460 vdd.n1186 9.3005
R20105 vdd.n1190 vdd.n1187 9.3005
R20106 vdd.n2455 vdd.n1191 9.3005
R20107 vdd.n2454 vdd.n1192 9.3005
R20108 vdd.n2453 vdd.n1193 9.3005
R20109 vdd.n1197 vdd.n1194 9.3005
R20110 vdd.n2448 vdd.n1198 9.3005
R20111 vdd.n2447 vdd.n1199 9.3005
R20112 vdd.n2446 vdd.n1200 9.3005
R20113 vdd.n1204 vdd.n1201 9.3005
R20114 vdd.n2441 vdd.n1205 9.3005
R20115 vdd.n2440 vdd.n1206 9.3005
R20116 vdd.n2473 vdd.n2472 9.3005
R20117 vdd.n1182 vdd.n1181 9.3005
R20118 vdd.n2270 vdd.n2269 9.3005
R20119 vdd.n1579 vdd.n1578 9.3005
R20120 vdd.n2284 vdd.n2283 9.3005
R20121 vdd.n2285 vdd.n1577 9.3005
R20122 vdd.n2287 vdd.n2286 9.3005
R20123 vdd.n1568 vdd.n1567 9.3005
R20124 vdd.n2301 vdd.n2300 9.3005
R20125 vdd.n2302 vdd.n1566 9.3005
R20126 vdd.n2304 vdd.n2303 9.3005
R20127 vdd.n1557 vdd.n1556 9.3005
R20128 vdd.n2317 vdd.n2316 9.3005
R20129 vdd.n2318 vdd.n1555 9.3005
R20130 vdd.n2320 vdd.n2319 9.3005
R20131 vdd.n1545 vdd.n1544 9.3005
R20132 vdd.n2334 vdd.n2333 9.3005
R20133 vdd.n2335 vdd.n1543 9.3005
R20134 vdd.n2337 vdd.n2336 9.3005
R20135 vdd.n1533 vdd.n1532 9.3005
R20136 vdd.n2353 vdd.n2352 9.3005
R20137 vdd.n2354 vdd.n1531 9.3005
R20138 vdd.n2356 vdd.n2355 9.3005
R20139 vdd.n307 vdd.n306 9.3005
R20140 vdd.n302 vdd.n301 9.3005
R20141 vdd.n313 vdd.n312 9.3005
R20142 vdd.n315 vdd.n314 9.3005
R20143 vdd.n298 vdd.n297 9.3005
R20144 vdd.n321 vdd.n320 9.3005
R20145 vdd.n323 vdd.n322 9.3005
R20146 vdd.n295 vdd.n292 9.3005
R20147 vdd.n330 vdd.n329 9.3005
R20148 vdd.n248 vdd.n247 9.3005
R20149 vdd.n243 vdd.n242 9.3005
R20150 vdd.n254 vdd.n253 9.3005
R20151 vdd.n256 vdd.n255 9.3005
R20152 vdd.n239 vdd.n238 9.3005
R20153 vdd.n262 vdd.n261 9.3005
R20154 vdd.n264 vdd.n263 9.3005
R20155 vdd.n236 vdd.n233 9.3005
R20156 vdd.n271 vdd.n270 9.3005
R20157 vdd.n205 vdd.n204 9.3005
R20158 vdd.n200 vdd.n199 9.3005
R20159 vdd.n211 vdd.n210 9.3005
R20160 vdd.n213 vdd.n212 9.3005
R20161 vdd.n196 vdd.n195 9.3005
R20162 vdd.n219 vdd.n218 9.3005
R20163 vdd.n221 vdd.n220 9.3005
R20164 vdd.n193 vdd.n190 9.3005
R20165 vdd.n228 vdd.n227 9.3005
R20166 vdd.n146 vdd.n145 9.3005
R20167 vdd.n141 vdd.n140 9.3005
R20168 vdd.n152 vdd.n151 9.3005
R20169 vdd.n154 vdd.n153 9.3005
R20170 vdd.n137 vdd.n136 9.3005
R20171 vdd.n160 vdd.n159 9.3005
R20172 vdd.n162 vdd.n161 9.3005
R20173 vdd.n134 vdd.n131 9.3005
R20174 vdd.n169 vdd.n168 9.3005
R20175 vdd.n104 vdd.n103 9.3005
R20176 vdd.n99 vdd.n98 9.3005
R20177 vdd.n110 vdd.n109 9.3005
R20178 vdd.n112 vdd.n111 9.3005
R20179 vdd.n95 vdd.n94 9.3005
R20180 vdd.n118 vdd.n117 9.3005
R20181 vdd.n120 vdd.n119 9.3005
R20182 vdd.n92 vdd.n89 9.3005
R20183 vdd.n127 vdd.n126 9.3005
R20184 vdd.n45 vdd.n44 9.3005
R20185 vdd.n40 vdd.n39 9.3005
R20186 vdd.n51 vdd.n50 9.3005
R20187 vdd.n53 vdd.n52 9.3005
R20188 vdd.n36 vdd.n35 9.3005
R20189 vdd.n59 vdd.n58 9.3005
R20190 vdd.n61 vdd.n60 9.3005
R20191 vdd.n33 vdd.n30 9.3005
R20192 vdd.n68 vdd.n67 9.3005
R20193 vdd.n3410 vdd.n3409 9.3005
R20194 vdd.n3413 vdd.n766 9.3005
R20195 vdd.n3414 vdd.n765 9.3005
R20196 vdd.n3417 vdd.n764 9.3005
R20197 vdd.n3418 vdd.n763 9.3005
R20198 vdd.n3421 vdd.n762 9.3005
R20199 vdd.n3422 vdd.n761 9.3005
R20200 vdd.n3425 vdd.n760 9.3005
R20201 vdd.n3426 vdd.n759 9.3005
R20202 vdd.n3429 vdd.n758 9.3005
R20203 vdd.n3430 vdd.n757 9.3005
R20204 vdd.n3433 vdd.n756 9.3005
R20205 vdd.n3434 vdd.n755 9.3005
R20206 vdd.n3437 vdd.n754 9.3005
R20207 vdd.n3438 vdd.n753 9.3005
R20208 vdd.n3441 vdd.n752 9.3005
R20209 vdd.n3442 vdd.n751 9.3005
R20210 vdd.n3445 vdd.n750 9.3005
R20211 vdd.n3446 vdd.n749 9.3005
R20212 vdd.n3449 vdd.n748 9.3005
R20213 vdd.n3453 vdd.n3452 9.3005
R20214 vdd.n3454 vdd.n747 9.3005
R20215 vdd.n3458 vdd.n3455 9.3005
R20216 vdd.n3461 vdd.n746 9.3005
R20217 vdd.n3462 vdd.n745 9.3005
R20218 vdd.n3465 vdd.n744 9.3005
R20219 vdd.n3466 vdd.n743 9.3005
R20220 vdd.n3469 vdd.n742 9.3005
R20221 vdd.n3470 vdd.n741 9.3005
R20222 vdd.n3473 vdd.n740 9.3005
R20223 vdd.n3474 vdd.n739 9.3005
R20224 vdd.n3477 vdd.n738 9.3005
R20225 vdd.n3478 vdd.n737 9.3005
R20226 vdd.n3481 vdd.n736 9.3005
R20227 vdd.n3482 vdd.n735 9.3005
R20228 vdd.n3485 vdd.n730 9.3005
R20229 vdd.n3491 vdd.n727 9.3005
R20230 vdd.n3492 vdd.n726 9.3005
R20231 vdd.n3506 vdd.n3505 9.3005
R20232 vdd.n3507 vdd.n681 9.3005
R20233 vdd.n3509 vdd.n3508 9.3005
R20234 vdd.n671 vdd.n670 9.3005
R20235 vdd.n3523 vdd.n3522 9.3005
R20236 vdd.n3524 vdd.n669 9.3005
R20237 vdd.n3526 vdd.n3525 9.3005
R20238 vdd.n660 vdd.n659 9.3005
R20239 vdd.n3539 vdd.n3538 9.3005
R20240 vdd.n3540 vdd.n658 9.3005
R20241 vdd.n3542 vdd.n3541 9.3005
R20242 vdd.n648 vdd.n647 9.3005
R20243 vdd.n3556 vdd.n3555 9.3005
R20244 vdd.n3557 vdd.n646 9.3005
R20245 vdd.n3559 vdd.n3558 9.3005
R20246 vdd.n637 vdd.n636 9.3005
R20247 vdd.n3575 vdd.n3574 9.3005
R20248 vdd.n3576 vdd.n635 9.3005
R20249 vdd.n3578 vdd.n3577 9.3005
R20250 vdd.n336 vdd.n334 9.3005
R20251 vdd.n683 vdd.n682 9.3005
R20252 vdd.n3670 vdd.n3669 9.3005
R20253 vdd.n337 vdd.n335 9.3005
R20254 vdd.n3663 vdd.n346 9.3005
R20255 vdd.n3662 vdd.n347 9.3005
R20256 vdd.n3661 vdd.n348 9.3005
R20257 vdd.n355 vdd.n349 9.3005
R20258 vdd.n3655 vdd.n356 9.3005
R20259 vdd.n3654 vdd.n357 9.3005
R20260 vdd.n3653 vdd.n358 9.3005
R20261 vdd.n366 vdd.n359 9.3005
R20262 vdd.n3647 vdd.n367 9.3005
R20263 vdd.n3646 vdd.n368 9.3005
R20264 vdd.n3645 vdd.n369 9.3005
R20265 vdd.n377 vdd.n370 9.3005
R20266 vdd.n3639 vdd.n378 9.3005
R20267 vdd.n3638 vdd.n379 9.3005
R20268 vdd.n3637 vdd.n380 9.3005
R20269 vdd.n388 vdd.n381 9.3005
R20270 vdd.n3631 vdd.n389 9.3005
R20271 vdd.n3630 vdd.n390 9.3005
R20272 vdd.n3629 vdd.n391 9.3005
R20273 vdd.n466 vdd.n463 9.3005
R20274 vdd.n470 vdd.n469 9.3005
R20275 vdd.n471 vdd.n462 9.3005
R20276 vdd.n475 vdd.n472 9.3005
R20277 vdd.n476 vdd.n461 9.3005
R20278 vdd.n480 vdd.n479 9.3005
R20279 vdd.n481 vdd.n460 9.3005
R20280 vdd.n485 vdd.n482 9.3005
R20281 vdd.n486 vdd.n459 9.3005
R20282 vdd.n490 vdd.n489 9.3005
R20283 vdd.n491 vdd.n458 9.3005
R20284 vdd.n495 vdd.n492 9.3005
R20285 vdd.n496 vdd.n457 9.3005
R20286 vdd.n500 vdd.n499 9.3005
R20287 vdd.n501 vdd.n456 9.3005
R20288 vdd.n505 vdd.n502 9.3005
R20289 vdd.n506 vdd.n455 9.3005
R20290 vdd.n510 vdd.n509 9.3005
R20291 vdd.n511 vdd.n454 9.3005
R20292 vdd.n515 vdd.n512 9.3005
R20293 vdd.n516 vdd.n451 9.3005
R20294 vdd.n520 vdd.n519 9.3005
R20295 vdd.n521 vdd.n450 9.3005
R20296 vdd.n525 vdd.n522 9.3005
R20297 vdd.n526 vdd.n449 9.3005
R20298 vdd.n530 vdd.n529 9.3005
R20299 vdd.n531 vdd.n448 9.3005
R20300 vdd.n535 vdd.n532 9.3005
R20301 vdd.n536 vdd.n447 9.3005
R20302 vdd.n540 vdd.n539 9.3005
R20303 vdd.n541 vdd.n446 9.3005
R20304 vdd.n545 vdd.n542 9.3005
R20305 vdd.n546 vdd.n445 9.3005
R20306 vdd.n550 vdd.n549 9.3005
R20307 vdd.n551 vdd.n444 9.3005
R20308 vdd.n555 vdd.n552 9.3005
R20309 vdd.n556 vdd.n443 9.3005
R20310 vdd.n560 vdd.n559 9.3005
R20311 vdd.n561 vdd.n442 9.3005
R20312 vdd.n565 vdd.n562 9.3005
R20313 vdd.n566 vdd.n439 9.3005
R20314 vdd.n570 vdd.n569 9.3005
R20315 vdd.n571 vdd.n438 9.3005
R20316 vdd.n575 vdd.n572 9.3005
R20317 vdd.n576 vdd.n437 9.3005
R20318 vdd.n580 vdd.n579 9.3005
R20319 vdd.n581 vdd.n436 9.3005
R20320 vdd.n585 vdd.n582 9.3005
R20321 vdd.n586 vdd.n435 9.3005
R20322 vdd.n590 vdd.n589 9.3005
R20323 vdd.n591 vdd.n434 9.3005
R20324 vdd.n595 vdd.n592 9.3005
R20325 vdd.n596 vdd.n433 9.3005
R20326 vdd.n600 vdd.n599 9.3005
R20327 vdd.n601 vdd.n432 9.3005
R20328 vdd.n605 vdd.n602 9.3005
R20329 vdd.n606 vdd.n431 9.3005
R20330 vdd.n610 vdd.n609 9.3005
R20331 vdd.n611 vdd.n430 9.3005
R20332 vdd.n615 vdd.n612 9.3005
R20333 vdd.n617 vdd.n429 9.3005
R20334 vdd.n619 vdd.n618 9.3005
R20335 vdd.n3623 vdd.n3622 9.3005
R20336 vdd.n465 vdd.n464 9.3005
R20337 vdd.n3501 vdd.n3500 9.3005
R20338 vdd.n676 vdd.n675 9.3005
R20339 vdd.n3514 vdd.n3513 9.3005
R20340 vdd.n3515 vdd.n674 9.3005
R20341 vdd.n3517 vdd.n3516 9.3005
R20342 vdd.n666 vdd.n665 9.3005
R20343 vdd.n3531 vdd.n3530 9.3005
R20344 vdd.n3532 vdd.n664 9.3005
R20345 vdd.n3534 vdd.n3533 9.3005
R20346 vdd.n653 vdd.n652 9.3005
R20347 vdd.n3547 vdd.n3546 9.3005
R20348 vdd.n3548 vdd.n651 9.3005
R20349 vdd.n3550 vdd.n3549 9.3005
R20350 vdd.n642 vdd.n641 9.3005
R20351 vdd.n3564 vdd.n3563 9.3005
R20352 vdd.n3565 vdd.n640 9.3005
R20353 vdd.n3570 vdd.n3566 9.3005
R20354 vdd.n3569 vdd.n3568 9.3005
R20355 vdd.n3567 vdd.n631 9.3005
R20356 vdd.n3583 vdd.n630 9.3005
R20357 vdd.n3585 vdd.n3584 9.3005
R20358 vdd.n3586 vdd.n629 9.3005
R20359 vdd.n3588 vdd.n3587 9.3005
R20360 vdd.n3590 vdd.n628 9.3005
R20361 vdd.n3592 vdd.n3591 9.3005
R20362 vdd.n3593 vdd.n627 9.3005
R20363 vdd.n3595 vdd.n3594 9.3005
R20364 vdd.n3597 vdd.n626 9.3005
R20365 vdd.n3599 vdd.n3598 9.3005
R20366 vdd.n3600 vdd.n625 9.3005
R20367 vdd.n3602 vdd.n3601 9.3005
R20368 vdd.n3605 vdd.n624 9.3005
R20369 vdd.n3607 vdd.n3606 9.3005
R20370 vdd.n3608 vdd.n623 9.3005
R20371 vdd.n3610 vdd.n3609 9.3005
R20372 vdd.n3612 vdd.n622 9.3005
R20373 vdd.n3614 vdd.n3613 9.3005
R20374 vdd.n3615 vdd.n621 9.3005
R20375 vdd.n3617 vdd.n3616 9.3005
R20376 vdd.n3619 vdd.n620 9.3005
R20377 vdd.n3621 vdd.n3620 9.3005
R20378 vdd.n3499 vdd.n686 9.3005
R20379 vdd.n3498 vdd.n3497 9.3005
R20380 vdd.n3367 vdd.n687 9.3005
R20381 vdd.n3376 vdd.n783 9.3005
R20382 vdd.n3379 vdd.n782 9.3005
R20383 vdd.n3380 vdd.n781 9.3005
R20384 vdd.n3383 vdd.n780 9.3005
R20385 vdd.n3384 vdd.n779 9.3005
R20386 vdd.n3387 vdd.n778 9.3005
R20387 vdd.n3388 vdd.n777 9.3005
R20388 vdd.n3391 vdd.n776 9.3005
R20389 vdd.n3392 vdd.n775 9.3005
R20390 vdd.n3395 vdd.n774 9.3005
R20391 vdd.n3396 vdd.n773 9.3005
R20392 vdd.n3399 vdd.n772 9.3005
R20393 vdd.n3400 vdd.n771 9.3005
R20394 vdd.n3403 vdd.n770 9.3005
R20395 vdd.n3407 vdd.n3406 9.3005
R20396 vdd.n3408 vdd.n767 9.3005
R20397 vdd.n2366 vdd.n2365 9.3005
R20398 vdd.n2361 vdd.n1517 9.3005
R20399 vdd.n1885 vdd.n1884 9.3005
R20400 vdd.n1886 vdd.n1640 9.3005
R20401 vdd.n1888 vdd.n1887 9.3005
R20402 vdd.n1630 vdd.n1629 9.3005
R20403 vdd.n1902 vdd.n1901 9.3005
R20404 vdd.n1903 vdd.n1628 9.3005
R20405 vdd.n1905 vdd.n1904 9.3005
R20406 vdd.n1620 vdd.n1619 9.3005
R20407 vdd.n1919 vdd.n1918 9.3005
R20408 vdd.n1920 vdd.n1618 9.3005
R20409 vdd.n1922 vdd.n1921 9.3005
R20410 vdd.n1607 vdd.n1606 9.3005
R20411 vdd.n1935 vdd.n1934 9.3005
R20412 vdd.n1936 vdd.n1605 9.3005
R20413 vdd.n1938 vdd.n1937 9.3005
R20414 vdd.n1596 vdd.n1595 9.3005
R20415 vdd.n1952 vdd.n1951 9.3005
R20416 vdd.n1953 vdd.n1594 9.3005
R20417 vdd.n1955 vdd.n1954 9.3005
R20418 vdd.n1585 vdd.n1584 9.3005
R20419 vdd.n2275 vdd.n2274 9.3005
R20420 vdd.n2276 vdd.n1583 9.3005
R20421 vdd.n2278 vdd.n2277 9.3005
R20422 vdd.n1573 vdd.n1572 9.3005
R20423 vdd.n2292 vdd.n2291 9.3005
R20424 vdd.n2293 vdd.n1571 9.3005
R20425 vdd.n2295 vdd.n2294 9.3005
R20426 vdd.n1563 vdd.n1562 9.3005
R20427 vdd.n2309 vdd.n2308 9.3005
R20428 vdd.n2310 vdd.n1561 9.3005
R20429 vdd.n2312 vdd.n2311 9.3005
R20430 vdd.n1550 vdd.n1549 9.3005
R20431 vdd.n2325 vdd.n2324 9.3005
R20432 vdd.n2326 vdd.n1548 9.3005
R20433 vdd.n2328 vdd.n2327 9.3005
R20434 vdd.n1540 vdd.n1539 9.3005
R20435 vdd.n2342 vdd.n2341 9.3005
R20436 vdd.n2343 vdd.n1537 9.3005
R20437 vdd.n2347 vdd.n2346 9.3005
R20438 vdd.n2345 vdd.n1538 9.3005
R20439 vdd.n2344 vdd.n1528 9.3005
R20440 vdd.n1642 vdd.n1641 9.3005
R20441 vdd.n1778 vdd.n1777 9.3005
R20442 vdd.n1779 vdd.n1768 9.3005
R20443 vdd.n1781 vdd.n1780 9.3005
R20444 vdd.n1782 vdd.n1767 9.3005
R20445 vdd.n1784 vdd.n1783 9.3005
R20446 vdd.n1785 vdd.n1762 9.3005
R20447 vdd.n1787 vdd.n1786 9.3005
R20448 vdd.n1788 vdd.n1761 9.3005
R20449 vdd.n1790 vdd.n1789 9.3005
R20450 vdd.n1791 vdd.n1756 9.3005
R20451 vdd.n1793 vdd.n1792 9.3005
R20452 vdd.n1794 vdd.n1755 9.3005
R20453 vdd.n1796 vdd.n1795 9.3005
R20454 vdd.n1797 vdd.n1750 9.3005
R20455 vdd.n1799 vdd.n1798 9.3005
R20456 vdd.n1800 vdd.n1749 9.3005
R20457 vdd.n1802 vdd.n1801 9.3005
R20458 vdd.n1803 vdd.n1744 9.3005
R20459 vdd.n1805 vdd.n1804 9.3005
R20460 vdd.n1806 vdd.n1743 9.3005
R20461 vdd.n1808 vdd.n1807 9.3005
R20462 vdd.n1812 vdd.n1739 9.3005
R20463 vdd.n1814 vdd.n1813 9.3005
R20464 vdd.n1815 vdd.n1738 9.3005
R20465 vdd.n1817 vdd.n1816 9.3005
R20466 vdd.n1818 vdd.n1733 9.3005
R20467 vdd.n1820 vdd.n1819 9.3005
R20468 vdd.n1821 vdd.n1732 9.3005
R20469 vdd.n1823 vdd.n1822 9.3005
R20470 vdd.n1824 vdd.n1727 9.3005
R20471 vdd.n1826 vdd.n1825 9.3005
R20472 vdd.n1827 vdd.n1726 9.3005
R20473 vdd.n1829 vdd.n1828 9.3005
R20474 vdd.n1830 vdd.n1721 9.3005
R20475 vdd.n1832 vdd.n1831 9.3005
R20476 vdd.n1833 vdd.n1720 9.3005
R20477 vdd.n1835 vdd.n1834 9.3005
R20478 vdd.n1836 vdd.n1715 9.3005
R20479 vdd.n1838 vdd.n1837 9.3005
R20480 vdd.n1839 vdd.n1714 9.3005
R20481 vdd.n1841 vdd.n1840 9.3005
R20482 vdd.n1842 vdd.n1709 9.3005
R20483 vdd.n1844 vdd.n1843 9.3005
R20484 vdd.n1845 vdd.n1708 9.3005
R20485 vdd.n1847 vdd.n1846 9.3005
R20486 vdd.n1848 vdd.n1701 9.3005
R20487 vdd.n1850 vdd.n1849 9.3005
R20488 vdd.n1851 vdd.n1700 9.3005
R20489 vdd.n1853 vdd.n1852 9.3005
R20490 vdd.n1854 vdd.n1695 9.3005
R20491 vdd.n1856 vdd.n1855 9.3005
R20492 vdd.n1857 vdd.n1694 9.3005
R20493 vdd.n1859 vdd.n1858 9.3005
R20494 vdd.n1860 vdd.n1689 9.3005
R20495 vdd.n1862 vdd.n1861 9.3005
R20496 vdd.n1863 vdd.n1688 9.3005
R20497 vdd.n1865 vdd.n1864 9.3005
R20498 vdd.n1866 vdd.n1683 9.3005
R20499 vdd.n1868 vdd.n1867 9.3005
R20500 vdd.n1869 vdd.n1682 9.3005
R20501 vdd.n1871 vdd.n1870 9.3005
R20502 vdd.n1647 vdd.n1646 9.3005
R20503 vdd.n1877 vdd.n1876 9.3005
R20504 vdd.n1776 vdd.n1775 9.3005
R20505 vdd.n1880 vdd.n1879 9.3005
R20506 vdd.n1636 vdd.n1635 9.3005
R20507 vdd.n1894 vdd.n1893 9.3005
R20508 vdd.n1895 vdd.n1634 9.3005
R20509 vdd.n1897 vdd.n1896 9.3005
R20510 vdd.n1625 vdd.n1624 9.3005
R20511 vdd.n1911 vdd.n1910 9.3005
R20512 vdd.n1912 vdd.n1623 9.3005
R20513 vdd.n1914 vdd.n1913 9.3005
R20514 vdd.n1614 vdd.n1613 9.3005
R20515 vdd.n1927 vdd.n1926 9.3005
R20516 vdd.n1928 vdd.n1612 9.3005
R20517 vdd.n1930 vdd.n1929 9.3005
R20518 vdd.n1602 vdd.n1601 9.3005
R20519 vdd.n1944 vdd.n1943 9.3005
R20520 vdd.n1945 vdd.n1600 9.3005
R20521 vdd.n1947 vdd.n1946 9.3005
R20522 vdd.n1591 vdd.n1590 9.3005
R20523 vdd.n1960 vdd.n1959 9.3005
R20524 vdd.n1961 vdd.n1589 9.3005
R20525 vdd.n1878 vdd.n1645 9.3005
R20526 vdd.n2181 vdd.n2180 9.3005
R20527 vdd.n2176 vdd.n2175 9.3005
R20528 vdd.n2187 vdd.n2186 9.3005
R20529 vdd.n2189 vdd.n2188 9.3005
R20530 vdd.n2172 vdd.n2171 9.3005
R20531 vdd.n2195 vdd.n2194 9.3005
R20532 vdd.n2197 vdd.n2196 9.3005
R20533 vdd.n2169 vdd.n2166 9.3005
R20534 vdd.n2204 vdd.n2203 9.3005
R20535 vdd.n2240 vdd.n2239 9.3005
R20536 vdd.n2235 vdd.n2234 9.3005
R20537 vdd.n2246 vdd.n2245 9.3005
R20538 vdd.n2248 vdd.n2247 9.3005
R20539 vdd.n2231 vdd.n2230 9.3005
R20540 vdd.n2254 vdd.n2253 9.3005
R20541 vdd.n2256 vdd.n2255 9.3005
R20542 vdd.n2228 vdd.n2225 9.3005
R20543 vdd.n2263 vdd.n2262 9.3005
R20544 vdd.n2079 vdd.n2078 9.3005
R20545 vdd.n2074 vdd.n2073 9.3005
R20546 vdd.n2085 vdd.n2084 9.3005
R20547 vdd.n2087 vdd.n2086 9.3005
R20548 vdd.n2070 vdd.n2069 9.3005
R20549 vdd.n2093 vdd.n2092 9.3005
R20550 vdd.n2095 vdd.n2094 9.3005
R20551 vdd.n2067 vdd.n2064 9.3005
R20552 vdd.n2102 vdd.n2101 9.3005
R20553 vdd.n2138 vdd.n2137 9.3005
R20554 vdd.n2133 vdd.n2132 9.3005
R20555 vdd.n2144 vdd.n2143 9.3005
R20556 vdd.n2146 vdd.n2145 9.3005
R20557 vdd.n2129 vdd.n2128 9.3005
R20558 vdd.n2152 vdd.n2151 9.3005
R20559 vdd.n2154 vdd.n2153 9.3005
R20560 vdd.n2126 vdd.n2123 9.3005
R20561 vdd.n2161 vdd.n2160 9.3005
R20562 vdd.n1978 vdd.n1977 9.3005
R20563 vdd.n1973 vdd.n1972 9.3005
R20564 vdd.n1984 vdd.n1983 9.3005
R20565 vdd.n1986 vdd.n1985 9.3005
R20566 vdd.n1969 vdd.n1968 9.3005
R20567 vdd.n1992 vdd.n1991 9.3005
R20568 vdd.n1994 vdd.n1993 9.3005
R20569 vdd.n1966 vdd.n1963 9.3005
R20570 vdd.n2001 vdd.n2000 9.3005
R20571 vdd.n2037 vdd.n2036 9.3005
R20572 vdd.n2032 vdd.n2031 9.3005
R20573 vdd.n2043 vdd.n2042 9.3005
R20574 vdd.n2045 vdd.n2044 9.3005
R20575 vdd.n2028 vdd.n2027 9.3005
R20576 vdd.n2051 vdd.n2050 9.3005
R20577 vdd.n2053 vdd.n2052 9.3005
R20578 vdd.n2025 vdd.n2022 9.3005
R20579 vdd.n2060 vdd.n2059 9.3005
R20580 vdd.n1916 vdd.t79 9.18308
R20581 vdd.n3603 vdd.t2 9.18308
R20582 vdd.n1610 vdd.t203 8.95635
R20583 vdd.n2358 vdd.t92 8.95635
R20584 vdd.n723 vdd.t109 8.95635
R20585 vdd.t51 vdd.n3657 8.95635
R20586 vdd.n312 vdd.n311 8.92171
R20587 vdd.n253 vdd.n252 8.92171
R20588 vdd.n210 vdd.n209 8.92171
R20589 vdd.n151 vdd.n150 8.92171
R20590 vdd.n109 vdd.n108 8.92171
R20591 vdd.n50 vdd.n49 8.92171
R20592 vdd.n2186 vdd.n2185 8.92171
R20593 vdd.n2245 vdd.n2244 8.92171
R20594 vdd.n2084 vdd.n2083 8.92171
R20595 vdd.n2143 vdd.n2142 8.92171
R20596 vdd.n1983 vdd.n1982 8.92171
R20597 vdd.n2042 vdd.n2041 8.92171
R20598 vdd.n231 vdd.n129 8.81535
R20599 vdd.n2164 vdd.n2062 8.81535
R20600 vdd.n1957 vdd.t75 8.72962
R20601 vdd.t70 vdd.n3666 8.72962
R20602 vdd.n2280 vdd.t167 8.50289
R20603 vdd.n3572 vdd.t77 8.50289
R20604 vdd.n28 vdd.n14 8.42249
R20605 vdd.n2306 vdd.t56 8.27616
R20606 vdd.t222 vdd.n656 8.27616
R20607 vdd.n3672 vdd.n3671 8.16225
R20608 vdd.n2268 vdd.n2267 8.16225
R20609 vdd.n308 vdd.n302 8.14595
R20610 vdd.n249 vdd.n243 8.14595
R20611 vdd.n206 vdd.n200 8.14595
R20612 vdd.n147 vdd.n141 8.14595
R20613 vdd.n105 vdd.n99 8.14595
R20614 vdd.n46 vdd.n40 8.14595
R20615 vdd.n2182 vdd.n2176 8.14595
R20616 vdd.n2241 vdd.n2235 8.14595
R20617 vdd.n2080 vdd.n2074 8.14595
R20618 vdd.n2139 vdd.n2133 8.14595
R20619 vdd.n1979 vdd.n1973 8.14595
R20620 vdd.n2038 vdd.n2032 8.14595
R20621 vdd.n1553 vdd.t35 8.04943
R20622 vdd.n3528 vdd.t27 8.04943
R20623 vdd.n2513 vdd.n1134 7.70933
R20624 vdd.n2513 vdd.n1137 7.70933
R20625 vdd.n2519 vdd.n1123 7.70933
R20626 vdd.n2525 vdd.n1123 7.70933
R20627 vdd.n2525 vdd.n1116 7.70933
R20628 vdd.n2531 vdd.n1116 7.70933
R20629 vdd.n2531 vdd.n1119 7.70933
R20630 vdd.n2537 vdd.n1112 7.70933
R20631 vdd.n2543 vdd.n1106 7.70933
R20632 vdd.n2549 vdd.n1093 7.70933
R20633 vdd.n2555 vdd.n1093 7.70933
R20634 vdd.n2561 vdd.n1087 7.70933
R20635 vdd.n2567 vdd.n1080 7.70933
R20636 vdd.n2567 vdd.n1083 7.70933
R20637 vdd.n2573 vdd.n1076 7.70933
R20638 vdd.n2580 vdd.n1062 7.70933
R20639 vdd.n2586 vdd.n1062 7.70933
R20640 vdd.n2592 vdd.n1056 7.70933
R20641 vdd.n2598 vdd.n1052 7.70933
R20642 vdd.n2604 vdd.n1046 7.70933
R20643 vdd.n2622 vdd.n1028 7.70933
R20644 vdd.n2622 vdd.n1021 7.70933
R20645 vdd.n2630 vdd.n1021 7.70933
R20646 vdd.n2712 vdd.n1005 7.70933
R20647 vdd.n3095 vdd.n957 7.70933
R20648 vdd.n3107 vdd.n946 7.70933
R20649 vdd.n3107 vdd.n940 7.70933
R20650 vdd.n3113 vdd.n940 7.70933
R20651 vdd.n3125 vdd.n931 7.70933
R20652 vdd.n3131 vdd.n925 7.70933
R20653 vdd.n3143 vdd.n912 7.70933
R20654 vdd.n3150 vdd.n905 7.70933
R20655 vdd.n3150 vdd.n908 7.70933
R20656 vdd.n3156 vdd.n901 7.70933
R20657 vdd.n3162 vdd.n887 7.70933
R20658 vdd.n3168 vdd.n887 7.70933
R20659 vdd.n3174 vdd.n881 7.70933
R20660 vdd.n3180 vdd.n874 7.70933
R20661 vdd.n3180 vdd.n877 7.70933
R20662 vdd.n3186 vdd.n870 7.70933
R20663 vdd.n3192 vdd.n864 7.70933
R20664 vdd.n3198 vdd.n851 7.70933
R20665 vdd.n3204 vdd.n851 7.70933
R20666 vdd.n3204 vdd.n843 7.70933
R20667 vdd.n3255 vdd.n843 7.70933
R20668 vdd.n3255 vdd.n846 7.70933
R20669 vdd.n3261 vdd.n805 7.70933
R20670 vdd.n3331 vdd.n805 7.70933
R20671 vdd.n307 vdd.n304 7.3702
R20672 vdd.n248 vdd.n245 7.3702
R20673 vdd.n205 vdd.n202 7.3702
R20674 vdd.n146 vdd.n143 7.3702
R20675 vdd.n104 vdd.n101 7.3702
R20676 vdd.n45 vdd.n42 7.3702
R20677 vdd.n2181 vdd.n2178 7.3702
R20678 vdd.n2240 vdd.n2237 7.3702
R20679 vdd.n2079 vdd.n2076 7.3702
R20680 vdd.n2138 vdd.n2135 7.3702
R20681 vdd.n1978 vdd.n1975 7.3702
R20682 vdd.n2037 vdd.n2034 7.3702
R20683 vdd.n1106 vdd.t289 7.36923
R20684 vdd.n3186 vdd.t266 7.36923
R20685 vdd.n2339 vdd.t47 7.1425
R20686 vdd.n2537 vdd.t243 7.1425
R20687 vdd.n1425 vdd.t237 7.1425
R20688 vdd.n3119 vdd.t242 7.1425
R20689 vdd.n864 vdd.t252 7.1425
R20690 vdd.n679 vdd.t31 7.1425
R20691 vdd.n1813 vdd.n1812 6.98232
R20692 vdd.n2401 vdd.n2400 6.98232
R20693 vdd.n566 vdd.n565 6.98232
R20694 vdd.n3413 vdd.n3410 6.98232
R20695 vdd.t174 vdd.n1552 6.91577
R20696 vdd.n3536 vdd.t54 6.91577
R20697 vdd.n1425 vdd.t238 6.80241
R20698 vdd.n3119 vdd.t282 6.80241
R20699 vdd.n2298 vdd.t161 6.68904
R20700 vdd.n3552 vdd.t33 6.68904
R20701 vdd.t72 vdd.n1581 6.46231
R20702 vdd.n2561 vdd.t250 6.46231
R20703 vdd.t253 vdd.n1056 6.46231
R20704 vdd.n3143 vdd.t258 6.46231
R20705 vdd.t274 vdd.n881 6.46231
R20706 vdd.n3580 vdd.t170 6.46231
R20707 vdd.n3672 vdd.n333 6.38151
R20708 vdd.n2267 vdd.n2266 6.38151
R20709 vdd.n2637 vdd.t286 6.34895
R20710 vdd.n3016 vdd.t271 6.34895
R20711 vdd.n3158 vdd.n897 6.2444
R20712 vdd.n2577 vdd.n2576 6.2444
R20713 vdd.n1949 vdd.t49 6.23558
R20714 vdd.t29 vdd.n344 6.23558
R20715 vdd.t4 vdd.n1609 6.00885
R20716 vdd.n3651 vdd.t6 6.00885
R20717 vdd.n2598 vdd.t279 5.89549
R20718 vdd.n925 vdd.t254 5.89549
R20719 vdd.n308 vdd.n307 5.81868
R20720 vdd.n249 vdd.n248 5.81868
R20721 vdd.n206 vdd.n205 5.81868
R20722 vdd.n147 vdd.n146 5.81868
R20723 vdd.n105 vdd.n104 5.81868
R20724 vdd.n46 vdd.n45 5.81868
R20725 vdd.n2182 vdd.n2181 5.81868
R20726 vdd.n2241 vdd.n2240 5.81868
R20727 vdd.n2080 vdd.n2079 5.81868
R20728 vdd.n2139 vdd.n2138 5.81868
R20729 vdd.n1979 vdd.n1978 5.81868
R20730 vdd.n2038 vdd.n2037 5.81868
R20731 vdd.n1908 vdd.t45 5.78212
R20732 vdd.n3642 vdd.t186 5.78212
R20733 vdd.n2720 vdd.n2719 5.77611
R20734 vdd.n1349 vdd.n1348 5.77611
R20735 vdd.n3028 vdd.n3027 5.77611
R20736 vdd.n3272 vdd.n3271 5.77611
R20737 vdd.n3336 vdd.n801 5.77611
R20738 vdd.n2891 vdd.n2825 5.77611
R20739 vdd.n2645 vdd.n1012 5.77611
R20740 vdd.n1485 vdd.n1317 5.77611
R20741 vdd.n1775 vdd.n1774 5.62474
R20742 vdd.n2364 vdd.n2361 5.62474
R20743 vdd.n3623 vdd.n428 5.62474
R20744 vdd.n3497 vdd.n690 5.62474
R20745 vdd.n1632 vdd.t45 5.55539
R20746 vdd.n2573 vdd.t268 5.55539
R20747 vdd.n901 vdd.t246 5.55539
R20748 vdd.t186 vdd.n3641 5.55539
R20749 vdd.n1924 vdd.t4 5.32866
R20750 vdd.t6 vdd.n3650 5.32866
R20751 vdd.n1940 vdd.t49 5.10193
R20752 vdd.n3659 vdd.t29 5.10193
R20753 vdd.n311 vdd.n302 5.04292
R20754 vdd.n252 vdd.n243 5.04292
R20755 vdd.n209 vdd.n200 5.04292
R20756 vdd.n150 vdd.n141 5.04292
R20757 vdd.n108 vdd.n99 5.04292
R20758 vdd.n49 vdd.n40 5.04292
R20759 vdd.n2185 vdd.n2176 5.04292
R20760 vdd.n2244 vdd.n2235 5.04292
R20761 vdd.n2083 vdd.n2074 5.04292
R20762 vdd.n2142 vdd.n2133 5.04292
R20763 vdd.n1982 vdd.n1973 5.04292
R20764 vdd.n2041 vdd.n2032 5.04292
R20765 vdd.n2272 vdd.t72 4.8752
R20766 vdd.t249 vdd.t260 4.8752
R20767 vdd.t290 vdd.t236 4.8752
R20768 vdd.t170 vdd.n340 4.8752
R20769 vdd.n2721 vdd.n2720 4.83952
R20770 vdd.n1348 vdd.n1347 4.83952
R20771 vdd.n3029 vdd.n3028 4.83952
R20772 vdd.n3273 vdd.n3272 4.83952
R20773 vdd.n801 vdd.n796 4.83952
R20774 vdd.n2888 vdd.n2825 4.83952
R20775 vdd.n2648 vdd.n1012 4.83952
R20776 vdd.n1488 vdd.n1317 4.83952
R20777 vdd.n1399 vdd.t256 4.76184
R20778 vdd.n3101 vdd.t244 4.76184
R20779 vdd.n2369 vdd.n2368 4.74817
R20780 vdd.n1521 vdd.n1516 4.74817
R20781 vdd.n1183 vdd.n1180 4.74817
R20782 vdd.n2462 vdd.n1179 4.74817
R20783 vdd.n2467 vdd.n1180 4.74817
R20784 vdd.n2466 vdd.n1179 4.74817
R20785 vdd.n3490 vdd.n3489 4.74817
R20786 vdd.n3487 vdd.n3486 4.74817
R20787 vdd.n3487 vdd.n732 4.74817
R20788 vdd.n3489 vdd.n729 4.74817
R20789 vdd.n3372 vdd.n784 4.74817
R20790 vdd.n3368 vdd.n3366 4.74817
R20791 vdd.n3371 vdd.n3366 4.74817
R20792 vdd.n3375 vdd.n784 4.74817
R20793 vdd.n2368 vdd.n1279 4.74817
R20794 vdd.n1518 vdd.n1516 4.74817
R20795 vdd.n333 vdd.n332 4.7074
R20796 vdd.n231 vdd.n230 4.7074
R20797 vdd.n2266 vdd.n2265 4.7074
R20798 vdd.n2164 vdd.n2163 4.7074
R20799 vdd.n1575 vdd.t161 4.64847
R20800 vdd.t251 vdd.n1087 4.64847
R20801 vdd.n2592 vdd.t288 4.64847
R20802 vdd.t277 vdd.n912 4.64847
R20803 vdd.n3174 vdd.t273 4.64847
R20804 vdd.n3561 vdd.t33 4.64847
R20805 vdd.n1076 vdd.t140 4.53511
R20806 vdd.n3156 vdd.t113 4.53511
R20807 vdd.n2314 vdd.t174 4.42174
R20808 vdd.n2519 vdd.t88 4.42174
R20809 vdd.n1399 vdd.t129 4.42174
R20810 vdd.n3101 vdd.t136 4.42174
R20811 vdd.n846 vdd.t84 4.42174
R20812 vdd.t54 vdd.n655 4.42174
R20813 vdd.n3147 vdd.n897 4.37123
R20814 vdd.n2578 vdd.n2577 4.37123
R20815 vdd.n2616 vdd.t275 4.30838
R20816 vdd.n3004 vdd.t262 4.30838
R20817 vdd.n312 vdd.n300 4.26717
R20818 vdd.n253 vdd.n241 4.26717
R20819 vdd.n210 vdd.n198 4.26717
R20820 vdd.n151 vdd.n139 4.26717
R20821 vdd.n109 vdd.n97 4.26717
R20822 vdd.n50 vdd.n38 4.26717
R20823 vdd.n2186 vdd.n2174 4.26717
R20824 vdd.n2245 vdd.n2233 4.26717
R20825 vdd.n2084 vdd.n2072 4.26717
R20826 vdd.n2143 vdd.n2131 4.26717
R20827 vdd.n1983 vdd.n1971 4.26717
R20828 vdd.n2042 vdd.n2030 4.26717
R20829 vdd.n2330 vdd.t47 4.19501
R20830 vdd.n3520 vdd.t31 4.19501
R20831 vdd.n333 vdd.n231 4.10845
R20832 vdd.n2266 vdd.n2164 4.10845
R20833 vdd.n289 vdd.t233 4.06363
R20834 vdd.n289 vdd.t297 4.06363
R20835 vdd.n287 vdd.t42 4.06363
R20836 vdd.n287 vdd.t3 4.06363
R20837 vdd.n285 vdd.t52 4.06363
R20838 vdd.n285 vdd.t67 4.06363
R20839 vdd.n283 vdd.t40 4.06363
R20840 vdd.n283 vdd.t181 4.06363
R20841 vdd.n281 vdd.t191 4.06363
R20842 vdd.n281 vdd.t227 4.06363
R20843 vdd.n279 vdd.t78 4.06363
R20844 vdd.n279 vdd.t160 4.06363
R20845 vdd.n277 vdd.t26 4.06363
R20846 vdd.n277 vdd.t172 4.06363
R20847 vdd.n275 vdd.t55 4.06363
R20848 vdd.n275 vdd.t232 4.06363
R20849 vdd.n273 vdd.t235 4.06363
R20850 vdd.n273 vdd.t178 4.06363
R20851 vdd.n187 vdd.t53 4.06363
R20852 vdd.n187 vdd.t187 4.06363
R20853 vdd.n185 vdd.t64 4.06363
R20854 vdd.n185 vdd.t177 4.06363
R20855 vdd.n183 vdd.t173 4.06363
R20856 vdd.n183 vdd.t82 4.06363
R20857 vdd.n181 vdd.t69 4.06363
R20858 vdd.n181 vdd.t30 4.06363
R20859 vdd.n179 vdd.t300 4.06363
R20860 vdd.n179 vdd.t71 4.06363
R20861 vdd.n177 vdd.t200 4.06363
R20862 vdd.n177 vdd.t218 4.06363
R20863 vdd.n175 vdd.t41 4.06363
R20864 vdd.n175 vdd.t34 4.06363
R20865 vdd.n173 vdd.t74 4.06363
R20866 vdd.n173 vdd.t295 4.06363
R20867 vdd.n171 vdd.t205 4.06363
R20868 vdd.n171 vdd.t63 4.06363
R20869 vdd.n86 vdd.t1 4.06363
R20870 vdd.n86 vdd.t230 4.06363
R20871 vdd.n84 vdd.t7 4.06363
R20872 vdd.n84 vdd.t195 4.06363
R20873 vdd.n82 vdd.t190 4.06363
R20874 vdd.n82 vdd.t234 4.06363
R20875 vdd.n80 vdd.t188 4.06363
R20876 vdd.n80 vdd.t292 4.06363
R20877 vdd.n78 vdd.t171 4.06363
R20878 vdd.n78 vdd.t199 4.06363
R20879 vdd.n76 vdd.t302 4.06363
R20880 vdd.n76 vdd.t231 4.06363
R20881 vdd.n74 vdd.t25 4.06363
R20882 vdd.n74 vdd.t226 4.06363
R20883 vdd.n72 vdd.t197 4.06363
R20884 vdd.n72 vdd.t223 4.06363
R20885 vdd.n70 vdd.t28 4.06363
R20886 vdd.n70 vdd.t294 4.06363
R20887 vdd.n2206 vdd.t298 4.06363
R20888 vdd.n2206 vdd.t36 4.06363
R20889 vdd.n2208 vdd.t57 4.06363
R20890 vdd.n2208 vdd.t306 4.06363
R20891 vdd.n2210 vdd.t213 4.06363
R20892 vdd.n2210 vdd.t215 4.06363
R20893 vdd.n2212 vdd.t304 4.06363
R20894 vdd.n2212 vdd.t307 4.06363
R20895 vdd.n2214 vdd.t198 4.06363
R20896 vdd.n2214 vdd.t224 4.06363
R20897 vdd.n2216 vdd.t201 4.06363
R20898 vdd.n2216 vdd.t180 4.06363
R20899 vdd.n2218 vdd.t303 4.06363
R20900 vdd.n2218 vdd.t219 4.06363
R20901 vdd.n2220 vdd.t217 4.06363
R20902 vdd.n2220 vdd.t299 4.06363
R20903 vdd.n2222 vdd.t216 4.06363
R20904 vdd.n2222 vdd.t59 4.06363
R20905 vdd.n2104 vdd.t194 4.06363
R20906 vdd.n2104 vdd.t183 4.06363
R20907 vdd.n2106 vdd.t209 4.06363
R20908 vdd.n2106 vdd.t175 4.06363
R20909 vdd.n2108 vdd.t162 4.06363
R20910 vdd.n2108 vdd.t61 4.06363
R20911 vdd.n2110 vdd.t212 4.06363
R20912 vdd.n2110 vdd.t176 4.06363
R20913 vdd.n2112 vdd.t196 4.06363
R20914 vdd.n2112 vdd.t73 4.06363
R20915 vdd.n2114 vdd.t50 4.06363
R20916 vdd.n2114 vdd.t301 4.06363
R20917 vdd.n2116 vdd.t164 4.06363
R20918 vdd.n2116 vdd.t204 4.06363
R20919 vdd.n2118 vdd.t228 4.06363
R20920 vdd.n2118 vdd.t182 4.06363
R20921 vdd.n2120 vdd.t46 4.06363
R20922 vdd.n2120 vdd.t296 4.06363
R20923 vdd.n2003 vdd.t293 4.06363
R20924 vdd.n2003 vdd.t68 4.06363
R20925 vdd.n2005 vdd.t221 4.06363
R20926 vdd.n2005 vdd.t214 4.06363
R20927 vdd.n2007 vdd.t192 4.06363
R20928 vdd.n2007 vdd.t44 4.06363
R20929 vdd.n2009 vdd.t208 4.06363
R20930 vdd.n2009 vdd.t168 4.06363
R20931 vdd.n2011 vdd.t76 4.06363
R20932 vdd.n2011 vdd.t169 4.06363
R20933 vdd.n2013 vdd.t229 4.06363
R20934 vdd.n2013 vdd.t189 4.06363
R20935 vdd.n2015 vdd.t220 4.06363
R20936 vdd.n2015 vdd.t305 4.06363
R20937 vdd.n2017 vdd.t80 4.06363
R20938 vdd.n2017 vdd.t5 4.06363
R20939 vdd.n2019 vdd.t206 4.06363
R20940 vdd.n2019 vdd.t166 4.06363
R20941 vdd.n1112 vdd.t281 3.96828
R20942 vdd.n2610 vdd.t259 3.96828
R20943 vdd.n2998 vdd.t278 3.96828
R20944 vdd.n3192 vdd.t267 3.96828
R20945 vdd.n26 vdd.t20 3.9605
R20946 vdd.n26 vdd.t23 3.9605
R20947 vdd.n23 vdd.t19 3.9605
R20948 vdd.n23 vdd.t13 3.9605
R20949 vdd.n21 vdd.t9 3.9605
R20950 vdd.n21 vdd.t18 3.9605
R20951 vdd.n20 vdd.t8 3.9605
R20952 vdd.n20 vdd.t22 3.9605
R20953 vdd.n15 vdd.t14 3.9605
R20954 vdd.n15 vdd.t10 3.9605
R20955 vdd.n16 vdd.t16 3.9605
R20956 vdd.n16 vdd.t11 3.9605
R20957 vdd.n18 vdd.t21 3.9605
R20958 vdd.n18 vdd.t17 3.9605
R20959 vdd.n25 vdd.t12 3.9605
R20960 vdd.n25 vdd.t15 3.9605
R20961 vdd.n2543 vdd.t281 3.74155
R20962 vdd.n1046 vdd.t259 3.74155
R20963 vdd.n3125 vdd.t278 3.74155
R20964 vdd.n870 vdd.t267 3.74155
R20965 vdd.n7 vdd.t291 3.61217
R20966 vdd.n7 vdd.t255 3.61217
R20967 vdd.n8 vdd.t263 3.61217
R20968 vdd.n8 vdd.t283 3.61217
R20969 vdd.n10 vdd.t272 3.61217
R20970 vdd.n10 vdd.t245 3.61217
R20971 vdd.n12 vdd.t241 3.61217
R20972 vdd.n12 vdd.t270 3.61217
R20973 vdd.n5 vdd.t285 3.61217
R20974 vdd.n5 vdd.t265 3.61217
R20975 vdd.n3 vdd.t257 3.61217
R20976 vdd.n3 vdd.t287 3.61217
R20977 vdd.n1 vdd.t239 3.61217
R20978 vdd.n1 vdd.t276 3.61217
R20979 vdd.n0 vdd.t280 3.61217
R20980 vdd.n0 vdd.t261 3.61217
R20981 vdd.n316 vdd.n315 3.49141
R20982 vdd.n257 vdd.n256 3.49141
R20983 vdd.n214 vdd.n213 3.49141
R20984 vdd.n155 vdd.n154 3.49141
R20985 vdd.n113 vdd.n112 3.49141
R20986 vdd.n54 vdd.n53 3.49141
R20987 vdd.n2190 vdd.n2189 3.49141
R20988 vdd.n2249 vdd.n2248 3.49141
R20989 vdd.n2088 vdd.n2087 3.49141
R20990 vdd.n2147 vdd.n2146 3.49141
R20991 vdd.n1987 vdd.n1986 3.49141
R20992 vdd.n2046 vdd.n2045 3.49141
R20993 vdd.t275 vdd.n1028 3.40145
R20994 vdd.n2784 vdd.t284 3.40145
R20995 vdd.n3088 vdd.t269 3.40145
R20996 vdd.n3113 vdd.t262 3.40145
R20997 vdd.n2331 vdd.t35 3.28809
R20998 vdd.n1137 vdd.t88 3.28809
R20999 vdd.n2637 vdd.t129 3.28809
R21000 vdd.n3016 vdd.t136 3.28809
R21001 vdd.n3261 vdd.t84 3.28809
R21002 vdd.n3519 vdd.t27 3.28809
R21003 vdd.t56 vdd.n1559 3.06136
R21004 vdd.n2555 vdd.t251 3.06136
R21005 vdd.n1437 vdd.t288 3.06136
R21006 vdd.n3137 vdd.t277 3.06136
R21007 vdd.t273 vdd.n874 3.06136
R21008 vdd.n3544 vdd.t222 3.06136
R21009 vdd.n2630 vdd.t256 2.94799
R21010 vdd.t244 vdd.n946 2.94799
R21011 vdd.n2289 vdd.t167 2.83463
R21012 vdd.n644 vdd.t77 2.83463
R21013 vdd.n319 vdd.n298 2.71565
R21014 vdd.n260 vdd.n239 2.71565
R21015 vdd.n217 vdd.n196 2.71565
R21016 vdd.n158 vdd.n137 2.71565
R21017 vdd.n116 vdd.n95 2.71565
R21018 vdd.n57 vdd.n36 2.71565
R21019 vdd.n2193 vdd.n2172 2.71565
R21020 vdd.n2252 vdd.n2231 2.71565
R21021 vdd.n2091 vdd.n2070 2.71565
R21022 vdd.n2150 vdd.n2129 2.71565
R21023 vdd.n1990 vdd.n1969 2.71565
R21024 vdd.n2049 vdd.n2028 2.71565
R21025 vdd.t75 vdd.n1587 2.6079
R21026 vdd.n3667 vdd.t70 2.6079
R21027 vdd.n2604 vdd.t260 2.49453
R21028 vdd.n931 vdd.t290 2.49453
R21029 vdd.n306 vdd.n305 2.4129
R21030 vdd.n247 vdd.n246 2.4129
R21031 vdd.n204 vdd.n203 2.4129
R21032 vdd.n145 vdd.n144 2.4129
R21033 vdd.n103 vdd.n102 2.4129
R21034 vdd.n44 vdd.n43 2.4129
R21035 vdd.n2180 vdd.n2179 2.4129
R21036 vdd.n2239 vdd.n2238 2.4129
R21037 vdd.n2078 vdd.n2077 2.4129
R21038 vdd.n2137 vdd.n2136 2.4129
R21039 vdd.n1977 vdd.n1976 2.4129
R21040 vdd.n2036 vdd.n2035 2.4129
R21041 vdd.n1941 vdd.t203 2.38117
R21042 vdd.n2349 vdd.t92 2.38117
R21043 vdd.n3503 vdd.t109 2.38117
R21044 vdd.n3658 vdd.t51 2.38117
R21045 vdd.n2474 vdd.n1180 2.27742
R21046 vdd.n2474 vdd.n1179 2.27742
R21047 vdd.n3488 vdd.n3487 2.27742
R21048 vdd.n3489 vdd.n3488 2.27742
R21049 vdd.n3366 vdd.n3365 2.27742
R21050 vdd.n3365 vdd.n784 2.27742
R21051 vdd.n2368 vdd.n2367 2.27742
R21052 vdd.n2367 vdd.n1516 2.27742
R21053 vdd.t79 vdd.n1616 2.15444
R21054 vdd.n1083 vdd.t268 2.15444
R21055 vdd.n2580 vdd.t248 2.15444
R21056 vdd.n908 vdd.t247 2.15444
R21057 vdd.n3162 vdd.t246 2.15444
R21058 vdd.n3649 vdd.t2 2.15444
R21059 vdd.n320 vdd.n296 1.93989
R21060 vdd.n261 vdd.n237 1.93989
R21061 vdd.n218 vdd.n194 1.93989
R21062 vdd.n159 vdd.n135 1.93989
R21063 vdd.n117 vdd.n93 1.93989
R21064 vdd.n58 vdd.n34 1.93989
R21065 vdd.n2194 vdd.n2170 1.93989
R21066 vdd.n2253 vdd.n2229 1.93989
R21067 vdd.n2092 vdd.n2068 1.93989
R21068 vdd.n2151 vdd.n2127 1.93989
R21069 vdd.n1991 vdd.n1967 1.93989
R21070 vdd.n2050 vdd.n2026 1.93989
R21071 vdd.n1899 vdd.t37 1.92771
R21072 vdd.t184 vdd.n375 1.92771
R21073 vdd.n1437 vdd.t279 1.81434
R21074 vdd.n3137 vdd.t254 1.81434
R21075 vdd.n1907 vdd.t58 1.70098
R21076 vdd.n3643 vdd.t0 1.70098
R21077 vdd.n1932 vdd.t163 1.47425
R21078 vdd.n361 vdd.t66 1.47425
R21079 vdd.t286 vdd.n1005 1.36088
R21080 vdd.n3095 vdd.t271 1.36088
R21081 vdd.n1598 vdd.t179 1.24752
R21082 vdd.t250 vdd.n1080 1.24752
R21083 vdd.n2586 vdd.t253 1.24752
R21084 vdd.t258 vdd.n905 1.24752
R21085 vdd.n3168 vdd.t274 1.24752
R21086 vdd.t39 vdd.n3665 1.24752
R21087 vdd.n2267 vdd.n28 1.21639
R21088 vdd vdd.n3672 1.20856
R21089 vdd.n331 vdd.n291 1.16414
R21090 vdd.n324 vdd.n323 1.16414
R21091 vdd.n272 vdd.n232 1.16414
R21092 vdd.n265 vdd.n264 1.16414
R21093 vdd.n229 vdd.n189 1.16414
R21094 vdd.n222 vdd.n221 1.16414
R21095 vdd.n170 vdd.n130 1.16414
R21096 vdd.n163 vdd.n162 1.16414
R21097 vdd.n128 vdd.n88 1.16414
R21098 vdd.n121 vdd.n120 1.16414
R21099 vdd.n69 vdd.n29 1.16414
R21100 vdd.n62 vdd.n61 1.16414
R21101 vdd.n2205 vdd.n2165 1.16414
R21102 vdd.n2198 vdd.n2197 1.16414
R21103 vdd.n2264 vdd.n2224 1.16414
R21104 vdd.n2257 vdd.n2256 1.16414
R21105 vdd.n2103 vdd.n2063 1.16414
R21106 vdd.n2096 vdd.n2095 1.16414
R21107 vdd.n2162 vdd.n2122 1.16414
R21108 vdd.n2155 vdd.n2154 1.16414
R21109 vdd.n2002 vdd.n1962 1.16414
R21110 vdd.n1995 vdd.n1994 1.16414
R21111 vdd.n2061 vdd.n2021 1.16414
R21112 vdd.n2054 vdd.n2053 1.16414
R21113 vdd.n2281 vdd.t207 1.02079
R21114 vdd.t140 vdd.t248 1.02079
R21115 vdd.t247 vdd.t113 1.02079
R21116 vdd.t159 vdd.n633 1.02079
R21117 vdd.n1778 vdd.n1774 0.970197
R21118 vdd.n2365 vdd.n2364 0.970197
R21119 vdd.n618 vdd.n428 0.970197
R21120 vdd.n3367 vdd.n690 0.970197
R21121 vdd.n2610 vdd.t238 0.907421
R21122 vdd.n2998 vdd.t282 0.907421
R21123 vdd.n2297 vdd.t43 0.794056
R21124 vdd.n3553 vdd.t24 0.794056
R21125 vdd.n2322 vdd.t193 0.567326
R21126 vdd.n1119 vdd.t243 0.567326
R21127 vdd.n2616 vdd.t237 0.567326
R21128 vdd.n3004 vdd.t242 0.567326
R21129 vdd.n3198 vdd.t252 0.567326
R21130 vdd.t62 vdd.n662 0.567326
R21131 vdd.n2355 vdd.n1181 0.530988
R21132 vdd.n726 vdd.n682 0.530988
R21133 vdd.n464 vdd.n391 0.530988
R21134 vdd.n3622 vdd.n3621 0.530988
R21135 vdd.n3499 vdd.n3498 0.530988
R21136 vdd.n2344 vdd.n1517 0.530988
R21137 vdd.n1776 vdd.n1641 0.530988
R21138 vdd.n1878 vdd.n1877 0.530988
R21139 vdd.n4 vdd.n2 0.459552
R21140 vdd.n11 vdd.n9 0.459552
R21141 vdd.n329 vdd.n328 0.388379
R21142 vdd.n295 vdd.n293 0.388379
R21143 vdd.n270 vdd.n269 0.388379
R21144 vdd.n236 vdd.n234 0.388379
R21145 vdd.n227 vdd.n226 0.388379
R21146 vdd.n193 vdd.n191 0.388379
R21147 vdd.n168 vdd.n167 0.388379
R21148 vdd.n134 vdd.n132 0.388379
R21149 vdd.n126 vdd.n125 0.388379
R21150 vdd.n92 vdd.n90 0.388379
R21151 vdd.n67 vdd.n66 0.388379
R21152 vdd.n33 vdd.n31 0.388379
R21153 vdd.n2203 vdd.n2202 0.388379
R21154 vdd.n2169 vdd.n2167 0.388379
R21155 vdd.n2262 vdd.n2261 0.388379
R21156 vdd.n2228 vdd.n2226 0.388379
R21157 vdd.n2101 vdd.n2100 0.388379
R21158 vdd.n2067 vdd.n2065 0.388379
R21159 vdd.n2160 vdd.n2159 0.388379
R21160 vdd.n2126 vdd.n2124 0.388379
R21161 vdd.n2000 vdd.n1999 0.388379
R21162 vdd.n1966 vdd.n1964 0.388379
R21163 vdd.n2059 vdd.n2058 0.388379
R21164 vdd.n2025 vdd.n2023 0.388379
R21165 vdd.n19 vdd.n17 0.387128
R21166 vdd.n24 vdd.n22 0.387128
R21167 vdd.n6 vdd.n4 0.358259
R21168 vdd.n13 vdd.n11 0.358259
R21169 vdd.n276 vdd.n274 0.358259
R21170 vdd.n278 vdd.n276 0.358259
R21171 vdd.n280 vdd.n278 0.358259
R21172 vdd.n282 vdd.n280 0.358259
R21173 vdd.n284 vdd.n282 0.358259
R21174 vdd.n286 vdd.n284 0.358259
R21175 vdd.n288 vdd.n286 0.358259
R21176 vdd.n290 vdd.n288 0.358259
R21177 vdd.n332 vdd.n290 0.358259
R21178 vdd.n174 vdd.n172 0.358259
R21179 vdd.n176 vdd.n174 0.358259
R21180 vdd.n178 vdd.n176 0.358259
R21181 vdd.n180 vdd.n178 0.358259
R21182 vdd.n182 vdd.n180 0.358259
R21183 vdd.n184 vdd.n182 0.358259
R21184 vdd.n186 vdd.n184 0.358259
R21185 vdd.n188 vdd.n186 0.358259
R21186 vdd.n230 vdd.n188 0.358259
R21187 vdd.n73 vdd.n71 0.358259
R21188 vdd.n75 vdd.n73 0.358259
R21189 vdd.n77 vdd.n75 0.358259
R21190 vdd.n79 vdd.n77 0.358259
R21191 vdd.n81 vdd.n79 0.358259
R21192 vdd.n83 vdd.n81 0.358259
R21193 vdd.n85 vdd.n83 0.358259
R21194 vdd.n87 vdd.n85 0.358259
R21195 vdd.n129 vdd.n87 0.358259
R21196 vdd.n2265 vdd.n2223 0.358259
R21197 vdd.n2223 vdd.n2221 0.358259
R21198 vdd.n2221 vdd.n2219 0.358259
R21199 vdd.n2219 vdd.n2217 0.358259
R21200 vdd.n2217 vdd.n2215 0.358259
R21201 vdd.n2215 vdd.n2213 0.358259
R21202 vdd.n2213 vdd.n2211 0.358259
R21203 vdd.n2211 vdd.n2209 0.358259
R21204 vdd.n2209 vdd.n2207 0.358259
R21205 vdd.n2163 vdd.n2121 0.358259
R21206 vdd.n2121 vdd.n2119 0.358259
R21207 vdd.n2119 vdd.n2117 0.358259
R21208 vdd.n2117 vdd.n2115 0.358259
R21209 vdd.n2115 vdd.n2113 0.358259
R21210 vdd.n2113 vdd.n2111 0.358259
R21211 vdd.n2111 vdd.n2109 0.358259
R21212 vdd.n2109 vdd.n2107 0.358259
R21213 vdd.n2107 vdd.n2105 0.358259
R21214 vdd.n2062 vdd.n2020 0.358259
R21215 vdd.n2020 vdd.n2018 0.358259
R21216 vdd.n2018 vdd.n2016 0.358259
R21217 vdd.n2016 vdd.n2014 0.358259
R21218 vdd.n2014 vdd.n2012 0.358259
R21219 vdd.n2012 vdd.n2010 0.358259
R21220 vdd.n2010 vdd.n2008 0.358259
R21221 vdd.n2008 vdd.n2006 0.358259
R21222 vdd.n2006 vdd.n2004 0.358259
R21223 vdd.n2549 vdd.t289 0.340595
R21224 vdd.n1052 vdd.t249 0.340595
R21225 vdd.n3131 vdd.t236 0.340595
R21226 vdd.n877 vdd.t266 0.340595
R21227 vdd.n14 vdd.n6 0.334552
R21228 vdd.n14 vdd.n13 0.334552
R21229 vdd.n27 vdd.n19 0.21707
R21230 vdd.n27 vdd.n24 0.21707
R21231 vdd.n330 vdd.n292 0.155672
R21232 vdd.n322 vdd.n292 0.155672
R21233 vdd.n322 vdd.n321 0.155672
R21234 vdd.n321 vdd.n297 0.155672
R21235 vdd.n314 vdd.n297 0.155672
R21236 vdd.n314 vdd.n313 0.155672
R21237 vdd.n313 vdd.n301 0.155672
R21238 vdd.n306 vdd.n301 0.155672
R21239 vdd.n271 vdd.n233 0.155672
R21240 vdd.n263 vdd.n233 0.155672
R21241 vdd.n263 vdd.n262 0.155672
R21242 vdd.n262 vdd.n238 0.155672
R21243 vdd.n255 vdd.n238 0.155672
R21244 vdd.n255 vdd.n254 0.155672
R21245 vdd.n254 vdd.n242 0.155672
R21246 vdd.n247 vdd.n242 0.155672
R21247 vdd.n228 vdd.n190 0.155672
R21248 vdd.n220 vdd.n190 0.155672
R21249 vdd.n220 vdd.n219 0.155672
R21250 vdd.n219 vdd.n195 0.155672
R21251 vdd.n212 vdd.n195 0.155672
R21252 vdd.n212 vdd.n211 0.155672
R21253 vdd.n211 vdd.n199 0.155672
R21254 vdd.n204 vdd.n199 0.155672
R21255 vdd.n169 vdd.n131 0.155672
R21256 vdd.n161 vdd.n131 0.155672
R21257 vdd.n161 vdd.n160 0.155672
R21258 vdd.n160 vdd.n136 0.155672
R21259 vdd.n153 vdd.n136 0.155672
R21260 vdd.n153 vdd.n152 0.155672
R21261 vdd.n152 vdd.n140 0.155672
R21262 vdd.n145 vdd.n140 0.155672
R21263 vdd.n127 vdd.n89 0.155672
R21264 vdd.n119 vdd.n89 0.155672
R21265 vdd.n119 vdd.n118 0.155672
R21266 vdd.n118 vdd.n94 0.155672
R21267 vdd.n111 vdd.n94 0.155672
R21268 vdd.n111 vdd.n110 0.155672
R21269 vdd.n110 vdd.n98 0.155672
R21270 vdd.n103 vdd.n98 0.155672
R21271 vdd.n68 vdd.n30 0.155672
R21272 vdd.n60 vdd.n30 0.155672
R21273 vdd.n60 vdd.n59 0.155672
R21274 vdd.n59 vdd.n35 0.155672
R21275 vdd.n52 vdd.n35 0.155672
R21276 vdd.n52 vdd.n51 0.155672
R21277 vdd.n51 vdd.n39 0.155672
R21278 vdd.n44 vdd.n39 0.155672
R21279 vdd.n2204 vdd.n2166 0.155672
R21280 vdd.n2196 vdd.n2166 0.155672
R21281 vdd.n2196 vdd.n2195 0.155672
R21282 vdd.n2195 vdd.n2171 0.155672
R21283 vdd.n2188 vdd.n2171 0.155672
R21284 vdd.n2188 vdd.n2187 0.155672
R21285 vdd.n2187 vdd.n2175 0.155672
R21286 vdd.n2180 vdd.n2175 0.155672
R21287 vdd.n2263 vdd.n2225 0.155672
R21288 vdd.n2255 vdd.n2225 0.155672
R21289 vdd.n2255 vdd.n2254 0.155672
R21290 vdd.n2254 vdd.n2230 0.155672
R21291 vdd.n2247 vdd.n2230 0.155672
R21292 vdd.n2247 vdd.n2246 0.155672
R21293 vdd.n2246 vdd.n2234 0.155672
R21294 vdd.n2239 vdd.n2234 0.155672
R21295 vdd.n2102 vdd.n2064 0.155672
R21296 vdd.n2094 vdd.n2064 0.155672
R21297 vdd.n2094 vdd.n2093 0.155672
R21298 vdd.n2093 vdd.n2069 0.155672
R21299 vdd.n2086 vdd.n2069 0.155672
R21300 vdd.n2086 vdd.n2085 0.155672
R21301 vdd.n2085 vdd.n2073 0.155672
R21302 vdd.n2078 vdd.n2073 0.155672
R21303 vdd.n2161 vdd.n2123 0.155672
R21304 vdd.n2153 vdd.n2123 0.155672
R21305 vdd.n2153 vdd.n2152 0.155672
R21306 vdd.n2152 vdd.n2128 0.155672
R21307 vdd.n2145 vdd.n2128 0.155672
R21308 vdd.n2145 vdd.n2144 0.155672
R21309 vdd.n2144 vdd.n2132 0.155672
R21310 vdd.n2137 vdd.n2132 0.155672
R21311 vdd.n2001 vdd.n1963 0.155672
R21312 vdd.n1993 vdd.n1963 0.155672
R21313 vdd.n1993 vdd.n1992 0.155672
R21314 vdd.n1992 vdd.n1968 0.155672
R21315 vdd.n1985 vdd.n1968 0.155672
R21316 vdd.n1985 vdd.n1984 0.155672
R21317 vdd.n1984 vdd.n1972 0.155672
R21318 vdd.n1977 vdd.n1972 0.155672
R21319 vdd.n2060 vdd.n2022 0.155672
R21320 vdd.n2052 vdd.n2022 0.155672
R21321 vdd.n2052 vdd.n2051 0.155672
R21322 vdd.n2051 vdd.n2027 0.155672
R21323 vdd.n2044 vdd.n2027 0.155672
R21324 vdd.n2044 vdd.n2043 0.155672
R21325 vdd.n2043 vdd.n2031 0.155672
R21326 vdd.n2036 vdd.n2031 0.155672
R21327 vdd.n1186 vdd.n1178 0.152939
R21328 vdd.n1190 vdd.n1186 0.152939
R21329 vdd.n1191 vdd.n1190 0.152939
R21330 vdd.n1192 vdd.n1191 0.152939
R21331 vdd.n1193 vdd.n1192 0.152939
R21332 vdd.n1197 vdd.n1193 0.152939
R21333 vdd.n1198 vdd.n1197 0.152939
R21334 vdd.n1199 vdd.n1198 0.152939
R21335 vdd.n1200 vdd.n1199 0.152939
R21336 vdd.n1204 vdd.n1200 0.152939
R21337 vdd.n1205 vdd.n1204 0.152939
R21338 vdd.n1206 vdd.n1205 0.152939
R21339 vdd.n2438 vdd.n1206 0.152939
R21340 vdd.n2438 vdd.n2437 0.152939
R21341 vdd.n2437 vdd.n2436 0.152939
R21342 vdd.n2436 vdd.n1212 0.152939
R21343 vdd.n1217 vdd.n1212 0.152939
R21344 vdd.n1218 vdd.n1217 0.152939
R21345 vdd.n1219 vdd.n1218 0.152939
R21346 vdd.n1223 vdd.n1219 0.152939
R21347 vdd.n1224 vdd.n1223 0.152939
R21348 vdd.n1225 vdd.n1224 0.152939
R21349 vdd.n1226 vdd.n1225 0.152939
R21350 vdd.n1230 vdd.n1226 0.152939
R21351 vdd.n1231 vdd.n1230 0.152939
R21352 vdd.n1232 vdd.n1231 0.152939
R21353 vdd.n1233 vdd.n1232 0.152939
R21354 vdd.n1237 vdd.n1233 0.152939
R21355 vdd.n1238 vdd.n1237 0.152939
R21356 vdd.n1239 vdd.n1238 0.152939
R21357 vdd.n1240 vdd.n1239 0.152939
R21358 vdd.n1244 vdd.n1240 0.152939
R21359 vdd.n1245 vdd.n1244 0.152939
R21360 vdd.n1246 vdd.n1245 0.152939
R21361 vdd.n2399 vdd.n1246 0.152939
R21362 vdd.n2399 vdd.n2398 0.152939
R21363 vdd.n2398 vdd.n2397 0.152939
R21364 vdd.n2397 vdd.n1252 0.152939
R21365 vdd.n1257 vdd.n1252 0.152939
R21366 vdd.n1258 vdd.n1257 0.152939
R21367 vdd.n1259 vdd.n1258 0.152939
R21368 vdd.n1263 vdd.n1259 0.152939
R21369 vdd.n1264 vdd.n1263 0.152939
R21370 vdd.n1265 vdd.n1264 0.152939
R21371 vdd.n1266 vdd.n1265 0.152939
R21372 vdd.n1270 vdd.n1266 0.152939
R21373 vdd.n1271 vdd.n1270 0.152939
R21374 vdd.n1272 vdd.n1271 0.152939
R21375 vdd.n1273 vdd.n1272 0.152939
R21376 vdd.n1277 vdd.n1273 0.152939
R21377 vdd.n1278 vdd.n1277 0.152939
R21378 vdd.n2473 vdd.n1181 0.152939
R21379 vdd.n2269 vdd.n1578 0.152939
R21380 vdd.n2284 vdd.n1578 0.152939
R21381 vdd.n2285 vdd.n2284 0.152939
R21382 vdd.n2286 vdd.n2285 0.152939
R21383 vdd.n2286 vdd.n1567 0.152939
R21384 vdd.n2301 vdd.n1567 0.152939
R21385 vdd.n2302 vdd.n2301 0.152939
R21386 vdd.n2303 vdd.n2302 0.152939
R21387 vdd.n2303 vdd.n1556 0.152939
R21388 vdd.n2317 vdd.n1556 0.152939
R21389 vdd.n2318 vdd.n2317 0.152939
R21390 vdd.n2319 vdd.n2318 0.152939
R21391 vdd.n2319 vdd.n1544 0.152939
R21392 vdd.n2334 vdd.n1544 0.152939
R21393 vdd.n2335 vdd.n2334 0.152939
R21394 vdd.n2336 vdd.n2335 0.152939
R21395 vdd.n2336 vdd.n1532 0.152939
R21396 vdd.n2353 vdd.n1532 0.152939
R21397 vdd.n2354 vdd.n2353 0.152939
R21398 vdd.n2355 vdd.n2354 0.152939
R21399 vdd.n735 vdd.n730 0.152939
R21400 vdd.n736 vdd.n735 0.152939
R21401 vdd.n737 vdd.n736 0.152939
R21402 vdd.n738 vdd.n737 0.152939
R21403 vdd.n739 vdd.n738 0.152939
R21404 vdd.n740 vdd.n739 0.152939
R21405 vdd.n741 vdd.n740 0.152939
R21406 vdd.n742 vdd.n741 0.152939
R21407 vdd.n743 vdd.n742 0.152939
R21408 vdd.n744 vdd.n743 0.152939
R21409 vdd.n745 vdd.n744 0.152939
R21410 vdd.n746 vdd.n745 0.152939
R21411 vdd.n3455 vdd.n746 0.152939
R21412 vdd.n3455 vdd.n3454 0.152939
R21413 vdd.n3454 vdd.n3453 0.152939
R21414 vdd.n3453 vdd.n748 0.152939
R21415 vdd.n749 vdd.n748 0.152939
R21416 vdd.n750 vdd.n749 0.152939
R21417 vdd.n751 vdd.n750 0.152939
R21418 vdd.n752 vdd.n751 0.152939
R21419 vdd.n753 vdd.n752 0.152939
R21420 vdd.n754 vdd.n753 0.152939
R21421 vdd.n755 vdd.n754 0.152939
R21422 vdd.n756 vdd.n755 0.152939
R21423 vdd.n757 vdd.n756 0.152939
R21424 vdd.n758 vdd.n757 0.152939
R21425 vdd.n759 vdd.n758 0.152939
R21426 vdd.n760 vdd.n759 0.152939
R21427 vdd.n761 vdd.n760 0.152939
R21428 vdd.n762 vdd.n761 0.152939
R21429 vdd.n763 vdd.n762 0.152939
R21430 vdd.n764 vdd.n763 0.152939
R21431 vdd.n765 vdd.n764 0.152939
R21432 vdd.n766 vdd.n765 0.152939
R21433 vdd.n3409 vdd.n766 0.152939
R21434 vdd.n3409 vdd.n3408 0.152939
R21435 vdd.n3408 vdd.n3407 0.152939
R21436 vdd.n3407 vdd.n770 0.152939
R21437 vdd.n771 vdd.n770 0.152939
R21438 vdd.n772 vdd.n771 0.152939
R21439 vdd.n773 vdd.n772 0.152939
R21440 vdd.n774 vdd.n773 0.152939
R21441 vdd.n775 vdd.n774 0.152939
R21442 vdd.n776 vdd.n775 0.152939
R21443 vdd.n777 vdd.n776 0.152939
R21444 vdd.n778 vdd.n777 0.152939
R21445 vdd.n779 vdd.n778 0.152939
R21446 vdd.n780 vdd.n779 0.152939
R21447 vdd.n781 vdd.n780 0.152939
R21448 vdd.n782 vdd.n781 0.152939
R21449 vdd.n783 vdd.n782 0.152939
R21450 vdd.n727 vdd.n726 0.152939
R21451 vdd.n3506 vdd.n682 0.152939
R21452 vdd.n3507 vdd.n3506 0.152939
R21453 vdd.n3508 vdd.n3507 0.152939
R21454 vdd.n3508 vdd.n670 0.152939
R21455 vdd.n3523 vdd.n670 0.152939
R21456 vdd.n3524 vdd.n3523 0.152939
R21457 vdd.n3525 vdd.n3524 0.152939
R21458 vdd.n3525 vdd.n659 0.152939
R21459 vdd.n3539 vdd.n659 0.152939
R21460 vdd.n3540 vdd.n3539 0.152939
R21461 vdd.n3541 vdd.n3540 0.152939
R21462 vdd.n3541 vdd.n647 0.152939
R21463 vdd.n3556 vdd.n647 0.152939
R21464 vdd.n3557 vdd.n3556 0.152939
R21465 vdd.n3558 vdd.n3557 0.152939
R21466 vdd.n3558 vdd.n636 0.152939
R21467 vdd.n3575 vdd.n636 0.152939
R21468 vdd.n3576 vdd.n3575 0.152939
R21469 vdd.n3577 vdd.n3576 0.152939
R21470 vdd.n3577 vdd.n334 0.152939
R21471 vdd.n3670 vdd.n335 0.152939
R21472 vdd.n346 vdd.n335 0.152939
R21473 vdd.n347 vdd.n346 0.152939
R21474 vdd.n348 vdd.n347 0.152939
R21475 vdd.n355 vdd.n348 0.152939
R21476 vdd.n356 vdd.n355 0.152939
R21477 vdd.n357 vdd.n356 0.152939
R21478 vdd.n358 vdd.n357 0.152939
R21479 vdd.n366 vdd.n358 0.152939
R21480 vdd.n367 vdd.n366 0.152939
R21481 vdd.n368 vdd.n367 0.152939
R21482 vdd.n369 vdd.n368 0.152939
R21483 vdd.n377 vdd.n369 0.152939
R21484 vdd.n378 vdd.n377 0.152939
R21485 vdd.n379 vdd.n378 0.152939
R21486 vdd.n380 vdd.n379 0.152939
R21487 vdd.n388 vdd.n380 0.152939
R21488 vdd.n389 vdd.n388 0.152939
R21489 vdd.n390 vdd.n389 0.152939
R21490 vdd.n391 vdd.n390 0.152939
R21491 vdd.n464 vdd.n463 0.152939
R21492 vdd.n470 vdd.n463 0.152939
R21493 vdd.n471 vdd.n470 0.152939
R21494 vdd.n472 vdd.n471 0.152939
R21495 vdd.n472 vdd.n461 0.152939
R21496 vdd.n480 vdd.n461 0.152939
R21497 vdd.n481 vdd.n480 0.152939
R21498 vdd.n482 vdd.n481 0.152939
R21499 vdd.n482 vdd.n459 0.152939
R21500 vdd.n490 vdd.n459 0.152939
R21501 vdd.n491 vdd.n490 0.152939
R21502 vdd.n492 vdd.n491 0.152939
R21503 vdd.n492 vdd.n457 0.152939
R21504 vdd.n500 vdd.n457 0.152939
R21505 vdd.n501 vdd.n500 0.152939
R21506 vdd.n502 vdd.n501 0.152939
R21507 vdd.n502 vdd.n455 0.152939
R21508 vdd.n510 vdd.n455 0.152939
R21509 vdd.n511 vdd.n510 0.152939
R21510 vdd.n512 vdd.n511 0.152939
R21511 vdd.n512 vdd.n451 0.152939
R21512 vdd.n520 vdd.n451 0.152939
R21513 vdd.n521 vdd.n520 0.152939
R21514 vdd.n522 vdd.n521 0.152939
R21515 vdd.n522 vdd.n449 0.152939
R21516 vdd.n530 vdd.n449 0.152939
R21517 vdd.n531 vdd.n530 0.152939
R21518 vdd.n532 vdd.n531 0.152939
R21519 vdd.n532 vdd.n447 0.152939
R21520 vdd.n540 vdd.n447 0.152939
R21521 vdd.n541 vdd.n540 0.152939
R21522 vdd.n542 vdd.n541 0.152939
R21523 vdd.n542 vdd.n445 0.152939
R21524 vdd.n550 vdd.n445 0.152939
R21525 vdd.n551 vdd.n550 0.152939
R21526 vdd.n552 vdd.n551 0.152939
R21527 vdd.n552 vdd.n443 0.152939
R21528 vdd.n560 vdd.n443 0.152939
R21529 vdd.n561 vdd.n560 0.152939
R21530 vdd.n562 vdd.n561 0.152939
R21531 vdd.n562 vdd.n439 0.152939
R21532 vdd.n570 vdd.n439 0.152939
R21533 vdd.n571 vdd.n570 0.152939
R21534 vdd.n572 vdd.n571 0.152939
R21535 vdd.n572 vdd.n437 0.152939
R21536 vdd.n580 vdd.n437 0.152939
R21537 vdd.n581 vdd.n580 0.152939
R21538 vdd.n582 vdd.n581 0.152939
R21539 vdd.n582 vdd.n435 0.152939
R21540 vdd.n590 vdd.n435 0.152939
R21541 vdd.n591 vdd.n590 0.152939
R21542 vdd.n592 vdd.n591 0.152939
R21543 vdd.n592 vdd.n433 0.152939
R21544 vdd.n600 vdd.n433 0.152939
R21545 vdd.n601 vdd.n600 0.152939
R21546 vdd.n602 vdd.n601 0.152939
R21547 vdd.n602 vdd.n431 0.152939
R21548 vdd.n610 vdd.n431 0.152939
R21549 vdd.n611 vdd.n610 0.152939
R21550 vdd.n612 vdd.n611 0.152939
R21551 vdd.n612 vdd.n429 0.152939
R21552 vdd.n619 vdd.n429 0.152939
R21553 vdd.n3622 vdd.n619 0.152939
R21554 vdd.n3500 vdd.n3499 0.152939
R21555 vdd.n3500 vdd.n675 0.152939
R21556 vdd.n3514 vdd.n675 0.152939
R21557 vdd.n3515 vdd.n3514 0.152939
R21558 vdd.n3516 vdd.n3515 0.152939
R21559 vdd.n3516 vdd.n665 0.152939
R21560 vdd.n3531 vdd.n665 0.152939
R21561 vdd.n3532 vdd.n3531 0.152939
R21562 vdd.n3533 vdd.n3532 0.152939
R21563 vdd.n3533 vdd.n652 0.152939
R21564 vdd.n3547 vdd.n652 0.152939
R21565 vdd.n3548 vdd.n3547 0.152939
R21566 vdd.n3549 vdd.n3548 0.152939
R21567 vdd.n3549 vdd.n641 0.152939
R21568 vdd.n3564 vdd.n641 0.152939
R21569 vdd.n3565 vdd.n3564 0.152939
R21570 vdd.n3566 vdd.n3565 0.152939
R21571 vdd.n3568 vdd.n3566 0.152939
R21572 vdd.n3568 vdd.n3567 0.152939
R21573 vdd.n3567 vdd.n630 0.152939
R21574 vdd.n3585 vdd.n630 0.152939
R21575 vdd.n3586 vdd.n3585 0.152939
R21576 vdd.n3587 vdd.n3586 0.152939
R21577 vdd.n3587 vdd.n628 0.152939
R21578 vdd.n3592 vdd.n628 0.152939
R21579 vdd.n3593 vdd.n3592 0.152939
R21580 vdd.n3594 vdd.n3593 0.152939
R21581 vdd.n3594 vdd.n626 0.152939
R21582 vdd.n3599 vdd.n626 0.152939
R21583 vdd.n3600 vdd.n3599 0.152939
R21584 vdd.n3601 vdd.n3600 0.152939
R21585 vdd.n3601 vdd.n624 0.152939
R21586 vdd.n3607 vdd.n624 0.152939
R21587 vdd.n3608 vdd.n3607 0.152939
R21588 vdd.n3609 vdd.n3608 0.152939
R21589 vdd.n3609 vdd.n622 0.152939
R21590 vdd.n3614 vdd.n622 0.152939
R21591 vdd.n3615 vdd.n3614 0.152939
R21592 vdd.n3616 vdd.n3615 0.152939
R21593 vdd.n3616 vdd.n620 0.152939
R21594 vdd.n3621 vdd.n620 0.152939
R21595 vdd.n3498 vdd.n687 0.152939
R21596 vdd.n2366 vdd.n1517 0.152939
R21597 vdd.n1885 vdd.n1641 0.152939
R21598 vdd.n1886 vdd.n1885 0.152939
R21599 vdd.n1887 vdd.n1886 0.152939
R21600 vdd.n1887 vdd.n1629 0.152939
R21601 vdd.n1902 vdd.n1629 0.152939
R21602 vdd.n1903 vdd.n1902 0.152939
R21603 vdd.n1904 vdd.n1903 0.152939
R21604 vdd.n1904 vdd.n1619 0.152939
R21605 vdd.n1919 vdd.n1619 0.152939
R21606 vdd.n1920 vdd.n1919 0.152939
R21607 vdd.n1921 vdd.n1920 0.152939
R21608 vdd.n1921 vdd.n1606 0.152939
R21609 vdd.n1935 vdd.n1606 0.152939
R21610 vdd.n1936 vdd.n1935 0.152939
R21611 vdd.n1937 vdd.n1936 0.152939
R21612 vdd.n1937 vdd.n1595 0.152939
R21613 vdd.n1952 vdd.n1595 0.152939
R21614 vdd.n1953 vdd.n1952 0.152939
R21615 vdd.n1954 vdd.n1953 0.152939
R21616 vdd.n1954 vdd.n1584 0.152939
R21617 vdd.n2275 vdd.n1584 0.152939
R21618 vdd.n2276 vdd.n2275 0.152939
R21619 vdd.n2277 vdd.n2276 0.152939
R21620 vdd.n2277 vdd.n1572 0.152939
R21621 vdd.n2292 vdd.n1572 0.152939
R21622 vdd.n2293 vdd.n2292 0.152939
R21623 vdd.n2294 vdd.n2293 0.152939
R21624 vdd.n2294 vdd.n1562 0.152939
R21625 vdd.n2309 vdd.n1562 0.152939
R21626 vdd.n2310 vdd.n2309 0.152939
R21627 vdd.n2311 vdd.n2310 0.152939
R21628 vdd.n2311 vdd.n1549 0.152939
R21629 vdd.n2325 vdd.n1549 0.152939
R21630 vdd.n2326 vdd.n2325 0.152939
R21631 vdd.n2327 vdd.n2326 0.152939
R21632 vdd.n2327 vdd.n1539 0.152939
R21633 vdd.n2342 vdd.n1539 0.152939
R21634 vdd.n2343 vdd.n2342 0.152939
R21635 vdd.n2346 vdd.n2343 0.152939
R21636 vdd.n2346 vdd.n2345 0.152939
R21637 vdd.n2345 vdd.n2344 0.152939
R21638 vdd.n1877 vdd.n1646 0.152939
R21639 vdd.n1870 vdd.n1646 0.152939
R21640 vdd.n1870 vdd.n1869 0.152939
R21641 vdd.n1869 vdd.n1868 0.152939
R21642 vdd.n1868 vdd.n1683 0.152939
R21643 vdd.n1864 vdd.n1683 0.152939
R21644 vdd.n1864 vdd.n1863 0.152939
R21645 vdd.n1863 vdd.n1862 0.152939
R21646 vdd.n1862 vdd.n1689 0.152939
R21647 vdd.n1858 vdd.n1689 0.152939
R21648 vdd.n1858 vdd.n1857 0.152939
R21649 vdd.n1857 vdd.n1856 0.152939
R21650 vdd.n1856 vdd.n1695 0.152939
R21651 vdd.n1852 vdd.n1695 0.152939
R21652 vdd.n1852 vdd.n1851 0.152939
R21653 vdd.n1851 vdd.n1850 0.152939
R21654 vdd.n1850 vdd.n1701 0.152939
R21655 vdd.n1846 vdd.n1701 0.152939
R21656 vdd.n1846 vdd.n1845 0.152939
R21657 vdd.n1845 vdd.n1844 0.152939
R21658 vdd.n1844 vdd.n1709 0.152939
R21659 vdd.n1840 vdd.n1709 0.152939
R21660 vdd.n1840 vdd.n1839 0.152939
R21661 vdd.n1839 vdd.n1838 0.152939
R21662 vdd.n1838 vdd.n1715 0.152939
R21663 vdd.n1834 vdd.n1715 0.152939
R21664 vdd.n1834 vdd.n1833 0.152939
R21665 vdd.n1833 vdd.n1832 0.152939
R21666 vdd.n1832 vdd.n1721 0.152939
R21667 vdd.n1828 vdd.n1721 0.152939
R21668 vdd.n1828 vdd.n1827 0.152939
R21669 vdd.n1827 vdd.n1826 0.152939
R21670 vdd.n1826 vdd.n1727 0.152939
R21671 vdd.n1822 vdd.n1727 0.152939
R21672 vdd.n1822 vdd.n1821 0.152939
R21673 vdd.n1821 vdd.n1820 0.152939
R21674 vdd.n1820 vdd.n1733 0.152939
R21675 vdd.n1816 vdd.n1733 0.152939
R21676 vdd.n1816 vdd.n1815 0.152939
R21677 vdd.n1815 vdd.n1814 0.152939
R21678 vdd.n1814 vdd.n1739 0.152939
R21679 vdd.n1807 vdd.n1739 0.152939
R21680 vdd.n1807 vdd.n1806 0.152939
R21681 vdd.n1806 vdd.n1805 0.152939
R21682 vdd.n1805 vdd.n1744 0.152939
R21683 vdd.n1801 vdd.n1744 0.152939
R21684 vdd.n1801 vdd.n1800 0.152939
R21685 vdd.n1800 vdd.n1799 0.152939
R21686 vdd.n1799 vdd.n1750 0.152939
R21687 vdd.n1795 vdd.n1750 0.152939
R21688 vdd.n1795 vdd.n1794 0.152939
R21689 vdd.n1794 vdd.n1793 0.152939
R21690 vdd.n1793 vdd.n1756 0.152939
R21691 vdd.n1789 vdd.n1756 0.152939
R21692 vdd.n1789 vdd.n1788 0.152939
R21693 vdd.n1788 vdd.n1787 0.152939
R21694 vdd.n1787 vdd.n1762 0.152939
R21695 vdd.n1783 vdd.n1762 0.152939
R21696 vdd.n1783 vdd.n1782 0.152939
R21697 vdd.n1782 vdd.n1781 0.152939
R21698 vdd.n1781 vdd.n1768 0.152939
R21699 vdd.n1777 vdd.n1768 0.152939
R21700 vdd.n1777 vdd.n1776 0.152939
R21701 vdd.n1879 vdd.n1878 0.152939
R21702 vdd.n1879 vdd.n1635 0.152939
R21703 vdd.n1894 vdd.n1635 0.152939
R21704 vdd.n1895 vdd.n1894 0.152939
R21705 vdd.n1896 vdd.n1895 0.152939
R21706 vdd.n1896 vdd.n1624 0.152939
R21707 vdd.n1911 vdd.n1624 0.152939
R21708 vdd.n1912 vdd.n1911 0.152939
R21709 vdd.n1913 vdd.n1912 0.152939
R21710 vdd.n1913 vdd.n1613 0.152939
R21711 vdd.n1927 vdd.n1613 0.152939
R21712 vdd.n1928 vdd.n1927 0.152939
R21713 vdd.n1929 vdd.n1928 0.152939
R21714 vdd.n1929 vdd.n1601 0.152939
R21715 vdd.n1944 vdd.n1601 0.152939
R21716 vdd.n1945 vdd.n1944 0.152939
R21717 vdd.n1946 vdd.n1945 0.152939
R21718 vdd.n1946 vdd.n1590 0.152939
R21719 vdd.n1960 vdd.n1590 0.152939
R21720 vdd.n1961 vdd.n1960 0.152939
R21721 vdd.n1882 vdd.t147 0.113865
R21722 vdd.t96 vdd.n386 0.113865
R21723 vdd.n2474 vdd.n2473 0.110256
R21724 vdd.n3488 vdd.n727 0.110256
R21725 vdd.n3365 vdd.n687 0.110256
R21726 vdd.n2367 vdd.n2366 0.110256
R21727 vdd.n2269 vdd.n2268 0.0695946
R21728 vdd.n3671 vdd.n334 0.0695946
R21729 vdd.n3671 vdd.n3670 0.0695946
R21730 vdd.n2268 vdd.n1961 0.0695946
R21731 vdd.n2474 vdd.n1178 0.0431829
R21732 vdd.n2367 vdd.n1278 0.0431829
R21733 vdd.n3488 vdd.n730 0.0431829
R21734 vdd.n3365 vdd.n783 0.0431829
R21735 vdd vdd.n28 0.00833333
R21736 a_n2804_13878.n2 a_n2804_13878.n0 98.9633
R21737 a_n2804_13878.n5 a_n2804_13878.n3 98.7517
R21738 a_n2804_13878.n25 a_n2804_13878.n24 98.6055
R21739 a_n2804_13878.n27 a_n2804_13878.n26 98.6055
R21740 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R21741 a_n2804_13878.n13 a_n2804_13878.n12 98.6055
R21742 a_n2804_13878.n11 a_n2804_13878.n10 98.6055
R21743 a_n2804_13878.n9 a_n2804_13878.n8 98.6055
R21744 a_n2804_13878.n7 a_n2804_13878.n6 98.6055
R21745 a_n2804_13878.n5 a_n2804_13878.n4 98.6055
R21746 a_n2804_13878.n29 a_n2804_13878.n28 98.6054
R21747 a_n2804_13878.n23 a_n2804_13878.n22 98.6054
R21748 a_n2804_13878.n15 a_n2804_13878.t1 74.6477
R21749 a_n2804_13878.n20 a_n2804_13878.t2 74.2899
R21750 a_n2804_13878.n17 a_n2804_13878.t3 74.2899
R21751 a_n2804_13878.n16 a_n2804_13878.t0 74.2899
R21752 a_n2804_13878.n19 a_n2804_13878.n18 70.6783
R21753 a_n2804_13878.n15 a_n2804_13878.n14 70.6783
R21754 a_n2804_13878.n21 a_n2804_13878.n13 15.7159
R21755 a_n2804_13878.n23 a_n2804_13878.n21 12.6495
R21756 a_n2804_13878.n21 a_n2804_13878.n20 8.38735
R21757 a_n2804_13878.n22 a_n2804_13878.t15 3.61217
R21758 a_n2804_13878.n22 a_n2804_13878.t24 3.61217
R21759 a_n2804_13878.n24 a_n2804_13878.t28 3.61217
R21760 a_n2804_13878.n24 a_n2804_13878.t14 3.61217
R21761 a_n2804_13878.n26 a_n2804_13878.t18 3.61217
R21762 a_n2804_13878.n26 a_n2804_13878.t19 3.61217
R21763 a_n2804_13878.n1 a_n2804_13878.t8 3.61217
R21764 a_n2804_13878.n1 a_n2804_13878.t20 3.61217
R21765 a_n2804_13878.n0 a_n2804_13878.t25 3.61217
R21766 a_n2804_13878.n0 a_n2804_13878.t31 3.61217
R21767 a_n2804_13878.n18 a_n2804_13878.t6 3.61217
R21768 a_n2804_13878.n18 a_n2804_13878.t7 3.61217
R21769 a_n2804_13878.n14 a_n2804_13878.t4 3.61217
R21770 a_n2804_13878.n14 a_n2804_13878.t5 3.61217
R21771 a_n2804_13878.n12 a_n2804_13878.t21 3.61217
R21772 a_n2804_13878.n12 a_n2804_13878.t9 3.61217
R21773 a_n2804_13878.n10 a_n2804_13878.t26 3.61217
R21774 a_n2804_13878.n10 a_n2804_13878.t11 3.61217
R21775 a_n2804_13878.n8 a_n2804_13878.t10 3.61217
R21776 a_n2804_13878.n8 a_n2804_13878.t13 3.61217
R21777 a_n2804_13878.n6 a_n2804_13878.t23 3.61217
R21778 a_n2804_13878.n6 a_n2804_13878.t16 3.61217
R21779 a_n2804_13878.n4 a_n2804_13878.t27 3.61217
R21780 a_n2804_13878.n4 a_n2804_13878.t17 3.61217
R21781 a_n2804_13878.n3 a_n2804_13878.t12 3.61217
R21782 a_n2804_13878.n3 a_n2804_13878.t22 3.61217
R21783 a_n2804_13878.n29 a_n2804_13878.t29 3.61217
R21784 a_n2804_13878.t30 a_n2804_13878.n29 3.61217
R21785 a_n2804_13878.n16 a_n2804_13878.n15 0.358259
R21786 a_n2804_13878.n19 a_n2804_13878.n17 0.358259
R21787 a_n2804_13878.n20 a_n2804_13878.n19 0.358259
R21788 a_n2804_13878.n28 a_n2804_13878.n2 0.358259
R21789 a_n2804_13878.n28 a_n2804_13878.n27 0.358259
R21790 a_n2804_13878.n27 a_n2804_13878.n25 0.358259
R21791 a_n2804_13878.n25 a_n2804_13878.n23 0.358259
R21792 a_n2804_13878.n7 a_n2804_13878.n5 0.146627
R21793 a_n2804_13878.n9 a_n2804_13878.n7 0.146627
R21794 a_n2804_13878.n11 a_n2804_13878.n9 0.146627
R21795 a_n2804_13878.n13 a_n2804_13878.n11 0.146627
R21796 a_n2804_13878.n17 a_n2804_13878.n16 0.101793
R21797 a_n9628_8799.n225 a_n9628_8799.t137 485.149
R21798 a_n9628_8799.n244 a_n9628_8799.t152 485.149
R21799 a_n9628_8799.n264 a_n9628_8799.t75 485.149
R21800 a_n9628_8799.n164 a_n9628_8799.t89 485.149
R21801 a_n9628_8799.n183 a_n9628_8799.t102 485.149
R21802 a_n9628_8799.n203 a_n9628_8799.t73 485.149
R21803 a_n9628_8799.n56 a_n9628_8799.t46 485.135
R21804 a_n9628_8799.n237 a_n9628_8799.t45 464.166
R21805 a_n9628_8799.n219 a_n9628_8799.t131 464.166
R21806 a_n9628_8799.n236 a_n9628_8799.t67 464.166
R21807 a_n9628_8799.n235 a_n9628_8799.t50 464.166
R21808 a_n9628_8799.n220 a_n9628_8799.t139 464.166
R21809 a_n9628_8799.n234 a_n9628_8799.t94 464.166
R21810 a_n9628_8799.n233 a_n9628_8799.t68 464.166
R21811 a_n9628_8799.n221 a_n9628_8799.t156 464.166
R21812 a_n9628_8799.n232 a_n9628_8799.t111 464.166
R21813 a_n9628_8799.n231 a_n9628_8799.t71 464.166
R21814 a_n9628_8799.n222 a_n9628_8799.t150 464.166
R21815 a_n9628_8799.n230 a_n9628_8799.t113 464.166
R21816 a_n9628_8799.n229 a_n9628_8799.t85 464.166
R21817 a_n9628_8799.n223 a_n9628_8799.t47 464.166
R21818 a_n9628_8799.n228 a_n9628_8799.t134 464.166
R21819 a_n9628_8799.n227 a_n9628_8799.t117 464.166
R21820 a_n9628_8799.n224 a_n9628_8799.t51 464.166
R21821 a_n9628_8799.n226 a_n9628_8799.t141 464.166
R21822 a_n9628_8799.n71 a_n9628_8799.t58 485.135
R21823 a_n9628_8799.n256 a_n9628_8799.t57 464.166
R21824 a_n9628_8799.n238 a_n9628_8799.t148 464.166
R21825 a_n9628_8799.n255 a_n9628_8799.t76 464.166
R21826 a_n9628_8799.n254 a_n9628_8799.t65 464.166
R21827 a_n9628_8799.n239 a_n9628_8799.t151 464.166
R21828 a_n9628_8799.n253 a_n9628_8799.t107 464.166
R21829 a_n9628_8799.n252 a_n9628_8799.t79 464.166
R21830 a_n9628_8799.n240 a_n9628_8799.t49 464.166
R21831 a_n9628_8799.n251 a_n9628_8799.t124 464.166
R21832 a_n9628_8799.n250 a_n9628_8799.t80 464.166
R21833 a_n9628_8799.n241 a_n9628_8799.t41 464.166
R21834 a_n9628_8799.n249 a_n9628_8799.t129 464.166
R21835 a_n9628_8799.n248 a_n9628_8799.t95 464.166
R21836 a_n9628_8799.n242 a_n9628_8799.t59 464.166
R21837 a_n9628_8799.n247 a_n9628_8799.t149 464.166
R21838 a_n9628_8799.n246 a_n9628_8799.t130 464.166
R21839 a_n9628_8799.n243 a_n9628_8799.t66 464.166
R21840 a_n9628_8799.n245 a_n9628_8799.t153 464.166
R21841 a_n9628_8799.n86 a_n9628_8799.t106 485.135
R21842 a_n9628_8799.n276 a_n9628_8799.t128 464.166
R21843 a_n9628_8799.n258 a_n9628_8799.t64 464.166
R21844 a_n9628_8799.n275 a_n9628_8799.t146 464.166
R21845 a_n9628_8799.n274 a_n9628_8799.t83 464.166
R21846 a_n9628_8799.n259 a_n9628_8799.t138 464.166
R21847 a_n9628_8799.n273 a_n9628_8799.t70 464.166
R21848 a_n9628_8799.n272 a_n9628_8799.t118 464.166
R21849 a_n9628_8799.n260 a_n9628_8799.t55 464.166
R21850 a_n9628_8799.n271 a_n9628_8799.t101 464.166
R21851 a_n9628_8799.n270 a_n9628_8799.t78 464.166
R21852 a_n9628_8799.n261 a_n9628_8799.t126 464.166
R21853 a_n9628_8799.n269 a_n9628_8799.t62 464.166
R21854 a_n9628_8799.n268 a_n9628_8799.t110 464.166
R21855 a_n9628_8799.n262 a_n9628_8799.t44 464.166
R21856 a_n9628_8799.n267 a_n9628_8799.t93 464.166
R21857 a_n9628_8799.n266 a_n9628_8799.t158 464.166
R21858 a_n9628_8799.n263 a_n9628_8799.t116 464.166
R21859 a_n9628_8799.n265 a_n9628_8799.t54 464.166
R21860 a_n9628_8799.n165 a_n9628_8799.t91 464.166
R21861 a_n9628_8799.n166 a_n9628_8799.t123 464.166
R21862 a_n9628_8799.n167 a_n9628_8799.t48 464.166
R21863 a_n9628_8799.n168 a_n9628_8799.t87 464.166
R21864 a_n9628_8799.n163 a_n9628_8799.t119 464.166
R21865 a_n9628_8799.n169 a_n9628_8799.t42 464.166
R21866 a_n9628_8799.n170 a_n9628_8799.t74 464.166
R21867 a_n9628_8799.n171 a_n9628_8799.t112 464.166
R21868 a_n9628_8799.n172 a_n9628_8799.t147 464.166
R21869 a_n9628_8799.n162 a_n9628_8799.t72 464.166
R21870 a_n9628_8799.n173 a_n9628_8799.t108 464.166
R21871 a_n9628_8799.n161 a_n9628_8799.t143 464.166
R21872 a_n9628_8799.n174 a_n9628_8799.t144 464.166
R21873 a_n9628_8799.n175 a_n9628_8799.t90 464.166
R21874 a_n9628_8799.n176 a_n9628_8799.t122 464.166
R21875 a_n9628_8799.n177 a_n9628_8799.t142 464.166
R21876 a_n9628_8799.n160 a_n9628_8799.t86 464.166
R21877 a_n9628_8799.n178 a_n9628_8799.t88 464.166
R21878 a_n9628_8799.n184 a_n9628_8799.t104 464.166
R21879 a_n9628_8799.n185 a_n9628_8799.t140 464.166
R21880 a_n9628_8799.n186 a_n9628_8799.t60 464.166
R21881 a_n9628_8799.n187 a_n9628_8799.t98 464.166
R21882 a_n9628_8799.n182 a_n9628_8799.t132 464.166
R21883 a_n9628_8799.n188 a_n9628_8799.t56 464.166
R21884 a_n9628_8799.n189 a_n9628_8799.t84 464.166
R21885 a_n9628_8799.n190 a_n9628_8799.t125 464.166
R21886 a_n9628_8799.n191 a_n9628_8799.t159 464.166
R21887 a_n9628_8799.n181 a_n9628_8799.t81 464.166
R21888 a_n9628_8799.n192 a_n9628_8799.t121 464.166
R21889 a_n9628_8799.n180 a_n9628_8799.t155 464.166
R21890 a_n9628_8799.n193 a_n9628_8799.t157 464.166
R21891 a_n9628_8799.n194 a_n9628_8799.t103 464.166
R21892 a_n9628_8799.n195 a_n9628_8799.t136 464.166
R21893 a_n9628_8799.n196 a_n9628_8799.t154 464.166
R21894 a_n9628_8799.n179 a_n9628_8799.t97 464.166
R21895 a_n9628_8799.n197 a_n9628_8799.t99 464.166
R21896 a_n9628_8799.n204 a_n9628_8799.t52 464.166
R21897 a_n9628_8799.n205 a_n9628_8799.t114 464.166
R21898 a_n9628_8799.n206 a_n9628_8799.t69 464.166
R21899 a_n9628_8799.n207 a_n9628_8799.t92 464.166
R21900 a_n9628_8799.n202 a_n9628_8799.t43 464.166
R21901 a_n9628_8799.n208 a_n9628_8799.t109 464.166
R21902 a_n9628_8799.n209 a_n9628_8799.t61 464.166
R21903 a_n9628_8799.n210 a_n9628_8799.t127 464.166
R21904 a_n9628_8799.n211 a_n9628_8799.t77 464.166
R21905 a_n9628_8799.n201 a_n9628_8799.t100 464.166
R21906 a_n9628_8799.n212 a_n9628_8799.t53 464.166
R21907 a_n9628_8799.n200 a_n9628_8799.t115 464.166
R21908 a_n9628_8799.n213 a_n9628_8799.t96 464.166
R21909 a_n9628_8799.n214 a_n9628_8799.t135 464.166
R21910 a_n9628_8799.n215 a_n9628_8799.t82 464.166
R21911 a_n9628_8799.n216 a_n9628_8799.t145 464.166
R21912 a_n9628_8799.n199 a_n9628_8799.t63 464.166
R21913 a_n9628_8799.n217 a_n9628_8799.t40 464.166
R21914 a_n9628_8799.n44 a_n9628_8799.n70 71.7212
R21915 a_n9628_8799.n70 a_n9628_8799.n224 17.8606
R21916 a_n9628_8799.n69 a_n9628_8799.n44 76.9909
R21917 a_n9628_8799.n227 a_n9628_8799.n69 7.32118
R21918 a_n9628_8799.n68 a_n9628_8799.n43 78.3454
R21919 a_n9628_8799.n43 a_n9628_8799.n67 72.8951
R21920 a_n9628_8799.n66 a_n9628_8799.n45 70.1674
R21921 a_n9628_8799.n230 a_n9628_8799.n66 20.9683
R21922 a_n9628_8799.n45 a_n9628_8799.n65 72.3034
R21923 a_n9628_8799.n65 a_n9628_8799.n222 16.6962
R21924 a_n9628_8799.n64 a_n9628_8799.n46 77.6622
R21925 a_n9628_8799.n231 a_n9628_8799.n64 5.97853
R21926 a_n9628_8799.n63 a_n9628_8799.n46 77.6622
R21927 a_n9628_8799.n47 a_n9628_8799.n62 72.3034
R21928 a_n9628_8799.n61 a_n9628_8799.n47 70.1674
R21929 a_n9628_8799.n234 a_n9628_8799.n61 20.9683
R21930 a_n9628_8799.n49 a_n9628_8799.n60 72.8951
R21931 a_n9628_8799.n60 a_n9628_8799.n220 15.5127
R21932 a_n9628_8799.n59 a_n9628_8799.n49 78.3454
R21933 a_n9628_8799.n235 a_n9628_8799.n59 4.61226
R21934 a_n9628_8799.n58 a_n9628_8799.n48 76.9909
R21935 a_n9628_8799.n48 a_n9628_8799.n57 71.7212
R21936 a_n9628_8799.n237 a_n9628_8799.n56 20.9683
R21937 a_n9628_8799.n50 a_n9628_8799.n56 70.1674
R21938 a_n9628_8799.n36 a_n9628_8799.n85 71.7212
R21939 a_n9628_8799.n85 a_n9628_8799.n243 17.8606
R21940 a_n9628_8799.n84 a_n9628_8799.n36 76.9909
R21941 a_n9628_8799.n246 a_n9628_8799.n84 7.32118
R21942 a_n9628_8799.n83 a_n9628_8799.n35 78.3454
R21943 a_n9628_8799.n35 a_n9628_8799.n82 72.8951
R21944 a_n9628_8799.n81 a_n9628_8799.n37 70.1674
R21945 a_n9628_8799.n249 a_n9628_8799.n81 20.9683
R21946 a_n9628_8799.n37 a_n9628_8799.n80 72.3034
R21947 a_n9628_8799.n80 a_n9628_8799.n241 16.6962
R21948 a_n9628_8799.n79 a_n9628_8799.n38 77.6622
R21949 a_n9628_8799.n250 a_n9628_8799.n79 5.97853
R21950 a_n9628_8799.n78 a_n9628_8799.n38 77.6622
R21951 a_n9628_8799.n39 a_n9628_8799.n77 72.3034
R21952 a_n9628_8799.n76 a_n9628_8799.n39 70.1674
R21953 a_n9628_8799.n253 a_n9628_8799.n76 20.9683
R21954 a_n9628_8799.n41 a_n9628_8799.n75 72.8951
R21955 a_n9628_8799.n75 a_n9628_8799.n239 15.5127
R21956 a_n9628_8799.n74 a_n9628_8799.n41 78.3454
R21957 a_n9628_8799.n254 a_n9628_8799.n74 4.61226
R21958 a_n9628_8799.n73 a_n9628_8799.n40 76.9909
R21959 a_n9628_8799.n40 a_n9628_8799.n72 71.7212
R21960 a_n9628_8799.n256 a_n9628_8799.n71 20.9683
R21961 a_n9628_8799.n42 a_n9628_8799.n71 70.1674
R21962 a_n9628_8799.n28 a_n9628_8799.n100 71.7212
R21963 a_n9628_8799.n100 a_n9628_8799.n263 17.8606
R21964 a_n9628_8799.n99 a_n9628_8799.n28 76.9909
R21965 a_n9628_8799.n266 a_n9628_8799.n99 7.32118
R21966 a_n9628_8799.n98 a_n9628_8799.n27 78.3454
R21967 a_n9628_8799.n27 a_n9628_8799.n97 72.8951
R21968 a_n9628_8799.n96 a_n9628_8799.n29 70.1674
R21969 a_n9628_8799.n269 a_n9628_8799.n96 20.9683
R21970 a_n9628_8799.n29 a_n9628_8799.n95 72.3034
R21971 a_n9628_8799.n95 a_n9628_8799.n261 16.6962
R21972 a_n9628_8799.n94 a_n9628_8799.n30 77.6622
R21973 a_n9628_8799.n270 a_n9628_8799.n94 5.97853
R21974 a_n9628_8799.n93 a_n9628_8799.n30 77.6622
R21975 a_n9628_8799.n31 a_n9628_8799.n92 72.3034
R21976 a_n9628_8799.n91 a_n9628_8799.n31 70.1674
R21977 a_n9628_8799.n273 a_n9628_8799.n91 20.9683
R21978 a_n9628_8799.n33 a_n9628_8799.n90 72.8951
R21979 a_n9628_8799.n90 a_n9628_8799.n259 15.5127
R21980 a_n9628_8799.n89 a_n9628_8799.n33 78.3454
R21981 a_n9628_8799.n274 a_n9628_8799.n89 4.61226
R21982 a_n9628_8799.n88 a_n9628_8799.n32 76.9909
R21983 a_n9628_8799.n32 a_n9628_8799.n87 71.7212
R21984 a_n9628_8799.n276 a_n9628_8799.n86 20.9683
R21985 a_n9628_8799.n34 a_n9628_8799.n86 70.1674
R21986 a_n9628_8799.n20 a_n9628_8799.n115 70.1674
R21987 a_n9628_8799.n178 a_n9628_8799.n115 20.9683
R21988 a_n9628_8799.n114 a_n9628_8799.n20 71.7212
R21989 a_n9628_8799.n114 a_n9628_8799.n160 17.8606
R21990 a_n9628_8799.n19 a_n9628_8799.n113 76.9909
R21991 a_n9628_8799.n177 a_n9628_8799.n113 7.32118
R21992 a_n9628_8799.n112 a_n9628_8799.n19 78.3454
R21993 a_n9628_8799.n21 a_n9628_8799.n111 72.8951
R21994 a_n9628_8799.n110 a_n9628_8799.n21 70.1674
R21995 a_n9628_8799.n110 a_n9628_8799.n161 20.9683
R21996 a_n9628_8799.n22 a_n9628_8799.n109 72.3034
R21997 a_n9628_8799.n173 a_n9628_8799.n109 16.6962
R21998 a_n9628_8799.n108 a_n9628_8799.n22 77.6622
R21999 a_n9628_8799.n108 a_n9628_8799.n162 5.97853
R22000 a_n9628_8799.n23 a_n9628_8799.n107 77.6622
R22001 a_n9628_8799.n106 a_n9628_8799.n23 72.3034
R22002 a_n9628_8799.n24 a_n9628_8799.n105 70.1674
R22003 a_n9628_8799.n169 a_n9628_8799.n105 20.9683
R22004 a_n9628_8799.n104 a_n9628_8799.n24 72.8951
R22005 a_n9628_8799.n104 a_n9628_8799.n163 15.5127
R22006 a_n9628_8799.n25 a_n9628_8799.n103 78.3454
R22007 a_n9628_8799.n168 a_n9628_8799.n103 4.61226
R22008 a_n9628_8799.n102 a_n9628_8799.n25 76.9909
R22009 a_n9628_8799.n101 a_n9628_8799.n166 17.8606
R22010 a_n9628_8799.n101 a_n9628_8799.n26 71.7212
R22011 a_n9628_8799.n12 a_n9628_8799.n130 70.1674
R22012 a_n9628_8799.n197 a_n9628_8799.n130 20.9683
R22013 a_n9628_8799.n129 a_n9628_8799.n12 71.7212
R22014 a_n9628_8799.n129 a_n9628_8799.n179 17.8606
R22015 a_n9628_8799.n11 a_n9628_8799.n128 76.9909
R22016 a_n9628_8799.n196 a_n9628_8799.n128 7.32118
R22017 a_n9628_8799.n127 a_n9628_8799.n11 78.3454
R22018 a_n9628_8799.n13 a_n9628_8799.n126 72.8951
R22019 a_n9628_8799.n125 a_n9628_8799.n13 70.1674
R22020 a_n9628_8799.n125 a_n9628_8799.n180 20.9683
R22021 a_n9628_8799.n14 a_n9628_8799.n124 72.3034
R22022 a_n9628_8799.n192 a_n9628_8799.n124 16.6962
R22023 a_n9628_8799.n123 a_n9628_8799.n14 77.6622
R22024 a_n9628_8799.n123 a_n9628_8799.n181 5.97853
R22025 a_n9628_8799.n15 a_n9628_8799.n122 77.6622
R22026 a_n9628_8799.n121 a_n9628_8799.n15 72.3034
R22027 a_n9628_8799.n16 a_n9628_8799.n120 70.1674
R22028 a_n9628_8799.n188 a_n9628_8799.n120 20.9683
R22029 a_n9628_8799.n119 a_n9628_8799.n16 72.8951
R22030 a_n9628_8799.n119 a_n9628_8799.n182 15.5127
R22031 a_n9628_8799.n17 a_n9628_8799.n118 78.3454
R22032 a_n9628_8799.n187 a_n9628_8799.n118 4.61226
R22033 a_n9628_8799.n117 a_n9628_8799.n17 76.9909
R22034 a_n9628_8799.n116 a_n9628_8799.n185 17.8606
R22035 a_n9628_8799.n116 a_n9628_8799.n18 71.7212
R22036 a_n9628_8799.n4 a_n9628_8799.n145 70.1674
R22037 a_n9628_8799.n217 a_n9628_8799.n145 20.9683
R22038 a_n9628_8799.n144 a_n9628_8799.n4 71.7212
R22039 a_n9628_8799.n144 a_n9628_8799.n199 17.8606
R22040 a_n9628_8799.n3 a_n9628_8799.n143 76.9909
R22041 a_n9628_8799.n216 a_n9628_8799.n143 7.32118
R22042 a_n9628_8799.n142 a_n9628_8799.n3 78.3454
R22043 a_n9628_8799.n5 a_n9628_8799.n141 72.8951
R22044 a_n9628_8799.n140 a_n9628_8799.n5 70.1674
R22045 a_n9628_8799.n140 a_n9628_8799.n200 20.9683
R22046 a_n9628_8799.n6 a_n9628_8799.n139 72.3034
R22047 a_n9628_8799.n212 a_n9628_8799.n139 16.6962
R22048 a_n9628_8799.n138 a_n9628_8799.n6 77.6622
R22049 a_n9628_8799.n138 a_n9628_8799.n201 5.97853
R22050 a_n9628_8799.n7 a_n9628_8799.n137 77.6622
R22051 a_n9628_8799.n136 a_n9628_8799.n7 72.3034
R22052 a_n9628_8799.n8 a_n9628_8799.n135 70.1674
R22053 a_n9628_8799.n208 a_n9628_8799.n135 20.9683
R22054 a_n9628_8799.n134 a_n9628_8799.n8 72.8951
R22055 a_n9628_8799.n134 a_n9628_8799.n202 15.5127
R22056 a_n9628_8799.n9 a_n9628_8799.n133 78.3454
R22057 a_n9628_8799.n207 a_n9628_8799.n133 4.61226
R22058 a_n9628_8799.n132 a_n9628_8799.n9 76.9909
R22059 a_n9628_8799.n131 a_n9628_8799.n205 17.8606
R22060 a_n9628_8799.n131 a_n9628_8799.n10 71.7212
R22061 a_n9628_8799.n51 a_n9628_8799.n146 98.9633
R22062 a_n9628_8799.n54 a_n9628_8799.n281 98.9631
R22063 a_n9628_8799.n54 a_n9628_8799.n282 98.6055
R22064 a_n9628_8799.n54 a_n9628_8799.n283 98.6055
R22065 a_n9628_8799.n55 a_n9628_8799.n284 98.6055
R22066 a_n9628_8799.n55 a_n9628_8799.n285 98.6055
R22067 a_n9628_8799.n53 a_n9628_8799.n151 98.6055
R22068 a_n9628_8799.n53 a_n9628_8799.n150 98.6055
R22069 a_n9628_8799.n52 a_n9628_8799.n149 98.6055
R22070 a_n9628_8799.n52 a_n9628_8799.n148 98.6055
R22071 a_n9628_8799.n51 a_n9628_8799.n147 98.6055
R22072 a_n9628_8799.n287 a_n9628_8799.n286 98.6054
R22073 a_n9628_8799.n1 a_n9628_8799.n152 81.4626
R22074 a_n9628_8799.n2 a_n9628_8799.n156 81.4626
R22075 a_n9628_8799.n2 a_n9628_8799.n154 81.4626
R22076 a_n9628_8799.n0 a_n9628_8799.n158 80.9324
R22077 a_n9628_8799.n1 a_n9628_8799.n159 80.9324
R22078 a_n9628_8799.n1 a_n9628_8799.n153 80.9324
R22079 a_n9628_8799.n2 a_n9628_8799.n157 80.9324
R22080 a_n9628_8799.n2 a_n9628_8799.n155 80.9324
R22081 a_n9628_8799.n44 a_n9628_8799.n225 70.4033
R22082 a_n9628_8799.n36 a_n9628_8799.n244 70.4033
R22083 a_n9628_8799.n28 a_n9628_8799.n264 70.4033
R22084 a_n9628_8799.n164 a_n9628_8799.n26 70.4033
R22085 a_n9628_8799.n183 a_n9628_8799.n18 70.4033
R22086 a_n9628_8799.n203 a_n9628_8799.n10 70.4033
R22087 a_n9628_8799.n236 a_n9628_8799.n235 48.2005
R22088 a_n9628_8799.n61 a_n9628_8799.n233 20.9683
R22089 a_n9628_8799.n232 a_n9628_8799.n231 48.2005
R22090 a_n9628_8799.n66 a_n9628_8799.n229 20.9683
R22091 a_n9628_8799.n228 a_n9628_8799.n227 48.2005
R22092 a_n9628_8799.n255 a_n9628_8799.n254 48.2005
R22093 a_n9628_8799.n76 a_n9628_8799.n252 20.9683
R22094 a_n9628_8799.n251 a_n9628_8799.n250 48.2005
R22095 a_n9628_8799.n81 a_n9628_8799.n248 20.9683
R22096 a_n9628_8799.n247 a_n9628_8799.n246 48.2005
R22097 a_n9628_8799.n275 a_n9628_8799.n274 48.2005
R22098 a_n9628_8799.n91 a_n9628_8799.n272 20.9683
R22099 a_n9628_8799.n271 a_n9628_8799.n270 48.2005
R22100 a_n9628_8799.n96 a_n9628_8799.n268 20.9683
R22101 a_n9628_8799.n267 a_n9628_8799.n266 48.2005
R22102 a_n9628_8799.n168 a_n9628_8799.n167 48.2005
R22103 a_n9628_8799.n170 a_n9628_8799.n105 20.9683
R22104 a_n9628_8799.n172 a_n9628_8799.n162 48.2005
R22105 a_n9628_8799.n174 a_n9628_8799.n110 20.9683
R22106 a_n9628_8799.n177 a_n9628_8799.n176 48.2005
R22107 a_n9628_8799.t120 a_n9628_8799.n115 485.135
R22108 a_n9628_8799.n187 a_n9628_8799.n186 48.2005
R22109 a_n9628_8799.n189 a_n9628_8799.n120 20.9683
R22110 a_n9628_8799.n191 a_n9628_8799.n181 48.2005
R22111 a_n9628_8799.n193 a_n9628_8799.n125 20.9683
R22112 a_n9628_8799.n196 a_n9628_8799.n195 48.2005
R22113 a_n9628_8799.t133 a_n9628_8799.n130 485.135
R22114 a_n9628_8799.n207 a_n9628_8799.n206 48.2005
R22115 a_n9628_8799.n209 a_n9628_8799.n135 20.9683
R22116 a_n9628_8799.n211 a_n9628_8799.n201 48.2005
R22117 a_n9628_8799.n213 a_n9628_8799.n140 20.9683
R22118 a_n9628_8799.n216 a_n9628_8799.n215 48.2005
R22119 a_n9628_8799.t105 a_n9628_8799.n145 485.135
R22120 a_n9628_8799.n57 a_n9628_8799.n219 17.8606
R22121 a_n9628_8799.n226 a_n9628_8799.n70 25.894
R22122 a_n9628_8799.n72 a_n9628_8799.n238 17.8606
R22123 a_n9628_8799.n245 a_n9628_8799.n85 25.894
R22124 a_n9628_8799.n87 a_n9628_8799.n258 17.8606
R22125 a_n9628_8799.n265 a_n9628_8799.n100 25.894
R22126 a_n9628_8799.n178 a_n9628_8799.n114 25.894
R22127 a_n9628_8799.n197 a_n9628_8799.n129 25.894
R22128 a_n9628_8799.n217 a_n9628_8799.n144 25.894
R22129 a_n9628_8799.n68 a_n9628_8799.n223 43.3183
R22130 a_n9628_8799.n83 a_n9628_8799.n242 43.3183
R22131 a_n9628_8799.n98 a_n9628_8799.n262 43.3183
R22132 a_n9628_8799.n175 a_n9628_8799.n112 43.3183
R22133 a_n9628_8799.n194 a_n9628_8799.n127 43.3183
R22134 a_n9628_8799.n214 a_n9628_8799.n142 43.3183
R22135 a_n9628_8799.n62 a_n9628_8799.n221 16.6962
R22136 a_n9628_8799.n230 a_n9628_8799.n65 27.6507
R22137 a_n9628_8799.n77 a_n9628_8799.n240 16.6962
R22138 a_n9628_8799.n249 a_n9628_8799.n80 27.6507
R22139 a_n9628_8799.n92 a_n9628_8799.n260 16.6962
R22140 a_n9628_8799.n269 a_n9628_8799.n95 27.6507
R22141 a_n9628_8799.n171 a_n9628_8799.n106 16.6962
R22142 a_n9628_8799.n161 a_n9628_8799.n109 27.6507
R22143 a_n9628_8799.n190 a_n9628_8799.n121 16.6962
R22144 a_n9628_8799.n180 a_n9628_8799.n124 27.6507
R22145 a_n9628_8799.n210 a_n9628_8799.n136 16.6962
R22146 a_n9628_8799.n200 a_n9628_8799.n139 27.6507
R22147 a_n9628_8799.n63 a_n9628_8799.n221 41.7634
R22148 a_n9628_8799.n78 a_n9628_8799.n240 41.7634
R22149 a_n9628_8799.n93 a_n9628_8799.n260 41.7634
R22150 a_n9628_8799.n107 a_n9628_8799.n171 41.7634
R22151 a_n9628_8799.n122 a_n9628_8799.n190 41.7634
R22152 a_n9628_8799.n137 a_n9628_8799.n210 41.7634
R22153 a_n9628_8799.n234 a_n9628_8799.n60 29.3885
R22154 a_n9628_8799.n67 a_n9628_8799.n223 15.5127
R22155 a_n9628_8799.n253 a_n9628_8799.n75 29.3885
R22156 a_n9628_8799.n82 a_n9628_8799.n242 15.5127
R22157 a_n9628_8799.n273 a_n9628_8799.n90 29.3885
R22158 a_n9628_8799.n97 a_n9628_8799.n262 15.5127
R22159 a_n9628_8799.n169 a_n9628_8799.n104 29.3885
R22160 a_n9628_8799.n175 a_n9628_8799.n111 15.5127
R22161 a_n9628_8799.n188 a_n9628_8799.n119 29.3885
R22162 a_n9628_8799.n194 a_n9628_8799.n126 15.5127
R22163 a_n9628_8799.n208 a_n9628_8799.n134 29.3885
R22164 a_n9628_8799.n214 a_n9628_8799.n141 15.5127
R22165 a_n9628_8799.n286 a_n9628_8799.n280 33.8838
R22166 a_n9628_8799.n58 a_n9628_8799.n219 40.1848
R22167 a_n9628_8799.n73 a_n9628_8799.n238 40.1848
R22168 a_n9628_8799.n88 a_n9628_8799.n258 40.1848
R22169 a_n9628_8799.n166 a_n9628_8799.n102 40.1848
R22170 a_n9628_8799.n185 a_n9628_8799.n117 40.1848
R22171 a_n9628_8799.n205 a_n9628_8799.n132 40.1848
R22172 a_n9628_8799.n280 a_n9628_8799.n53 21.0055
R22173 a_n9628_8799.n226 a_n9628_8799.n225 20.9576
R22174 a_n9628_8799.n245 a_n9628_8799.n244 20.9576
R22175 a_n9628_8799.n265 a_n9628_8799.n264 20.9576
R22176 a_n9628_8799.n165 a_n9628_8799.n164 20.9576
R22177 a_n9628_8799.n184 a_n9628_8799.n183 20.9576
R22178 a_n9628_8799.n204 a_n9628_8799.n203 20.9576
R22179 a_n9628_8799.n58 a_n9628_8799.n236 7.32118
R22180 a_n9628_8799.n69 a_n9628_8799.n224 40.1848
R22181 a_n9628_8799.n73 a_n9628_8799.n255 7.32118
R22182 a_n9628_8799.n84 a_n9628_8799.n243 40.1848
R22183 a_n9628_8799.n88 a_n9628_8799.n275 7.32118
R22184 a_n9628_8799.n99 a_n9628_8799.n263 40.1848
R22185 a_n9628_8799.n167 a_n9628_8799.n102 7.32118
R22186 a_n9628_8799.n160 a_n9628_8799.n113 40.1848
R22187 a_n9628_8799.n186 a_n9628_8799.n117 7.32118
R22188 a_n9628_8799.n179 a_n9628_8799.n128 40.1848
R22189 a_n9628_8799.n206 a_n9628_8799.n132 7.32118
R22190 a_n9628_8799.n199 a_n9628_8799.n143 40.1848
R22191 a_n9628_8799.n229 a_n9628_8799.n67 29.3885
R22192 a_n9628_8799.n248 a_n9628_8799.n82 29.3885
R22193 a_n9628_8799.n268 a_n9628_8799.n97 29.3885
R22194 a_n9628_8799.n111 a_n9628_8799.n174 29.3885
R22195 a_n9628_8799.n126 a_n9628_8799.n193 29.3885
R22196 a_n9628_8799.n141 a_n9628_8799.n213 29.3885
R22197 a_n9628_8799.n63 a_n9628_8799.n232 5.97853
R22198 a_n9628_8799.n64 a_n9628_8799.n222 41.7634
R22199 a_n9628_8799.n78 a_n9628_8799.n251 5.97853
R22200 a_n9628_8799.n79 a_n9628_8799.n241 41.7634
R22201 a_n9628_8799.n93 a_n9628_8799.n271 5.97853
R22202 a_n9628_8799.n94 a_n9628_8799.n261 41.7634
R22203 a_n9628_8799.n172 a_n9628_8799.n107 5.97853
R22204 a_n9628_8799.n173 a_n9628_8799.n108 41.7634
R22205 a_n9628_8799.n191 a_n9628_8799.n122 5.97853
R22206 a_n9628_8799.n192 a_n9628_8799.n123 41.7634
R22207 a_n9628_8799.n211 a_n9628_8799.n137 5.97853
R22208 a_n9628_8799.n212 a_n9628_8799.n138 41.7634
R22209 a_n9628_8799.n279 a_n9628_8799.n1 12.3339
R22210 a_n9628_8799.n280 a_n9628_8799.n279 11.4887
R22211 a_n9628_8799.n233 a_n9628_8799.n62 27.6507
R22212 a_n9628_8799.n252 a_n9628_8799.n77 27.6507
R22213 a_n9628_8799.n272 a_n9628_8799.n92 27.6507
R22214 a_n9628_8799.n170 a_n9628_8799.n106 27.6507
R22215 a_n9628_8799.n189 a_n9628_8799.n121 27.6507
R22216 a_n9628_8799.n209 a_n9628_8799.n136 27.6507
R22217 a_n9628_8799.n59 a_n9628_8799.n220 43.3183
R22218 a_n9628_8799.n68 a_n9628_8799.n228 4.61226
R22219 a_n9628_8799.n74 a_n9628_8799.n239 43.3183
R22220 a_n9628_8799.n83 a_n9628_8799.n247 4.61226
R22221 a_n9628_8799.n89 a_n9628_8799.n259 43.3183
R22222 a_n9628_8799.n98 a_n9628_8799.n267 4.61226
R22223 a_n9628_8799.n163 a_n9628_8799.n103 43.3183
R22224 a_n9628_8799.n176 a_n9628_8799.n112 4.61226
R22225 a_n9628_8799.n182 a_n9628_8799.n118 43.3183
R22226 a_n9628_8799.n195 a_n9628_8799.n127 4.61226
R22227 a_n9628_8799.n202 a_n9628_8799.n133 43.3183
R22228 a_n9628_8799.n0 a_n9628_8799.n2 33.2634
R22229 a_n9628_8799.n215 a_n9628_8799.n142 4.61226
R22230 a_n9628_8799.n257 a_n9628_8799.n50 9.04406
R22231 a_n9628_8799.n198 a_n9628_8799.n20 9.04406
R22232 a_n9628_8799.n237 a_n9628_8799.n57 25.894
R22233 a_n9628_8799.n256 a_n9628_8799.n72 25.894
R22234 a_n9628_8799.n276 a_n9628_8799.n87 25.894
R22235 a_n9628_8799.n101 a_n9628_8799.n165 25.894
R22236 a_n9628_8799.n116 a_n9628_8799.n184 25.894
R22237 a_n9628_8799.n131 a_n9628_8799.n204 25.894
R22238 a_n9628_8799.n278 a_n9628_8799.n218 7.17472
R22239 a_n9628_8799.n278 a_n9628_8799.n277 6.83225
R22240 a_n9628_8799.n257 a_n9628_8799.n42 4.93611
R22241 a_n9628_8799.n277 a_n9628_8799.n34 4.93611
R22242 a_n9628_8799.n198 a_n9628_8799.n12 4.93611
R22243 a_n9628_8799.n218 a_n9628_8799.n4 4.93611
R22244 a_n9628_8799.n277 a_n9628_8799.n257 4.10845
R22245 a_n9628_8799.n218 a_n9628_8799.n198 4.10845
R22246 a_n9628_8799.n281 a_n9628_8799.t34 3.61217
R22247 a_n9628_8799.n281 a_n9628_8799.t27 3.61217
R22248 a_n9628_8799.n282 a_n9628_8799.t26 3.61217
R22249 a_n9628_8799.n282 a_n9628_8799.t39 3.61217
R22250 a_n9628_8799.n283 a_n9628_8799.t31 3.61217
R22251 a_n9628_8799.n283 a_n9628_8799.t30 3.61217
R22252 a_n9628_8799.n284 a_n9628_8799.t28 3.61217
R22253 a_n9628_8799.n284 a_n9628_8799.t29 3.61217
R22254 a_n9628_8799.n285 a_n9628_8799.t20 3.61217
R22255 a_n9628_8799.n285 a_n9628_8799.t35 3.61217
R22256 a_n9628_8799.n151 a_n9628_8799.t37 3.61217
R22257 a_n9628_8799.n151 a_n9628_8799.t22 3.61217
R22258 a_n9628_8799.n150 a_n9628_8799.t19 3.61217
R22259 a_n9628_8799.n150 a_n9628_8799.t38 3.61217
R22260 a_n9628_8799.n149 a_n9628_8799.t25 3.61217
R22261 a_n9628_8799.n149 a_n9628_8799.t33 3.61217
R22262 a_n9628_8799.n148 a_n9628_8799.t21 3.61217
R22263 a_n9628_8799.n148 a_n9628_8799.t24 3.61217
R22264 a_n9628_8799.n147 a_n9628_8799.t18 3.61217
R22265 a_n9628_8799.n147 a_n9628_8799.t17 3.61217
R22266 a_n9628_8799.n146 a_n9628_8799.t36 3.61217
R22267 a_n9628_8799.n146 a_n9628_8799.t32 3.61217
R22268 a_n9628_8799.n287 a_n9628_8799.t23 3.61217
R22269 a_n9628_8799.t16 a_n9628_8799.n287 3.61217
R22270 a_n9628_8799.n279 a_n9628_8799.n278 3.4105
R22271 a_n9628_8799.n158 a_n9628_8799.t3 2.82907
R22272 a_n9628_8799.n158 a_n9628_8799.t2 2.82907
R22273 a_n9628_8799.n159 a_n9628_8799.t0 2.82907
R22274 a_n9628_8799.n159 a_n9628_8799.t13 2.82907
R22275 a_n9628_8799.n153 a_n9628_8799.t4 2.82907
R22276 a_n9628_8799.n153 a_n9628_8799.t12 2.82907
R22277 a_n9628_8799.n152 a_n9628_8799.t6 2.82907
R22278 a_n9628_8799.n152 a_n9628_8799.t1 2.82907
R22279 a_n9628_8799.n156 a_n9628_8799.t14 2.82907
R22280 a_n9628_8799.n156 a_n9628_8799.t7 2.82907
R22281 a_n9628_8799.n157 a_n9628_8799.t5 2.82907
R22282 a_n9628_8799.n157 a_n9628_8799.t9 2.82907
R22283 a_n9628_8799.n155 a_n9628_8799.t10 2.82907
R22284 a_n9628_8799.n155 a_n9628_8799.t8 2.82907
R22285 a_n9628_8799.n154 a_n9628_8799.t11 2.82907
R22286 a_n9628_8799.n154 a_n9628_8799.t15 2.82907
R22287 a_n9628_8799.n44 a_n9628_8799.n43 1.13686
R22288 a_n9628_8799.n36 a_n9628_8799.n35 1.13686
R22289 a_n9628_8799.n28 a_n9628_8799.n27 1.13686
R22290 a_n9628_8799.n20 a_n9628_8799.n19 1.13686
R22291 a_n9628_8799.n12 a_n9628_8799.n11 1.13686
R22292 a_n9628_8799.n4 a_n9628_8799.n3 1.13686
R22293 a_n9628_8799.n1 a_n9628_8799.n0 1.06084
R22294 a_n9628_8799.n49 a_n9628_8799.n48 0.758076
R22295 a_n9628_8799.n49 a_n9628_8799.n47 0.758076
R22296 a_n9628_8799.n47 a_n9628_8799.n46 0.758076
R22297 a_n9628_8799.n46 a_n9628_8799.n45 0.758076
R22298 a_n9628_8799.n43 a_n9628_8799.n45 0.758076
R22299 a_n9628_8799.n41 a_n9628_8799.n40 0.758076
R22300 a_n9628_8799.n41 a_n9628_8799.n39 0.758076
R22301 a_n9628_8799.n39 a_n9628_8799.n38 0.758076
R22302 a_n9628_8799.n38 a_n9628_8799.n37 0.758076
R22303 a_n9628_8799.n35 a_n9628_8799.n37 0.758076
R22304 a_n9628_8799.n33 a_n9628_8799.n32 0.758076
R22305 a_n9628_8799.n33 a_n9628_8799.n31 0.758076
R22306 a_n9628_8799.n31 a_n9628_8799.n30 0.758076
R22307 a_n9628_8799.n30 a_n9628_8799.n29 0.758076
R22308 a_n9628_8799.n27 a_n9628_8799.n29 0.758076
R22309 a_n9628_8799.n24 a_n9628_8799.n25 0.758076
R22310 a_n9628_8799.n23 a_n9628_8799.n24 0.758076
R22311 a_n9628_8799.n22 a_n9628_8799.n23 0.758076
R22312 a_n9628_8799.n21 a_n9628_8799.n22 0.758076
R22313 a_n9628_8799.n19 a_n9628_8799.n21 0.758076
R22314 a_n9628_8799.n16 a_n9628_8799.n17 0.758076
R22315 a_n9628_8799.n15 a_n9628_8799.n16 0.758076
R22316 a_n9628_8799.n14 a_n9628_8799.n15 0.758076
R22317 a_n9628_8799.n13 a_n9628_8799.n14 0.758076
R22318 a_n9628_8799.n11 a_n9628_8799.n13 0.758076
R22319 a_n9628_8799.n8 a_n9628_8799.n9 0.758076
R22320 a_n9628_8799.n7 a_n9628_8799.n8 0.758076
R22321 a_n9628_8799.n6 a_n9628_8799.n7 0.758076
R22322 a_n9628_8799.n5 a_n9628_8799.n6 0.758076
R22323 a_n9628_8799.n3 a_n9628_8799.n5 0.758076
R22324 a_n9628_8799.n55 a_n9628_8799.n54 0.716017
R22325 a_n9628_8799.n286 a_n9628_8799.n55 0.716017
R22326 a_n9628_8799.n53 a_n9628_8799.n52 0.716017
R22327 a_n9628_8799.n52 a_n9628_8799.n51 0.716017
R22328 a_n9628_8799.n9 a_n9628_8799.n10 0.568682
R22329 a_n9628_8799.n17 a_n9628_8799.n18 0.568682
R22330 a_n9628_8799.n25 a_n9628_8799.n26 0.568682
R22331 a_n9628_8799.n32 a_n9628_8799.n34 0.568682
R22332 a_n9628_8799.n40 a_n9628_8799.n42 0.568682
R22333 a_n9628_8799.n48 a_n9628_8799.n50 0.568682
R22334 output.n41 output.n15 289.615
R22335 output.n72 output.n46 289.615
R22336 output.n104 output.n78 289.615
R22337 output.n136 output.n110 289.615
R22338 output.n77 output.n45 197.26
R22339 output.n77 output.n76 196.298
R22340 output.n109 output.n108 196.298
R22341 output.n141 output.n140 196.298
R22342 output.n42 output.n41 185
R22343 output.n40 output.n39 185
R22344 output.n19 output.n18 185
R22345 output.n34 output.n33 185
R22346 output.n32 output.n31 185
R22347 output.n23 output.n22 185
R22348 output.n26 output.n25 185
R22349 output.n73 output.n72 185
R22350 output.n71 output.n70 185
R22351 output.n50 output.n49 185
R22352 output.n65 output.n64 185
R22353 output.n63 output.n62 185
R22354 output.n54 output.n53 185
R22355 output.n57 output.n56 185
R22356 output.n105 output.n104 185
R22357 output.n103 output.n102 185
R22358 output.n82 output.n81 185
R22359 output.n97 output.n96 185
R22360 output.n95 output.n94 185
R22361 output.n86 output.n85 185
R22362 output.n89 output.n88 185
R22363 output.n137 output.n136 185
R22364 output.n135 output.n134 185
R22365 output.n114 output.n113 185
R22366 output.n129 output.n128 185
R22367 output.n127 output.n126 185
R22368 output.n118 output.n117 185
R22369 output.n121 output.n120 185
R22370 output.t19 output.n24 147.661
R22371 output.t0 output.n55 147.661
R22372 output.t17 output.n87 147.661
R22373 output.t18 output.n119 147.661
R22374 output.n41 output.n40 104.615
R22375 output.n40 output.n18 104.615
R22376 output.n33 output.n18 104.615
R22377 output.n33 output.n32 104.615
R22378 output.n32 output.n22 104.615
R22379 output.n25 output.n22 104.615
R22380 output.n72 output.n71 104.615
R22381 output.n71 output.n49 104.615
R22382 output.n64 output.n49 104.615
R22383 output.n64 output.n63 104.615
R22384 output.n63 output.n53 104.615
R22385 output.n56 output.n53 104.615
R22386 output.n104 output.n103 104.615
R22387 output.n103 output.n81 104.615
R22388 output.n96 output.n81 104.615
R22389 output.n96 output.n95 104.615
R22390 output.n95 output.n85 104.615
R22391 output.n88 output.n85 104.615
R22392 output.n136 output.n135 104.615
R22393 output.n135 output.n113 104.615
R22394 output.n128 output.n113 104.615
R22395 output.n128 output.n127 104.615
R22396 output.n127 output.n117 104.615
R22397 output.n120 output.n117 104.615
R22398 output.n1 output.t9 77.056
R22399 output.n14 output.t11 76.6694
R22400 output.n1 output.n0 72.7095
R22401 output.n3 output.n2 72.7095
R22402 output.n5 output.n4 72.7095
R22403 output.n7 output.n6 72.7095
R22404 output.n9 output.n8 72.7095
R22405 output.n11 output.n10 72.7095
R22406 output.n13 output.n12 72.7095
R22407 output.n25 output.t19 52.3082
R22408 output.n56 output.t0 52.3082
R22409 output.n88 output.t17 52.3082
R22410 output.n120 output.t18 52.3082
R22411 output.n26 output.n24 15.6674
R22412 output.n57 output.n55 15.6674
R22413 output.n89 output.n87 15.6674
R22414 output.n121 output.n119 15.6674
R22415 output.n27 output.n23 12.8005
R22416 output.n58 output.n54 12.8005
R22417 output.n90 output.n86 12.8005
R22418 output.n122 output.n118 12.8005
R22419 output.n31 output.n30 12.0247
R22420 output.n62 output.n61 12.0247
R22421 output.n94 output.n93 12.0247
R22422 output.n126 output.n125 12.0247
R22423 output.n34 output.n21 11.249
R22424 output.n65 output.n52 11.249
R22425 output.n97 output.n84 11.249
R22426 output.n129 output.n116 11.249
R22427 output.n35 output.n19 10.4732
R22428 output.n66 output.n50 10.4732
R22429 output.n98 output.n82 10.4732
R22430 output.n130 output.n114 10.4732
R22431 output.n39 output.n38 9.69747
R22432 output.n70 output.n69 9.69747
R22433 output.n102 output.n101 9.69747
R22434 output.n134 output.n133 9.69747
R22435 output.n45 output.n44 9.45567
R22436 output.n76 output.n75 9.45567
R22437 output.n108 output.n107 9.45567
R22438 output.n140 output.n139 9.45567
R22439 output.n44 output.n43 9.3005
R22440 output.n17 output.n16 9.3005
R22441 output.n38 output.n37 9.3005
R22442 output.n36 output.n35 9.3005
R22443 output.n21 output.n20 9.3005
R22444 output.n30 output.n29 9.3005
R22445 output.n28 output.n27 9.3005
R22446 output.n75 output.n74 9.3005
R22447 output.n48 output.n47 9.3005
R22448 output.n69 output.n68 9.3005
R22449 output.n67 output.n66 9.3005
R22450 output.n52 output.n51 9.3005
R22451 output.n61 output.n60 9.3005
R22452 output.n59 output.n58 9.3005
R22453 output.n107 output.n106 9.3005
R22454 output.n80 output.n79 9.3005
R22455 output.n101 output.n100 9.3005
R22456 output.n99 output.n98 9.3005
R22457 output.n84 output.n83 9.3005
R22458 output.n93 output.n92 9.3005
R22459 output.n91 output.n90 9.3005
R22460 output.n139 output.n138 9.3005
R22461 output.n112 output.n111 9.3005
R22462 output.n133 output.n132 9.3005
R22463 output.n131 output.n130 9.3005
R22464 output.n116 output.n115 9.3005
R22465 output.n125 output.n124 9.3005
R22466 output.n123 output.n122 9.3005
R22467 output.n42 output.n17 8.92171
R22468 output.n73 output.n48 8.92171
R22469 output.n105 output.n80 8.92171
R22470 output.n137 output.n112 8.92171
R22471 output output.n141 8.15037
R22472 output.n43 output.n15 8.14595
R22473 output.n74 output.n46 8.14595
R22474 output.n106 output.n78 8.14595
R22475 output.n138 output.n110 8.14595
R22476 output.n45 output.n15 5.81868
R22477 output.n76 output.n46 5.81868
R22478 output.n108 output.n78 5.81868
R22479 output.n140 output.n110 5.81868
R22480 output.n43 output.n42 5.04292
R22481 output.n74 output.n73 5.04292
R22482 output.n106 output.n105 5.04292
R22483 output.n138 output.n137 5.04292
R22484 output.n28 output.n24 4.38594
R22485 output.n59 output.n55 4.38594
R22486 output.n91 output.n87 4.38594
R22487 output.n123 output.n119 4.38594
R22488 output.n39 output.n17 4.26717
R22489 output.n70 output.n48 4.26717
R22490 output.n102 output.n80 4.26717
R22491 output.n134 output.n112 4.26717
R22492 output.n0 output.t5 3.9605
R22493 output.n0 output.t3 3.9605
R22494 output.n2 output.t13 3.9605
R22495 output.n2 output.t15 3.9605
R22496 output.n4 output.t16 3.9605
R22497 output.n4 output.t7 3.9605
R22498 output.n6 output.t10 3.9605
R22499 output.n6 output.t14 3.9605
R22500 output.n8 output.t1 3.9605
R22501 output.n8 output.t6 3.9605
R22502 output.n10 output.t8 3.9605
R22503 output.n10 output.t12 3.9605
R22504 output.n12 output.t4 3.9605
R22505 output.n12 output.t2 3.9605
R22506 output.n38 output.n19 3.49141
R22507 output.n69 output.n50 3.49141
R22508 output.n101 output.n82 3.49141
R22509 output.n133 output.n114 3.49141
R22510 output.n35 output.n34 2.71565
R22511 output.n66 output.n65 2.71565
R22512 output.n98 output.n97 2.71565
R22513 output.n130 output.n129 2.71565
R22514 output.n31 output.n21 1.93989
R22515 output.n62 output.n52 1.93989
R22516 output.n94 output.n84 1.93989
R22517 output.n126 output.n116 1.93989
R22518 output.n30 output.n23 1.16414
R22519 output.n61 output.n54 1.16414
R22520 output.n93 output.n86 1.16414
R22521 output.n125 output.n118 1.16414
R22522 output.n141 output.n109 0.962709
R22523 output.n109 output.n77 0.962709
R22524 output.n27 output.n26 0.388379
R22525 output.n58 output.n57 0.388379
R22526 output.n90 output.n89 0.388379
R22527 output.n122 output.n121 0.388379
R22528 output.n14 output.n13 0.387128
R22529 output.n13 output.n11 0.387128
R22530 output.n11 output.n9 0.387128
R22531 output.n9 output.n7 0.387128
R22532 output.n7 output.n5 0.387128
R22533 output.n5 output.n3 0.387128
R22534 output.n3 output.n1 0.387128
R22535 output.n44 output.n16 0.155672
R22536 output.n37 output.n16 0.155672
R22537 output.n37 output.n36 0.155672
R22538 output.n36 output.n20 0.155672
R22539 output.n29 output.n20 0.155672
R22540 output.n29 output.n28 0.155672
R22541 output.n75 output.n47 0.155672
R22542 output.n68 output.n47 0.155672
R22543 output.n68 output.n67 0.155672
R22544 output.n67 output.n51 0.155672
R22545 output.n60 output.n51 0.155672
R22546 output.n60 output.n59 0.155672
R22547 output.n107 output.n79 0.155672
R22548 output.n100 output.n79 0.155672
R22549 output.n100 output.n99 0.155672
R22550 output.n99 output.n83 0.155672
R22551 output.n92 output.n83 0.155672
R22552 output.n92 output.n91 0.155672
R22553 output.n139 output.n111 0.155672
R22554 output.n132 output.n111 0.155672
R22555 output.n132 output.n131 0.155672
R22556 output.n131 output.n115 0.155672
R22557 output.n124 output.n115 0.155672
R22558 output.n124 output.n123 0.155672
R22559 output output.n14 0.126227
R22560 plus.n46 plus.t9 252.611
R22561 plus.n9 plus.t11 252.611
R22562 plus.n76 plus.t4 243.97
R22563 plus.n72 plus.t12 231.093
R22564 plus.n35 plus.t7 231.093
R22565 plus.n76 plus.n75 223.454
R22566 plus.n78 plus.n77 223.454
R22567 plus.n47 plus.t5 187.445
R22568 plus.n44 plus.t18 187.445
R22569 plus.n42 plus.t17 187.445
R22570 plus.n59 plus.t13 187.445
R22571 plus.n65 plus.t14 187.445
R22572 plus.n38 plus.t10 187.445
R22573 plus.n1 plus.t6 187.445
R22574 plus.n28 plus.t16 187.445
R22575 plus.n22 plus.t15 187.445
R22576 plus.n5 plus.t20 187.445
R22577 plus.n7 plus.t19 187.445
R22578 plus.n10 plus.t8 187.445
R22579 plus.n73 plus.n72 161.3
R22580 plus.n71 plus.n37 161.3
R22581 plus.n70 plus.n69 161.3
R22582 plus.n68 plus.n67 161.3
R22583 plus.n66 plus.n39 161.3
R22584 plus.n64 plus.n63 161.3
R22585 plus.n62 plus.n40 161.3
R22586 plus.n61 plus.n60 161.3
R22587 plus.n58 plus.n41 161.3
R22588 plus.n57 plus.n56 161.3
R22589 plus.n55 plus.n54 161.3
R22590 plus.n53 plus.n43 161.3
R22591 plus.n52 plus.n51 161.3
R22592 plus.n50 plus.n49 161.3
R22593 plus.n48 plus.n45 161.3
R22594 plus.n11 plus.n8 161.3
R22595 plus.n13 plus.n12 161.3
R22596 plus.n15 plus.n14 161.3
R22597 plus.n16 plus.n6 161.3
R22598 plus.n18 plus.n17 161.3
R22599 plus.n20 plus.n19 161.3
R22600 plus.n21 plus.n4 161.3
R22601 plus.n24 plus.n23 161.3
R22602 plus.n25 plus.n3 161.3
R22603 plus.n27 plus.n26 161.3
R22604 plus.n29 plus.n2 161.3
R22605 plus.n31 plus.n30 161.3
R22606 plus.n33 plus.n32 161.3
R22607 plus.n34 plus.n0 161.3
R22608 plus.n36 plus.n35 161.3
R22609 plus.n49 plus.n48 56.5617
R22610 plus.n58 plus.n57 56.5617
R22611 plus.n67 plus.n66 56.5617
R22612 plus.n30 plus.n29 56.5617
R22613 plus.n21 plus.n20 56.5617
R22614 plus.n12 plus.n11 56.5617
R22615 plus.n71 plus.n70 46.3896
R22616 plus.n34 plus.n33 46.3896
R22617 plus.n46 plus.n45 42.8164
R22618 plus.n9 plus.n8 42.8164
R22619 plus.n54 plus.n53 42.5146
R22620 plus.n60 plus.n40 42.5146
R22621 plus.n23 plus.n3 42.5146
R22622 plus.n17 plus.n16 42.5146
R22623 plus.n53 plus.n52 38.6395
R22624 plus.n64 plus.n40 38.6395
R22625 plus.n27 plus.n3 38.6395
R22626 plus.n16 plus.n15 38.6395
R22627 plus.n47 plus.n46 38.2514
R22628 plus.n10 plus.n9 38.2514
R22629 plus.n74 plus.n73 31.491
R22630 plus.n49 plus.n44 19.9199
R22631 plus.n66 plus.n65 19.9199
R22632 plus.n29 plus.n28 19.9199
R22633 plus.n12 plus.n7 19.9199
R22634 plus.n75 plus.t1 19.8005
R22635 plus.n75 plus.t2 19.8005
R22636 plus.n77 plus.t0 19.8005
R22637 plus.n77 plus.t3 19.8005
R22638 plus.n57 plus.n42 17.9525
R22639 plus.n59 plus.n58 17.9525
R22640 plus.n22 plus.n21 17.9525
R22641 plus.n20 plus.n5 17.9525
R22642 plus.n48 plus.n47 15.9852
R22643 plus.n67 plus.n38 15.9852
R22644 plus.n30 plus.n1 15.9852
R22645 plus.n11 plus.n10 15.9852
R22646 plus.n72 plus.n71 15.3369
R22647 plus.n35 plus.n34 15.3369
R22648 plus plus.n79 14.5081
R22649 plus.n74 plus.n36 11.9494
R22650 plus.n70 plus.n38 8.60764
R22651 plus.n33 plus.n1 8.60764
R22652 plus.n54 plus.n42 6.6403
R22653 plus.n60 plus.n59 6.6403
R22654 plus.n23 plus.n22 6.6403
R22655 plus.n17 plus.n5 6.6403
R22656 plus.n79 plus.n78 5.40567
R22657 plus.n52 plus.n44 4.67295
R22658 plus.n65 plus.n64 4.67295
R22659 plus.n28 plus.n27 4.67295
R22660 plus.n15 plus.n7 4.67295
R22661 plus.n79 plus.n74 1.188
R22662 plus.n78 plus.n76 0.716017
R22663 plus.n50 plus.n45 0.189894
R22664 plus.n51 plus.n50 0.189894
R22665 plus.n51 plus.n43 0.189894
R22666 plus.n55 plus.n43 0.189894
R22667 plus.n56 plus.n55 0.189894
R22668 plus.n56 plus.n41 0.189894
R22669 plus.n61 plus.n41 0.189894
R22670 plus.n62 plus.n61 0.189894
R22671 plus.n63 plus.n62 0.189894
R22672 plus.n63 plus.n39 0.189894
R22673 plus.n68 plus.n39 0.189894
R22674 plus.n69 plus.n68 0.189894
R22675 plus.n69 plus.n37 0.189894
R22676 plus.n73 plus.n37 0.189894
R22677 plus.n36 plus.n0 0.189894
R22678 plus.n32 plus.n0 0.189894
R22679 plus.n32 plus.n31 0.189894
R22680 plus.n31 plus.n2 0.189894
R22681 plus.n26 plus.n2 0.189894
R22682 plus.n26 plus.n25 0.189894
R22683 plus.n25 plus.n24 0.189894
R22684 plus.n24 plus.n4 0.189894
R22685 plus.n19 plus.n4 0.189894
R22686 plus.n19 plus.n18 0.189894
R22687 plus.n18 plus.n6 0.189894
R22688 plus.n14 plus.n6 0.189894
R22689 plus.n14 plus.n13 0.189894
R22690 plus.n13 plus.n8 0.189894
R22691 a_n2903_n3924.n0 a_n2903_n3924.t35 214.981
R22692 a_n2903_n3924.n2 a_n2903_n3924.t31 214.452
R22693 a_n2903_n3924.n11 a_n2903_n3924.t36 214.321
R22694 a_n2903_n3924.n12 a_n2903_n3924.t39 214.321
R22695 a_n2903_n3924.n13 a_n2903_n3924.t38 214.321
R22696 a_n2903_n3924.n14 a_n2903_n3924.t27 214.321
R22697 a_n2903_n3924.n15 a_n2903_n3924.t21 214.321
R22698 a_n2903_n3924.n0 a_n2903_n3924.t20 214.321
R22699 a_n2903_n3924.n1 a_n2903_n3924.t14 55.8337
R22700 a_n2903_n3924.n3 a_n2903_n3924.t22 55.8337
R22701 a_n2903_n3924.n10 a_n2903_n3924.t0 55.8337
R22702 a_n2903_n3924.n34 a_n2903_n3924.t11 55.8335
R22703 a_n2903_n3924.n32 a_n2903_n3924.t37 55.8335
R22704 a_n2903_n3924.n25 a_n2903_n3924.t2 55.8335
R22705 a_n2903_n3924.n24 a_n2903_n3924.t12 55.8335
R22706 a_n2903_n3924.n17 a_n2903_n3924.t16 55.8335
R22707 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0052
R22708 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0052
R22709 a_n2903_n3924.n5 a_n2903_n3924.n4 53.0052
R22710 a_n2903_n3924.n7 a_n2903_n3924.n6 53.0052
R22711 a_n2903_n3924.n9 a_n2903_n3924.n8 53.0052
R22712 a_n2903_n3924.n31 a_n2903_n3924.n30 53.0051
R22713 a_n2903_n3924.n29 a_n2903_n3924.n28 53.0051
R22714 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R22715 a_n2903_n3924.n23 a_n2903_n3924.n22 53.0051
R22716 a_n2903_n3924.n21 a_n2903_n3924.n20 53.0051
R22717 a_n2903_n3924.n19 a_n2903_n3924.n18 53.0051
R22718 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R22719 a_n2903_n3924.n16 a_n2903_n3924.n10 12.2417
R22720 a_n2903_n3924.n34 a_n2903_n3924.n33 12.2417
R22721 a_n2903_n3924.n17 a_n2903_n3924.n16 5.16214
R22722 a_n2903_n3924.n33 a_n2903_n3924.n32 5.16214
R22723 a_n2903_n3924.n35 a_n2903_n3924.t9 2.82907
R22724 a_n2903_n3924.n35 a_n2903_n3924.t13 2.82907
R22725 a_n2903_n3924.n37 a_n2903_n3924.t6 2.82907
R22726 a_n2903_n3924.n37 a_n2903_n3924.t10 2.82907
R22727 a_n2903_n3924.n4 a_n2903_n3924.t24 2.82907
R22728 a_n2903_n3924.n4 a_n2903_n3924.t19 2.82907
R22729 a_n2903_n3924.n6 a_n2903_n3924.t30 2.82907
R22730 a_n2903_n3924.n6 a_n2903_n3924.t32 2.82907
R22731 a_n2903_n3924.n8 a_n2903_n3924.t1 2.82907
R22732 a_n2903_n3924.n8 a_n2903_n3924.t29 2.82907
R22733 a_n2903_n3924.n30 a_n2903_n3924.t34 2.82907
R22734 a_n2903_n3924.n30 a_n2903_n3924.t28 2.82907
R22735 a_n2903_n3924.n28 a_n2903_n3924.t25 2.82907
R22736 a_n2903_n3924.n28 a_n2903_n3924.t33 2.82907
R22737 a_n2903_n3924.n26 a_n2903_n3924.t26 2.82907
R22738 a_n2903_n3924.n26 a_n2903_n3924.t23 2.82907
R22739 a_n2903_n3924.n22 a_n2903_n3924.t4 2.82907
R22740 a_n2903_n3924.n22 a_n2903_n3924.t15 2.82907
R22741 a_n2903_n3924.n20 a_n2903_n3924.t8 2.82907
R22742 a_n2903_n3924.n20 a_n2903_n3924.t3 2.82907
R22743 a_n2903_n3924.n18 a_n2903_n3924.t17 2.82907
R22744 a_n2903_n3924.n18 a_n2903_n3924.t7 2.82907
R22745 a_n2903_n3924.t18 a_n2903_n3924.n40 2.82907
R22746 a_n2903_n3924.n40 a_n2903_n3924.t5 2.82907
R22747 a_n2903_n3924.n33 a_n2903_n3924.n2 1.95694
R22748 a_n2903_n3924.n16 a_n2903_n3924.n0 1.95694
R22749 a_n2903_n3924.n0 a_n2903_n3924.n15 0.684366
R22750 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R22751 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R22752 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R22753 a_n2903_n3924.n12 a_n2903_n3924.n11 0.672012
R22754 a_n2903_n3924.n11 a_n2903_n3924.n2 0.541924
R22755 a_n2903_n3924.n19 a_n2903_n3924.n17 0.530672
R22756 a_n2903_n3924.n21 a_n2903_n3924.n19 0.530672
R22757 a_n2903_n3924.n23 a_n2903_n3924.n21 0.530672
R22758 a_n2903_n3924.n24 a_n2903_n3924.n23 0.530672
R22759 a_n2903_n3924.n27 a_n2903_n3924.n25 0.530672
R22760 a_n2903_n3924.n29 a_n2903_n3924.n27 0.530672
R22761 a_n2903_n3924.n31 a_n2903_n3924.n29 0.530672
R22762 a_n2903_n3924.n32 a_n2903_n3924.n31 0.530672
R22763 a_n2903_n3924.n10 a_n2903_n3924.n9 0.530672
R22764 a_n2903_n3924.n9 a_n2903_n3924.n7 0.530672
R22765 a_n2903_n3924.n7 a_n2903_n3924.n5 0.530672
R22766 a_n2903_n3924.n5 a_n2903_n3924.n3 0.530672
R22767 a_n2903_n3924.n39 a_n2903_n3924.n1 0.530672
R22768 a_n2903_n3924.n39 a_n2903_n3924.n38 0.530672
R22769 a_n2903_n3924.n38 a_n2903_n3924.n36 0.530672
R22770 a_n2903_n3924.n36 a_n2903_n3924.n34 0.530672
R22771 a_n2903_n3924.n25 a_n2903_n3924.n24 0.235414
R22772 a_n2903_n3924.n3 a_n2903_n3924.n1 0.235414
R22773 minus.n46 minus.t20 252.611
R22774 minus.n9 minus.t13 252.611
R22775 minus.n78 minus.t3 243.255
R22776 minus.n72 minus.t15 231.093
R22777 minus.n35 minus.t17 231.093
R22778 minus.n77 minus.n75 224.169
R22779 minus.n77 minus.n76 223.454
R22780 minus.n38 minus.t12 187.445
R22781 minus.n65 minus.t7 187.445
R22782 minus.n59 minus.t6 187.445
R22783 minus.n42 minus.t11 187.445
R22784 minus.n44 minus.t10 187.445
R22785 minus.n47 minus.t16 187.445
R22786 minus.n10 minus.t9 187.445
R22787 minus.n7 minus.t8 187.445
R22788 minus.n5 minus.t5 187.445
R22789 minus.n22 minus.t18 187.445
R22790 minus.n28 minus.t19 187.445
R22791 minus.n1 minus.t14 187.445
R22792 minus.n48 minus.n45 161.3
R22793 minus.n50 minus.n49 161.3
R22794 minus.n52 minus.n51 161.3
R22795 minus.n53 minus.n43 161.3
R22796 minus.n55 minus.n54 161.3
R22797 minus.n57 minus.n56 161.3
R22798 minus.n58 minus.n41 161.3
R22799 minus.n61 minus.n60 161.3
R22800 minus.n62 minus.n40 161.3
R22801 minus.n64 minus.n63 161.3
R22802 minus.n66 minus.n39 161.3
R22803 minus.n68 minus.n67 161.3
R22804 minus.n70 minus.n69 161.3
R22805 minus.n71 minus.n37 161.3
R22806 minus.n73 minus.n72 161.3
R22807 minus.n36 minus.n35 161.3
R22808 minus.n34 minus.n0 161.3
R22809 minus.n33 minus.n32 161.3
R22810 minus.n31 minus.n30 161.3
R22811 minus.n29 minus.n2 161.3
R22812 minus.n27 minus.n26 161.3
R22813 minus.n25 minus.n3 161.3
R22814 minus.n24 minus.n23 161.3
R22815 minus.n21 minus.n4 161.3
R22816 minus.n20 minus.n19 161.3
R22817 minus.n18 minus.n17 161.3
R22818 minus.n16 minus.n6 161.3
R22819 minus.n15 minus.n14 161.3
R22820 minus.n13 minus.n12 161.3
R22821 minus.n11 minus.n8 161.3
R22822 minus.n67 minus.n66 56.5617
R22823 minus.n58 minus.n57 56.5617
R22824 minus.n49 minus.n48 56.5617
R22825 minus.n12 minus.n11 56.5617
R22826 minus.n21 minus.n20 56.5617
R22827 minus.n30 minus.n29 56.5617
R22828 minus.n71 minus.n70 46.3896
R22829 minus.n34 minus.n33 46.3896
R22830 minus.n46 minus.n45 42.8164
R22831 minus.n9 minus.n8 42.8164
R22832 minus.n60 minus.n40 42.5146
R22833 minus.n54 minus.n53 42.5146
R22834 minus.n17 minus.n16 42.5146
R22835 minus.n23 minus.n3 42.5146
R22836 minus.n64 minus.n40 38.6395
R22837 minus.n53 minus.n52 38.6395
R22838 minus.n16 minus.n15 38.6395
R22839 minus.n27 minus.n3 38.6395
R22840 minus.n47 minus.n46 38.2514
R22841 minus.n10 minus.n9 38.2514
R22842 minus.n74 minus.n73 31.7069
R22843 minus.n66 minus.n65 19.9199
R22844 minus.n49 minus.n44 19.9199
R22845 minus.n12 minus.n7 19.9199
R22846 minus.n29 minus.n28 19.9199
R22847 minus.n76 minus.t2 19.8005
R22848 minus.n76 minus.t0 19.8005
R22849 minus.n75 minus.t1 19.8005
R22850 minus.n75 minus.t4 19.8005
R22851 minus.n59 minus.n58 17.9525
R22852 minus.n57 minus.n42 17.9525
R22853 minus.n20 minus.n5 17.9525
R22854 minus.n22 minus.n21 17.9525
R22855 minus.n67 minus.n38 15.9852
R22856 minus.n48 minus.n47 15.9852
R22857 minus.n11 minus.n10 15.9852
R22858 minus.n30 minus.n1 15.9852
R22859 minus.n72 minus.n71 15.3369
R22860 minus.n35 minus.n34 15.3369
R22861 minus.n74 minus.n36 12.1653
R22862 minus minus.n79 11.6359
R22863 minus.n70 minus.n38 8.60764
R22864 minus.n33 minus.n1 8.60764
R22865 minus.n60 minus.n59 6.6403
R22866 minus.n54 minus.n42 6.6403
R22867 minus.n17 minus.n5 6.6403
R22868 minus.n23 minus.n22 6.6403
R22869 minus.n79 minus.n78 4.80222
R22870 minus.n65 minus.n64 4.67295
R22871 minus.n52 minus.n44 4.67295
R22872 minus.n15 minus.n7 4.67295
R22873 minus.n28 minus.n27 4.67295
R22874 minus.n79 minus.n74 0.972091
R22875 minus.n78 minus.n77 0.716017
R22876 minus.n73 minus.n37 0.189894
R22877 minus.n69 minus.n37 0.189894
R22878 minus.n69 minus.n68 0.189894
R22879 minus.n68 minus.n39 0.189894
R22880 minus.n63 minus.n39 0.189894
R22881 minus.n63 minus.n62 0.189894
R22882 minus.n62 minus.n61 0.189894
R22883 minus.n61 minus.n41 0.189894
R22884 minus.n56 minus.n41 0.189894
R22885 minus.n56 minus.n55 0.189894
R22886 minus.n55 minus.n43 0.189894
R22887 minus.n51 minus.n43 0.189894
R22888 minus.n51 minus.n50 0.189894
R22889 minus.n50 minus.n45 0.189894
R22890 minus.n13 minus.n8 0.189894
R22891 minus.n14 minus.n13 0.189894
R22892 minus.n14 minus.n6 0.189894
R22893 minus.n18 minus.n6 0.189894
R22894 minus.n19 minus.n18 0.189894
R22895 minus.n19 minus.n4 0.189894
R22896 minus.n24 minus.n4 0.189894
R22897 minus.n25 minus.n24 0.189894
R22898 minus.n26 minus.n25 0.189894
R22899 minus.n26 minus.n2 0.189894
R22900 minus.n31 minus.n2 0.189894
R22901 minus.n32 minus.n31 0.189894
R22902 minus.n32 minus.n0 0.189894
R22903 minus.n36 minus.n0 0.189894
R22904 a_n2982_8322.n12 a_n2982_8322.t33 74.6477
R22905 a_n2982_8322.n1 a_n2982_8322.t12 74.6477
R22906 a_n2982_8322.n28 a_n2982_8322.t27 74.6474
R22907 a_n2982_8322.n20 a_n2982_8322.t7 74.2899
R22908 a_n2982_8322.n13 a_n2982_8322.t31 74.2899
R22909 a_n2982_8322.n14 a_n2982_8322.t34 74.2899
R22910 a_n2982_8322.n17 a_n2982_8322.t35 74.2899
R22911 a_n2982_8322.n10 a_n2982_8322.t6 74.2899
R22912 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R22913 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R22914 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R22915 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R22916 a_n2982_8322.n12 a_n2982_8322.n11 70.6783
R22917 a_n2982_8322.n16 a_n2982_8322.n15 70.6783
R22918 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R22919 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R22920 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R22921 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R22922 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R22923 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R22924 a_n2982_8322.n18 a_n2982_8322.n10 24.9022
R22925 a_n2982_8322.n19 a_n2982_8322.t0 9.69161
R22926 a_n2982_8322.n18 a_n2982_8322.n17 8.38735
R22927 a_n2982_8322.n20 a_n2982_8322.n19 6.90998
R22928 a_n2982_8322.n19 a_n2982_8322.n18 5.3452
R22929 a_n2982_8322.n27 a_n2982_8322.t20 3.61217
R22930 a_n2982_8322.n27 a_n2982_8322.t16 3.61217
R22931 a_n2982_8322.n25 a_n2982_8322.t26 3.61217
R22932 a_n2982_8322.n25 a_n2982_8322.t14 3.61217
R22933 a_n2982_8322.n23 a_n2982_8322.t11 3.61217
R22934 a_n2982_8322.n23 a_n2982_8322.t10 3.61217
R22935 a_n2982_8322.n21 a_n2982_8322.t24 3.61217
R22936 a_n2982_8322.n21 a_n2982_8322.t23 3.61217
R22937 a_n2982_8322.n11 a_n2982_8322.t37 3.61217
R22938 a_n2982_8322.n11 a_n2982_8322.t36 3.61217
R22939 a_n2982_8322.n15 a_n2982_8322.t32 3.61217
R22940 a_n2982_8322.n15 a_n2982_8322.t30 3.61217
R22941 a_n2982_8322.n0 a_n2982_8322.t25 3.61217
R22942 a_n2982_8322.n0 a_n2982_8322.t21 3.61217
R22943 a_n2982_8322.n2 a_n2982_8322.t28 3.61217
R22944 a_n2982_8322.n2 a_n2982_8322.t18 3.61217
R22945 a_n2982_8322.n4 a_n2982_8322.t9 3.61217
R22946 a_n2982_8322.n4 a_n2982_8322.t8 3.61217
R22947 a_n2982_8322.n6 a_n2982_8322.t22 3.61217
R22948 a_n2982_8322.n6 a_n2982_8322.t15 3.61217
R22949 a_n2982_8322.n8 a_n2982_8322.t19 3.61217
R22950 a_n2982_8322.n8 a_n2982_8322.t17 3.61217
R22951 a_n2982_8322.n30 a_n2982_8322.t13 3.61217
R22952 a_n2982_8322.t29 a_n2982_8322.n30 3.61217
R22953 a_n2982_8322.n17 a_n2982_8322.n16 0.358259
R22954 a_n2982_8322.n16 a_n2982_8322.n14 0.358259
R22955 a_n2982_8322.n13 a_n2982_8322.n12 0.358259
R22956 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R22957 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R22958 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R22959 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R22960 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R22961 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R22962 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R22963 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R22964 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R22965 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R22966 a_n2982_8322.n14 a_n2982_8322.n13 0.101793
R22967 a_n2982_8322.t5 a_n2982_8322.t1 0.0788333
R22968 a_n2982_8322.t4 a_n2982_8322.t2 0.0788333
R22969 a_n2982_8322.t0 a_n2982_8322.t3 0.0788333
R22970 a_n2982_8322.t4 a_n2982_8322.t5 0.0318333
R22971 a_n2982_8322.t0 a_n2982_8322.t2 0.0318333
R22972 a_n2982_8322.t1 a_n2982_8322.t2 0.0318333
R22973 a_n2982_8322.t3 a_n2982_8322.t4 0.0318333
R22974 outputibias.n27 outputibias.n1 289.615
R22975 outputibias.n58 outputibias.n32 289.615
R22976 outputibias.n90 outputibias.n64 289.615
R22977 outputibias.n122 outputibias.n96 289.615
R22978 outputibias.n28 outputibias.n27 185
R22979 outputibias.n26 outputibias.n25 185
R22980 outputibias.n5 outputibias.n4 185
R22981 outputibias.n20 outputibias.n19 185
R22982 outputibias.n18 outputibias.n17 185
R22983 outputibias.n9 outputibias.n8 185
R22984 outputibias.n12 outputibias.n11 185
R22985 outputibias.n59 outputibias.n58 185
R22986 outputibias.n57 outputibias.n56 185
R22987 outputibias.n36 outputibias.n35 185
R22988 outputibias.n51 outputibias.n50 185
R22989 outputibias.n49 outputibias.n48 185
R22990 outputibias.n40 outputibias.n39 185
R22991 outputibias.n43 outputibias.n42 185
R22992 outputibias.n91 outputibias.n90 185
R22993 outputibias.n89 outputibias.n88 185
R22994 outputibias.n68 outputibias.n67 185
R22995 outputibias.n83 outputibias.n82 185
R22996 outputibias.n81 outputibias.n80 185
R22997 outputibias.n72 outputibias.n71 185
R22998 outputibias.n75 outputibias.n74 185
R22999 outputibias.n123 outputibias.n122 185
R23000 outputibias.n121 outputibias.n120 185
R23001 outputibias.n100 outputibias.n99 185
R23002 outputibias.n115 outputibias.n114 185
R23003 outputibias.n113 outputibias.n112 185
R23004 outputibias.n104 outputibias.n103 185
R23005 outputibias.n107 outputibias.n106 185
R23006 outputibias.n0 outputibias.t10 178.945
R23007 outputibias.n133 outputibias.t9 177.018
R23008 outputibias.n132 outputibias.t11 177.018
R23009 outputibias.n0 outputibias.t8 177.018
R23010 outputibias.t7 outputibias.n10 147.661
R23011 outputibias.t1 outputibias.n41 147.661
R23012 outputibias.t5 outputibias.n73 147.661
R23013 outputibias.t3 outputibias.n105 147.661
R23014 outputibias.n128 outputibias.t6 132.363
R23015 outputibias.n128 outputibias.t0 130.436
R23016 outputibias.n129 outputibias.t4 130.436
R23017 outputibias.n130 outputibias.t2 130.436
R23018 outputibias.n27 outputibias.n26 104.615
R23019 outputibias.n26 outputibias.n4 104.615
R23020 outputibias.n19 outputibias.n4 104.615
R23021 outputibias.n19 outputibias.n18 104.615
R23022 outputibias.n18 outputibias.n8 104.615
R23023 outputibias.n11 outputibias.n8 104.615
R23024 outputibias.n58 outputibias.n57 104.615
R23025 outputibias.n57 outputibias.n35 104.615
R23026 outputibias.n50 outputibias.n35 104.615
R23027 outputibias.n50 outputibias.n49 104.615
R23028 outputibias.n49 outputibias.n39 104.615
R23029 outputibias.n42 outputibias.n39 104.615
R23030 outputibias.n90 outputibias.n89 104.615
R23031 outputibias.n89 outputibias.n67 104.615
R23032 outputibias.n82 outputibias.n67 104.615
R23033 outputibias.n82 outputibias.n81 104.615
R23034 outputibias.n81 outputibias.n71 104.615
R23035 outputibias.n74 outputibias.n71 104.615
R23036 outputibias.n122 outputibias.n121 104.615
R23037 outputibias.n121 outputibias.n99 104.615
R23038 outputibias.n114 outputibias.n99 104.615
R23039 outputibias.n114 outputibias.n113 104.615
R23040 outputibias.n113 outputibias.n103 104.615
R23041 outputibias.n106 outputibias.n103 104.615
R23042 outputibias.n63 outputibias.n31 95.6354
R23043 outputibias.n63 outputibias.n62 94.6732
R23044 outputibias.n95 outputibias.n94 94.6732
R23045 outputibias.n127 outputibias.n126 94.6732
R23046 outputibias.n11 outputibias.t7 52.3082
R23047 outputibias.n42 outputibias.t1 52.3082
R23048 outputibias.n74 outputibias.t5 52.3082
R23049 outputibias.n106 outputibias.t3 52.3082
R23050 outputibias.n12 outputibias.n10 15.6674
R23051 outputibias.n43 outputibias.n41 15.6674
R23052 outputibias.n75 outputibias.n73 15.6674
R23053 outputibias.n107 outputibias.n105 15.6674
R23054 outputibias.n13 outputibias.n9 12.8005
R23055 outputibias.n44 outputibias.n40 12.8005
R23056 outputibias.n76 outputibias.n72 12.8005
R23057 outputibias.n108 outputibias.n104 12.8005
R23058 outputibias.n17 outputibias.n16 12.0247
R23059 outputibias.n48 outputibias.n47 12.0247
R23060 outputibias.n80 outputibias.n79 12.0247
R23061 outputibias.n112 outputibias.n111 12.0247
R23062 outputibias.n20 outputibias.n7 11.249
R23063 outputibias.n51 outputibias.n38 11.249
R23064 outputibias.n83 outputibias.n70 11.249
R23065 outputibias.n115 outputibias.n102 11.249
R23066 outputibias.n21 outputibias.n5 10.4732
R23067 outputibias.n52 outputibias.n36 10.4732
R23068 outputibias.n84 outputibias.n68 10.4732
R23069 outputibias.n116 outputibias.n100 10.4732
R23070 outputibias.n25 outputibias.n24 9.69747
R23071 outputibias.n56 outputibias.n55 9.69747
R23072 outputibias.n88 outputibias.n87 9.69747
R23073 outputibias.n120 outputibias.n119 9.69747
R23074 outputibias.n31 outputibias.n30 9.45567
R23075 outputibias.n62 outputibias.n61 9.45567
R23076 outputibias.n94 outputibias.n93 9.45567
R23077 outputibias.n126 outputibias.n125 9.45567
R23078 outputibias.n30 outputibias.n29 9.3005
R23079 outputibias.n3 outputibias.n2 9.3005
R23080 outputibias.n24 outputibias.n23 9.3005
R23081 outputibias.n22 outputibias.n21 9.3005
R23082 outputibias.n7 outputibias.n6 9.3005
R23083 outputibias.n16 outputibias.n15 9.3005
R23084 outputibias.n14 outputibias.n13 9.3005
R23085 outputibias.n61 outputibias.n60 9.3005
R23086 outputibias.n34 outputibias.n33 9.3005
R23087 outputibias.n55 outputibias.n54 9.3005
R23088 outputibias.n53 outputibias.n52 9.3005
R23089 outputibias.n38 outputibias.n37 9.3005
R23090 outputibias.n47 outputibias.n46 9.3005
R23091 outputibias.n45 outputibias.n44 9.3005
R23092 outputibias.n93 outputibias.n92 9.3005
R23093 outputibias.n66 outputibias.n65 9.3005
R23094 outputibias.n87 outputibias.n86 9.3005
R23095 outputibias.n85 outputibias.n84 9.3005
R23096 outputibias.n70 outputibias.n69 9.3005
R23097 outputibias.n79 outputibias.n78 9.3005
R23098 outputibias.n77 outputibias.n76 9.3005
R23099 outputibias.n125 outputibias.n124 9.3005
R23100 outputibias.n98 outputibias.n97 9.3005
R23101 outputibias.n119 outputibias.n118 9.3005
R23102 outputibias.n117 outputibias.n116 9.3005
R23103 outputibias.n102 outputibias.n101 9.3005
R23104 outputibias.n111 outputibias.n110 9.3005
R23105 outputibias.n109 outputibias.n108 9.3005
R23106 outputibias.n28 outputibias.n3 8.92171
R23107 outputibias.n59 outputibias.n34 8.92171
R23108 outputibias.n91 outputibias.n66 8.92171
R23109 outputibias.n123 outputibias.n98 8.92171
R23110 outputibias.n29 outputibias.n1 8.14595
R23111 outputibias.n60 outputibias.n32 8.14595
R23112 outputibias.n92 outputibias.n64 8.14595
R23113 outputibias.n124 outputibias.n96 8.14595
R23114 outputibias.n31 outputibias.n1 5.81868
R23115 outputibias.n62 outputibias.n32 5.81868
R23116 outputibias.n94 outputibias.n64 5.81868
R23117 outputibias.n126 outputibias.n96 5.81868
R23118 outputibias.n131 outputibias.n130 5.20947
R23119 outputibias.n29 outputibias.n28 5.04292
R23120 outputibias.n60 outputibias.n59 5.04292
R23121 outputibias.n92 outputibias.n91 5.04292
R23122 outputibias.n124 outputibias.n123 5.04292
R23123 outputibias.n131 outputibias.n127 4.42209
R23124 outputibias.n14 outputibias.n10 4.38594
R23125 outputibias.n45 outputibias.n41 4.38594
R23126 outputibias.n77 outputibias.n73 4.38594
R23127 outputibias.n109 outputibias.n105 4.38594
R23128 outputibias.n132 outputibias.n131 4.28454
R23129 outputibias.n25 outputibias.n3 4.26717
R23130 outputibias.n56 outputibias.n34 4.26717
R23131 outputibias.n88 outputibias.n66 4.26717
R23132 outputibias.n120 outputibias.n98 4.26717
R23133 outputibias.n24 outputibias.n5 3.49141
R23134 outputibias.n55 outputibias.n36 3.49141
R23135 outputibias.n87 outputibias.n68 3.49141
R23136 outputibias.n119 outputibias.n100 3.49141
R23137 outputibias.n21 outputibias.n20 2.71565
R23138 outputibias.n52 outputibias.n51 2.71565
R23139 outputibias.n84 outputibias.n83 2.71565
R23140 outputibias.n116 outputibias.n115 2.71565
R23141 outputibias.n17 outputibias.n7 1.93989
R23142 outputibias.n48 outputibias.n38 1.93989
R23143 outputibias.n80 outputibias.n70 1.93989
R23144 outputibias.n112 outputibias.n102 1.93989
R23145 outputibias.n130 outputibias.n129 1.9266
R23146 outputibias.n129 outputibias.n128 1.9266
R23147 outputibias.n133 outputibias.n132 1.92658
R23148 outputibias.n134 outputibias.n133 1.29913
R23149 outputibias.n16 outputibias.n9 1.16414
R23150 outputibias.n47 outputibias.n40 1.16414
R23151 outputibias.n79 outputibias.n72 1.16414
R23152 outputibias.n111 outputibias.n104 1.16414
R23153 outputibias.n127 outputibias.n95 0.962709
R23154 outputibias.n95 outputibias.n63 0.962709
R23155 outputibias.n13 outputibias.n12 0.388379
R23156 outputibias.n44 outputibias.n43 0.388379
R23157 outputibias.n76 outputibias.n75 0.388379
R23158 outputibias.n108 outputibias.n107 0.388379
R23159 outputibias.n134 outputibias.n0 0.337251
R23160 outputibias outputibias.n134 0.302375
R23161 outputibias.n30 outputibias.n2 0.155672
R23162 outputibias.n23 outputibias.n2 0.155672
R23163 outputibias.n23 outputibias.n22 0.155672
R23164 outputibias.n22 outputibias.n6 0.155672
R23165 outputibias.n15 outputibias.n6 0.155672
R23166 outputibias.n15 outputibias.n14 0.155672
R23167 outputibias.n61 outputibias.n33 0.155672
R23168 outputibias.n54 outputibias.n33 0.155672
R23169 outputibias.n54 outputibias.n53 0.155672
R23170 outputibias.n53 outputibias.n37 0.155672
R23171 outputibias.n46 outputibias.n37 0.155672
R23172 outputibias.n46 outputibias.n45 0.155672
R23173 outputibias.n93 outputibias.n65 0.155672
R23174 outputibias.n86 outputibias.n65 0.155672
R23175 outputibias.n86 outputibias.n85 0.155672
R23176 outputibias.n85 outputibias.n69 0.155672
R23177 outputibias.n78 outputibias.n69 0.155672
R23178 outputibias.n78 outputibias.n77 0.155672
R23179 outputibias.n125 outputibias.n97 0.155672
R23180 outputibias.n118 outputibias.n97 0.155672
R23181 outputibias.n118 outputibias.n117 0.155672
R23182 outputibias.n117 outputibias.n101 0.155672
R23183 outputibias.n110 outputibias.n101 0.155672
R23184 outputibias.n110 outputibias.n109 0.155672
R23185 diffpairibias.n0 diffpairibias.t18 436.822
R23186 diffpairibias.n21 diffpairibias.t19 435.479
R23187 diffpairibias.n20 diffpairibias.t16 435.479
R23188 diffpairibias.n19 diffpairibias.t17 435.479
R23189 diffpairibias.n18 diffpairibias.t21 435.479
R23190 diffpairibias.n0 diffpairibias.t22 435.479
R23191 diffpairibias.n1 diffpairibias.t20 435.479
R23192 diffpairibias.n2 diffpairibias.t23 435.479
R23193 diffpairibias.n10 diffpairibias.t0 377.536
R23194 diffpairibias.n10 diffpairibias.t8 376.193
R23195 diffpairibias.n11 diffpairibias.t10 376.193
R23196 diffpairibias.n12 diffpairibias.t6 376.193
R23197 diffpairibias.n13 diffpairibias.t2 376.193
R23198 diffpairibias.n14 diffpairibias.t12 376.193
R23199 diffpairibias.n15 diffpairibias.t4 376.193
R23200 diffpairibias.n16 diffpairibias.t14 376.193
R23201 diffpairibias.n3 diffpairibias.t1 113.368
R23202 diffpairibias.n3 diffpairibias.t9 112.698
R23203 diffpairibias.n4 diffpairibias.t11 112.698
R23204 diffpairibias.n5 diffpairibias.t7 112.698
R23205 diffpairibias.n6 diffpairibias.t3 112.698
R23206 diffpairibias.n7 diffpairibias.t13 112.698
R23207 diffpairibias.n8 diffpairibias.t5 112.698
R23208 diffpairibias.n9 diffpairibias.t15 112.698
R23209 diffpairibias.n17 diffpairibias.n16 4.77242
R23210 diffpairibias.n17 diffpairibias.n9 4.30807
R23211 diffpairibias.n18 diffpairibias.n17 4.13945
R23212 diffpairibias.n16 diffpairibias.n15 1.34352
R23213 diffpairibias.n15 diffpairibias.n14 1.34352
R23214 diffpairibias.n14 diffpairibias.n13 1.34352
R23215 diffpairibias.n13 diffpairibias.n12 1.34352
R23216 diffpairibias.n12 diffpairibias.n11 1.34352
R23217 diffpairibias.n11 diffpairibias.n10 1.34352
R23218 diffpairibias.n2 diffpairibias.n1 1.34352
R23219 diffpairibias.n1 diffpairibias.n0 1.34352
R23220 diffpairibias.n19 diffpairibias.n18 1.34352
R23221 diffpairibias.n20 diffpairibias.n19 1.34352
R23222 diffpairibias.n21 diffpairibias.n20 1.34352
R23223 diffpairibias.n22 diffpairibias.n21 0.862419
R23224 diffpairibias diffpairibias.n22 0.684875
R23225 diffpairibias.n9 diffpairibias.n8 0.672012
R23226 diffpairibias.n8 diffpairibias.n7 0.672012
R23227 diffpairibias.n7 diffpairibias.n6 0.672012
R23228 diffpairibias.n6 diffpairibias.n5 0.672012
R23229 diffpairibias.n5 diffpairibias.n4 0.672012
R23230 diffpairibias.n4 diffpairibias.n3 0.672012
R23231 diffpairibias.n22 diffpairibias.n2 0.190907
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.142351p
C5 minus diffpairibias 3.46e-19
C6 commonsourceibias output 0.006829f
C7 CSoutput minus 2.84082f
C8 vdd plus 0.100764f
C9 commonsourceibias outputibias 0.003902f
C10 plus diffpairibias 2.47e-19
C11 vdd commonsourceibias 0.004262f
C12 CSoutput plus 0.861671f
C13 commonsourceibias diffpairibias 0.052851f
C14 CSoutput commonsourceibias 29.344599f
C15 minus plus 9.262711f
C16 minus commonsourceibias 0.323289f
C17 plus commonsourceibias 0.277692f
C18 diffpairibias gnd 48.96854f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.119336p
C22 plus gnd 32.908802f
C23 minus gnd 27.27192f
C24 CSoutput gnd 89.10971f
C25 vdd gnd 0.543041p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 outputibias.t8 gnd 0.11477f
C74 outputibias.t10 gnd 0.115567f
C75 outputibias.n0 gnd 0.130108f
C76 outputibias.n1 gnd 0.001372f
C77 outputibias.n2 gnd 9.76e-19
C78 outputibias.n3 gnd 5.24e-19
C79 outputibias.n4 gnd 0.001239f
C80 outputibias.n5 gnd 5.55e-19
C81 outputibias.n6 gnd 9.76e-19
C82 outputibias.n7 gnd 5.24e-19
C83 outputibias.n8 gnd 0.001239f
C84 outputibias.n9 gnd 5.55e-19
C85 outputibias.n10 gnd 0.004176f
C86 outputibias.t7 gnd 0.00202f
C87 outputibias.n11 gnd 9.3e-19
C88 outputibias.n12 gnd 7.32e-19
C89 outputibias.n13 gnd 5.24e-19
C90 outputibias.n14 gnd 0.02322f
C91 outputibias.n15 gnd 9.76e-19
C92 outputibias.n16 gnd 5.24e-19
C93 outputibias.n17 gnd 5.55e-19
C94 outputibias.n18 gnd 0.001239f
C95 outputibias.n19 gnd 0.001239f
C96 outputibias.n20 gnd 5.55e-19
C97 outputibias.n21 gnd 5.24e-19
C98 outputibias.n22 gnd 9.76e-19
C99 outputibias.n23 gnd 9.76e-19
C100 outputibias.n24 gnd 5.24e-19
C101 outputibias.n25 gnd 5.55e-19
C102 outputibias.n26 gnd 0.001239f
C103 outputibias.n27 gnd 0.002683f
C104 outputibias.n28 gnd 5.55e-19
C105 outputibias.n29 gnd 5.24e-19
C106 outputibias.n30 gnd 0.002256f
C107 outputibias.n31 gnd 0.005781f
C108 outputibias.n32 gnd 0.001372f
C109 outputibias.n33 gnd 9.76e-19
C110 outputibias.n34 gnd 5.24e-19
C111 outputibias.n35 gnd 0.001239f
C112 outputibias.n36 gnd 5.55e-19
C113 outputibias.n37 gnd 9.76e-19
C114 outputibias.n38 gnd 5.24e-19
C115 outputibias.n39 gnd 0.001239f
C116 outputibias.n40 gnd 5.55e-19
C117 outputibias.n41 gnd 0.004176f
C118 outputibias.t1 gnd 0.00202f
C119 outputibias.n42 gnd 9.3e-19
C120 outputibias.n43 gnd 7.32e-19
C121 outputibias.n44 gnd 5.24e-19
C122 outputibias.n45 gnd 0.02322f
C123 outputibias.n46 gnd 9.76e-19
C124 outputibias.n47 gnd 5.24e-19
C125 outputibias.n48 gnd 5.55e-19
C126 outputibias.n49 gnd 0.001239f
C127 outputibias.n50 gnd 0.001239f
C128 outputibias.n51 gnd 5.55e-19
C129 outputibias.n52 gnd 5.24e-19
C130 outputibias.n53 gnd 9.76e-19
C131 outputibias.n54 gnd 9.76e-19
C132 outputibias.n55 gnd 5.24e-19
C133 outputibias.n56 gnd 5.55e-19
C134 outputibias.n57 gnd 0.001239f
C135 outputibias.n58 gnd 0.002683f
C136 outputibias.n59 gnd 5.55e-19
C137 outputibias.n60 gnd 5.24e-19
C138 outputibias.n61 gnd 0.002256f
C139 outputibias.n62 gnd 0.005197f
C140 outputibias.n63 gnd 0.121892f
C141 outputibias.n64 gnd 0.001372f
C142 outputibias.n65 gnd 9.76e-19
C143 outputibias.n66 gnd 5.24e-19
C144 outputibias.n67 gnd 0.001239f
C145 outputibias.n68 gnd 5.55e-19
C146 outputibias.n69 gnd 9.76e-19
C147 outputibias.n70 gnd 5.24e-19
C148 outputibias.n71 gnd 0.001239f
C149 outputibias.n72 gnd 5.55e-19
C150 outputibias.n73 gnd 0.004176f
C151 outputibias.t5 gnd 0.00202f
C152 outputibias.n74 gnd 9.3e-19
C153 outputibias.n75 gnd 7.32e-19
C154 outputibias.n76 gnd 5.24e-19
C155 outputibias.n77 gnd 0.02322f
C156 outputibias.n78 gnd 9.76e-19
C157 outputibias.n79 gnd 5.24e-19
C158 outputibias.n80 gnd 5.55e-19
C159 outputibias.n81 gnd 0.001239f
C160 outputibias.n82 gnd 0.001239f
C161 outputibias.n83 gnd 5.55e-19
C162 outputibias.n84 gnd 5.24e-19
C163 outputibias.n85 gnd 9.76e-19
C164 outputibias.n86 gnd 9.76e-19
C165 outputibias.n87 gnd 5.24e-19
C166 outputibias.n88 gnd 5.55e-19
C167 outputibias.n89 gnd 0.001239f
C168 outputibias.n90 gnd 0.002683f
C169 outputibias.n91 gnd 5.55e-19
C170 outputibias.n92 gnd 5.24e-19
C171 outputibias.n93 gnd 0.002256f
C172 outputibias.n94 gnd 0.005197f
C173 outputibias.n95 gnd 0.064513f
C174 outputibias.n96 gnd 0.001372f
C175 outputibias.n97 gnd 9.76e-19
C176 outputibias.n98 gnd 5.24e-19
C177 outputibias.n99 gnd 0.001239f
C178 outputibias.n100 gnd 5.55e-19
C179 outputibias.n101 gnd 9.76e-19
C180 outputibias.n102 gnd 5.24e-19
C181 outputibias.n103 gnd 0.001239f
C182 outputibias.n104 gnd 5.55e-19
C183 outputibias.n105 gnd 0.004176f
C184 outputibias.t3 gnd 0.00202f
C185 outputibias.n106 gnd 9.3e-19
C186 outputibias.n107 gnd 7.32e-19
C187 outputibias.n108 gnd 5.24e-19
C188 outputibias.n109 gnd 0.02322f
C189 outputibias.n110 gnd 9.76e-19
C190 outputibias.n111 gnd 5.24e-19
C191 outputibias.n112 gnd 5.55e-19
C192 outputibias.n113 gnd 0.001239f
C193 outputibias.n114 gnd 0.001239f
C194 outputibias.n115 gnd 5.55e-19
C195 outputibias.n116 gnd 5.24e-19
C196 outputibias.n117 gnd 9.76e-19
C197 outputibias.n118 gnd 9.76e-19
C198 outputibias.n119 gnd 5.24e-19
C199 outputibias.n120 gnd 5.55e-19
C200 outputibias.n121 gnd 0.001239f
C201 outputibias.n122 gnd 0.002683f
C202 outputibias.n123 gnd 5.55e-19
C203 outputibias.n124 gnd 5.24e-19
C204 outputibias.n125 gnd 0.002256f
C205 outputibias.n126 gnd 0.005197f
C206 outputibias.n127 gnd 0.084814f
C207 outputibias.t2 gnd 0.108319f
C208 outputibias.t4 gnd 0.108319f
C209 outputibias.t0 gnd 0.108319f
C210 outputibias.t6 gnd 0.109238f
C211 outputibias.n128 gnd 0.134674f
C212 outputibias.n129 gnd 0.07244f
C213 outputibias.n130 gnd 0.079818f
C214 outputibias.n131 gnd 0.164901f
C215 outputibias.t11 gnd 0.11477f
C216 outputibias.n132 gnd 0.067481f
C217 outputibias.t9 gnd 0.11477f
C218 outputibias.n133 gnd 0.065115f
C219 outputibias.n134 gnd 0.029159f
C220 a_n2982_8322.t13 gnd 0.100161f
C221 a_n2982_8322.t2 gnd 20.7793f
C222 a_n2982_8322.t1 gnd 20.633598f
C223 a_n2982_8322.t5 gnd 20.633598f
C224 a_n2982_8322.t4 gnd 20.7793f
C225 a_n2982_8322.t3 gnd 20.633598f
C226 a_n2982_8322.t0 gnd 28.9697f
C227 a_n2982_8322.t12 gnd 0.937857f
C228 a_n2982_8322.t25 gnd 0.100161f
C229 a_n2982_8322.t21 gnd 0.100161f
C230 a_n2982_8322.n0 gnd 0.705534f
C231 a_n2982_8322.n1 gnd 0.78833f
C232 a_n2982_8322.t28 gnd 0.100161f
C233 a_n2982_8322.t18 gnd 0.100161f
C234 a_n2982_8322.n2 gnd 0.705534f
C235 a_n2982_8322.n3 gnd 0.40054f
C236 a_n2982_8322.t9 gnd 0.100161f
C237 a_n2982_8322.t8 gnd 0.100161f
C238 a_n2982_8322.n4 gnd 0.705534f
C239 a_n2982_8322.n5 gnd 0.40054f
C240 a_n2982_8322.t22 gnd 0.100161f
C241 a_n2982_8322.t15 gnd 0.100161f
C242 a_n2982_8322.n6 gnd 0.705534f
C243 a_n2982_8322.n7 gnd 0.40054f
C244 a_n2982_8322.t19 gnd 0.100161f
C245 a_n2982_8322.t17 gnd 0.100161f
C246 a_n2982_8322.n8 gnd 0.705534f
C247 a_n2982_8322.n9 gnd 0.40054f
C248 a_n2982_8322.t6 gnd 0.935989f
C249 a_n2982_8322.n10 gnd 1.87142f
C250 a_n2982_8322.t33 gnd 0.937857f
C251 a_n2982_8322.t37 gnd 0.100161f
C252 a_n2982_8322.t36 gnd 0.100161f
C253 a_n2982_8322.n11 gnd 0.705534f
C254 a_n2982_8322.n12 gnd 0.78833f
C255 a_n2982_8322.t31 gnd 0.935989f
C256 a_n2982_8322.n13 gnd 0.396699f
C257 a_n2982_8322.t34 gnd 0.935989f
C258 a_n2982_8322.n14 gnd 0.396699f
C259 a_n2982_8322.t32 gnd 0.100161f
C260 a_n2982_8322.t30 gnd 0.100161f
C261 a_n2982_8322.n15 gnd 0.705534f
C262 a_n2982_8322.n16 gnd 0.40054f
C263 a_n2982_8322.t35 gnd 0.935989f
C264 a_n2982_8322.n17 gnd 1.47142f
C265 a_n2982_8322.n18 gnd 2.35138f
C266 a_n2982_8322.n19 gnd 3.33814f
C267 a_n2982_8322.t7 gnd 0.935989f
C268 a_n2982_8322.n20 gnd 1.11148f
C269 a_n2982_8322.t24 gnd 0.100161f
C270 a_n2982_8322.t23 gnd 0.100161f
C271 a_n2982_8322.n21 gnd 0.705534f
C272 a_n2982_8322.n22 gnd 0.40054f
C273 a_n2982_8322.t11 gnd 0.100161f
C274 a_n2982_8322.t10 gnd 0.100161f
C275 a_n2982_8322.n23 gnd 0.705534f
C276 a_n2982_8322.n24 gnd 0.40054f
C277 a_n2982_8322.t26 gnd 0.100161f
C278 a_n2982_8322.t14 gnd 0.100161f
C279 a_n2982_8322.n25 gnd 0.705534f
C280 a_n2982_8322.n26 gnd 0.40054f
C281 a_n2982_8322.t27 gnd 0.937854f
C282 a_n2982_8322.t20 gnd 0.100161f
C283 a_n2982_8322.t16 gnd 0.100161f
C284 a_n2982_8322.n27 gnd 0.705534f
C285 a_n2982_8322.n28 gnd 0.788332f
C286 a_n2982_8322.n29 gnd 0.400539f
C287 a_n2982_8322.n30 gnd 0.705536f
C288 a_n2982_8322.t29 gnd 0.100161f
C289 minus.n0 gnd 0.029852f
C290 minus.t14 gnd 0.501953f
C291 minus.n1 gnd 0.203012f
C292 minus.n2 gnd 0.029852f
C293 minus.t19 gnd 0.501953f
C294 minus.n3 gnd 0.024263f
C295 minus.n4 gnd 0.029852f
C296 minus.t18 gnd 0.501953f
C297 minus.t5 gnd 0.501953f
C298 minus.n5 gnd 0.203012f
C299 minus.n6 gnd 0.029852f
C300 minus.t8 gnd 0.501953f
C301 minus.n7 gnd 0.203012f
C302 minus.n8 gnd 0.128142f
C303 minus.t9 gnd 0.501953f
C304 minus.t13 gnd 0.563561f
C305 minus.n9 gnd 0.23555f
C306 minus.n10 gnd 0.234447f
C307 minus.n11 gnd 0.037133f
C308 minus.n12 gnd 0.034898f
C309 minus.n13 gnd 0.029852f
C310 minus.n14 gnd 0.029852f
C311 minus.n15 gnd 0.037394f
C312 minus.n16 gnd 0.024263f
C313 minus.n17 gnd 0.038403f
C314 minus.n18 gnd 0.029852f
C315 minus.n19 gnd 0.029852f
C316 minus.n20 gnd 0.036016f
C317 minus.n21 gnd 0.036016f
C318 minus.n22 gnd 0.203012f
C319 minus.n23 gnd 0.038403f
C320 minus.n24 gnd 0.029852f
C321 minus.n25 gnd 0.029852f
C322 minus.n26 gnd 0.029852f
C323 minus.n27 gnd 0.037394f
C324 minus.n28 gnd 0.203012f
C325 minus.n29 gnd 0.034898f
C326 minus.n30 gnd 0.037133f
C327 minus.n31 gnd 0.029852f
C328 minus.n32 gnd 0.029852f
C329 minus.n33 gnd 0.038878f
C330 minus.n34 gnd 0.012364f
C331 minus.t17 gnd 0.542863f
C332 minus.n35 gnd 0.23579f
C333 minus.n36 gnd 0.350764f
C334 minus.n37 gnd 0.029852f
C335 minus.t15 gnd 0.542863f
C336 minus.t12 gnd 0.501953f
C337 minus.n38 gnd 0.203012f
C338 minus.n39 gnd 0.029852f
C339 minus.t7 gnd 0.501953f
C340 minus.n40 gnd 0.024263f
C341 minus.n41 gnd 0.029852f
C342 minus.t6 gnd 0.501953f
C343 minus.t11 gnd 0.501953f
C344 minus.n42 gnd 0.203012f
C345 minus.n43 gnd 0.029852f
C346 minus.t10 gnd 0.501953f
C347 minus.n44 gnd 0.203012f
C348 minus.n45 gnd 0.128142f
C349 minus.t16 gnd 0.501953f
C350 minus.t20 gnd 0.563561f
C351 minus.n46 gnd 0.23555f
C352 minus.n47 gnd 0.234447f
C353 minus.n48 gnd 0.037133f
C354 minus.n49 gnd 0.034898f
C355 minus.n50 gnd 0.029852f
C356 minus.n51 gnd 0.029852f
C357 minus.n52 gnd 0.037394f
C358 minus.n53 gnd 0.024263f
C359 minus.n54 gnd 0.038403f
C360 minus.n55 gnd 0.029852f
C361 minus.n56 gnd 0.029852f
C362 minus.n57 gnd 0.036016f
C363 minus.n58 gnd 0.036016f
C364 minus.n59 gnd 0.203012f
C365 minus.n60 gnd 0.038403f
C366 minus.n61 gnd 0.029852f
C367 minus.n62 gnd 0.029852f
C368 minus.n63 gnd 0.029852f
C369 minus.n64 gnd 0.037394f
C370 minus.n65 gnd 0.203012f
C371 minus.n66 gnd 0.034898f
C372 minus.n67 gnd 0.037133f
C373 minus.n68 gnd 0.029852f
C374 minus.n69 gnd 0.029852f
C375 minus.n70 gnd 0.038878f
C376 minus.n71 gnd 0.012364f
C377 minus.n72 gnd 0.23579f
C378 minus.n73 gnd 0.930168f
C379 minus.n74 gnd 1.39812f
C380 minus.t1 gnd 0.009202f
C381 minus.t4 gnd 0.009202f
C382 minus.n75 gnd 0.03026f
C383 minus.t2 gnd 0.009202f
C384 minus.t0 gnd 0.009202f
C385 minus.n76 gnd 0.029845f
C386 minus.n77 gnd 0.254715f
C387 minus.t3 gnd 0.05122f
C388 minus.n78 gnd 0.138995f
C389 minus.n79 gnd 1.93735f
C390 a_n2903_n3924.n0 gnd 1.45586f
C391 a_n2903_n3924.t5 gnd 0.088483f
C392 a_n2903_n3924.t14 gnd 0.919619f
C393 a_n2903_n3924.n1 gnd 0.347657f
C394 a_n2903_n3924.t31 gnd 1.14306f
C395 a_n2903_n3924.n2 gnd 1.19083f
C396 a_n2903_n3924.t22 gnd 0.919619f
C397 a_n2903_n3924.n3 gnd 0.347657f
C398 a_n2903_n3924.t24 gnd 0.088483f
C399 a_n2903_n3924.t19 gnd 0.088483f
C400 a_n2903_n3924.n4 gnd 0.722655f
C401 a_n2903_n3924.n5 gnd 0.364177f
C402 a_n2903_n3924.t30 gnd 0.088483f
C403 a_n2903_n3924.t32 gnd 0.088483f
C404 a_n2903_n3924.n6 gnd 0.722655f
C405 a_n2903_n3924.n7 gnd 0.364177f
C406 a_n2903_n3924.t1 gnd 0.088483f
C407 a_n2903_n3924.t29 gnd 0.088483f
C408 a_n2903_n3924.n8 gnd 0.722655f
C409 a_n2903_n3924.n9 gnd 0.364177f
C410 a_n2903_n3924.t0 gnd 0.919619f
C411 a_n2903_n3924.n10 gnd 0.860834f
C412 a_n2903_n3924.t35 gnd 1.14419f
C413 a_n2903_n3924.t36 gnd 1.14261f
C414 a_n2903_n3924.n11 gnd 0.745791f
C415 a_n2903_n3924.t39 gnd 1.14261f
C416 a_n2903_n3924.n12 gnd 0.804756f
C417 a_n2903_n3924.t38 gnd 1.14261f
C418 a_n2903_n3924.n13 gnd 0.804756f
C419 a_n2903_n3924.t27 gnd 1.14261f
C420 a_n2903_n3924.n14 gnd 0.804756f
C421 a_n2903_n3924.t21 gnd 1.14261f
C422 a_n2903_n3924.n15 gnd 0.804756f
C423 a_n2903_n3924.t20 gnd 1.14261f
C424 a_n2903_n3924.n16 gnd 0.834168f
C425 a_n2903_n3924.t16 gnd 0.919616f
C426 a_n2903_n3924.n17 gnd 0.571219f
C427 a_n2903_n3924.t17 gnd 0.088483f
C428 a_n2903_n3924.t7 gnd 0.088483f
C429 a_n2903_n3924.n18 gnd 0.722654f
C430 a_n2903_n3924.n19 gnd 0.364178f
C431 a_n2903_n3924.t8 gnd 0.088483f
C432 a_n2903_n3924.t3 gnd 0.088483f
C433 a_n2903_n3924.n20 gnd 0.722654f
C434 a_n2903_n3924.n21 gnd 0.364178f
C435 a_n2903_n3924.t4 gnd 0.088483f
C436 a_n2903_n3924.t15 gnd 0.088483f
C437 a_n2903_n3924.n22 gnd 0.722654f
C438 a_n2903_n3924.n23 gnd 0.364178f
C439 a_n2903_n3924.t12 gnd 0.919616f
C440 a_n2903_n3924.n24 gnd 0.347661f
C441 a_n2903_n3924.t2 gnd 0.919616f
C442 a_n2903_n3924.n25 gnd 0.347661f
C443 a_n2903_n3924.t26 gnd 0.088483f
C444 a_n2903_n3924.t23 gnd 0.088483f
C445 a_n2903_n3924.n26 gnd 0.722654f
C446 a_n2903_n3924.n27 gnd 0.364178f
C447 a_n2903_n3924.t25 gnd 0.088483f
C448 a_n2903_n3924.t33 gnd 0.088483f
C449 a_n2903_n3924.n28 gnd 0.722654f
C450 a_n2903_n3924.n29 gnd 0.364178f
C451 a_n2903_n3924.t34 gnd 0.088483f
C452 a_n2903_n3924.t28 gnd 0.088483f
C453 a_n2903_n3924.n30 gnd 0.722654f
C454 a_n2903_n3924.n31 gnd 0.364178f
C455 a_n2903_n3924.t37 gnd 0.919616f
C456 a_n2903_n3924.n32 gnd 0.571219f
C457 a_n2903_n3924.n33 gnd 0.834168f
C458 a_n2903_n3924.t11 gnd 0.919616f
C459 a_n2903_n3924.n34 gnd 0.860837f
C460 a_n2903_n3924.t9 gnd 0.088483f
C461 a_n2903_n3924.t13 gnd 0.088483f
C462 a_n2903_n3924.n35 gnd 0.722655f
C463 a_n2903_n3924.n36 gnd 0.364177f
C464 a_n2903_n3924.t6 gnd 0.088483f
C465 a_n2903_n3924.t10 gnd 0.088483f
C466 a_n2903_n3924.n37 gnd 0.722655f
C467 a_n2903_n3924.n38 gnd 0.364177f
C468 a_n2903_n3924.n39 gnd 0.364176f
C469 a_n2903_n3924.n40 gnd 0.722656f
C470 a_n2903_n3924.t18 gnd 0.088483f
C471 plus.n0 gnd 0.021954f
C472 plus.t7 gnd 0.399245f
C473 plus.t6 gnd 0.369159f
C474 plus.n1 gnd 0.149304f
C475 plus.n2 gnd 0.021954f
C476 plus.t16 gnd 0.369159f
C477 plus.n3 gnd 0.017844f
C478 plus.n4 gnd 0.021954f
C479 plus.t15 gnd 0.369159f
C480 plus.t20 gnd 0.369159f
C481 plus.n5 gnd 0.149304f
C482 plus.n6 gnd 0.021954f
C483 plus.t19 gnd 0.369159f
C484 plus.n7 gnd 0.149304f
C485 plus.n8 gnd 0.094241f
C486 plus.t8 gnd 0.369159f
C487 plus.t11 gnd 0.414468f
C488 plus.n9 gnd 0.173234f
C489 plus.n10 gnd 0.172423f
C490 plus.n11 gnd 0.027309f
C491 plus.n12 gnd 0.025666f
C492 plus.n13 gnd 0.021954f
C493 plus.n14 gnd 0.021954f
C494 plus.n15 gnd 0.027501f
C495 plus.n16 gnd 0.017844f
C496 plus.n17 gnd 0.028243f
C497 plus.n18 gnd 0.021954f
C498 plus.n19 gnd 0.021954f
C499 plus.n20 gnd 0.026487f
C500 plus.n21 gnd 0.026487f
C501 plus.n22 gnd 0.149304f
C502 plus.n23 gnd 0.028243f
C503 plus.n24 gnd 0.021954f
C504 plus.n25 gnd 0.021954f
C505 plus.n26 gnd 0.021954f
C506 plus.n27 gnd 0.027501f
C507 plus.n28 gnd 0.149304f
C508 plus.n29 gnd 0.025666f
C509 plus.n30 gnd 0.027309f
C510 plus.n31 gnd 0.021954f
C511 plus.n32 gnd 0.021954f
C512 plus.n33 gnd 0.028593f
C513 plus.n34 gnd 0.009093f
C514 plus.n35 gnd 0.17341f
C515 plus.n36 gnd 0.252321f
C516 plus.n37 gnd 0.021954f
C517 plus.t10 gnd 0.369159f
C518 plus.n38 gnd 0.149304f
C519 plus.n39 gnd 0.021954f
C520 plus.t14 gnd 0.369159f
C521 plus.n40 gnd 0.017844f
C522 plus.n41 gnd 0.021954f
C523 plus.t13 gnd 0.369159f
C524 plus.t17 gnd 0.369159f
C525 plus.n42 gnd 0.149304f
C526 plus.n43 gnd 0.021954f
C527 plus.t18 gnd 0.369159f
C528 plus.n44 gnd 0.149304f
C529 plus.n45 gnd 0.094241f
C530 plus.t5 gnd 0.369159f
C531 plus.t9 gnd 0.414468f
C532 plus.n46 gnd 0.173234f
C533 plus.n47 gnd 0.172423f
C534 plus.n48 gnd 0.027309f
C535 plus.n49 gnd 0.025666f
C536 plus.n50 gnd 0.021954f
C537 plus.n51 gnd 0.021954f
C538 plus.n52 gnd 0.027501f
C539 plus.n53 gnd 0.017844f
C540 plus.n54 gnd 0.028243f
C541 plus.n55 gnd 0.021954f
C542 plus.n56 gnd 0.021954f
C543 plus.n57 gnd 0.026487f
C544 plus.n58 gnd 0.026487f
C545 plus.n59 gnd 0.149304f
C546 plus.n60 gnd 0.028243f
C547 plus.n61 gnd 0.021954f
C548 plus.n62 gnd 0.021954f
C549 plus.n63 gnd 0.021954f
C550 plus.n64 gnd 0.027501f
C551 plus.n65 gnd 0.149304f
C552 plus.n66 gnd 0.025666f
C553 plus.n67 gnd 0.027309f
C554 plus.n68 gnd 0.021954f
C555 plus.n69 gnd 0.021954f
C556 plus.n70 gnd 0.028593f
C557 plus.n71 gnd 0.009093f
C558 plus.t12 gnd 0.399245f
C559 plus.n72 gnd 0.17341f
C560 plus.n73 gnd 0.67529f
C561 plus.n74 gnd 1.01953f
C562 plus.t4 gnd 0.0379f
C563 plus.t1 gnd 0.006768f
C564 plus.t2 gnd 0.006768f
C565 plus.n75 gnd 0.021949f
C566 plus.n76 gnd 0.170395f
C567 plus.t0 gnd 0.006768f
C568 plus.t3 gnd 0.006768f
C569 plus.n77 gnd 0.021949f
C570 plus.n78 gnd 0.127902f
C571 plus.n79 gnd 2.52333f
C572 output.t9 gnd 0.464308f
C573 output.t5 gnd 0.044422f
C574 output.t3 gnd 0.044422f
C575 output.n0 gnd 0.364624f
C576 output.n1 gnd 0.614102f
C577 output.t13 gnd 0.044422f
C578 output.t15 gnd 0.044422f
C579 output.n2 gnd 0.364624f
C580 output.n3 gnd 0.350265f
C581 output.t16 gnd 0.044422f
C582 output.t7 gnd 0.044422f
C583 output.n4 gnd 0.364624f
C584 output.n5 gnd 0.350265f
C585 output.t10 gnd 0.044422f
C586 output.t14 gnd 0.044422f
C587 output.n6 gnd 0.364624f
C588 output.n7 gnd 0.350265f
C589 output.t1 gnd 0.044422f
C590 output.t6 gnd 0.044422f
C591 output.n8 gnd 0.364624f
C592 output.n9 gnd 0.350265f
C593 output.t8 gnd 0.044422f
C594 output.t12 gnd 0.044422f
C595 output.n10 gnd 0.364624f
C596 output.n11 gnd 0.350265f
C597 output.t4 gnd 0.044422f
C598 output.t2 gnd 0.044422f
C599 output.n12 gnd 0.364624f
C600 output.n13 gnd 0.350265f
C601 output.t11 gnd 0.462979f
C602 output.n14 gnd 0.28994f
C603 output.n15 gnd 0.015803f
C604 output.n16 gnd 0.011243f
C605 output.n17 gnd 0.006041f
C606 output.n18 gnd 0.01428f
C607 output.n19 gnd 0.006397f
C608 output.n20 gnd 0.011243f
C609 output.n21 gnd 0.006041f
C610 output.n22 gnd 0.01428f
C611 output.n23 gnd 0.006397f
C612 output.n24 gnd 0.048111f
C613 output.t19 gnd 0.023274f
C614 output.n25 gnd 0.01071f
C615 output.n26 gnd 0.008435f
C616 output.n27 gnd 0.006041f
C617 output.n28 gnd 0.267512f
C618 output.n29 gnd 0.011243f
C619 output.n30 gnd 0.006041f
C620 output.n31 gnd 0.006397f
C621 output.n32 gnd 0.01428f
C622 output.n33 gnd 0.01428f
C623 output.n34 gnd 0.006397f
C624 output.n35 gnd 0.006041f
C625 output.n36 gnd 0.011243f
C626 output.n37 gnd 0.011243f
C627 output.n38 gnd 0.006041f
C628 output.n39 gnd 0.006397f
C629 output.n40 gnd 0.01428f
C630 output.n41 gnd 0.030913f
C631 output.n42 gnd 0.006397f
C632 output.n43 gnd 0.006041f
C633 output.n44 gnd 0.025987f
C634 output.n45 gnd 0.097665f
C635 output.n46 gnd 0.015803f
C636 output.n47 gnd 0.011243f
C637 output.n48 gnd 0.006041f
C638 output.n49 gnd 0.01428f
C639 output.n50 gnd 0.006397f
C640 output.n51 gnd 0.011243f
C641 output.n52 gnd 0.006041f
C642 output.n53 gnd 0.01428f
C643 output.n54 gnd 0.006397f
C644 output.n55 gnd 0.048111f
C645 output.t0 gnd 0.023274f
C646 output.n56 gnd 0.01071f
C647 output.n57 gnd 0.008435f
C648 output.n58 gnd 0.006041f
C649 output.n59 gnd 0.267512f
C650 output.n60 gnd 0.011243f
C651 output.n61 gnd 0.006041f
C652 output.n62 gnd 0.006397f
C653 output.n63 gnd 0.01428f
C654 output.n64 gnd 0.01428f
C655 output.n65 gnd 0.006397f
C656 output.n66 gnd 0.006041f
C657 output.n67 gnd 0.011243f
C658 output.n68 gnd 0.011243f
C659 output.n69 gnd 0.006041f
C660 output.n70 gnd 0.006397f
C661 output.n71 gnd 0.01428f
C662 output.n72 gnd 0.030913f
C663 output.n73 gnd 0.006397f
C664 output.n74 gnd 0.006041f
C665 output.n75 gnd 0.025987f
C666 output.n76 gnd 0.09306f
C667 output.n77 gnd 1.65264f
C668 output.n78 gnd 0.015803f
C669 output.n79 gnd 0.011243f
C670 output.n80 gnd 0.006041f
C671 output.n81 gnd 0.01428f
C672 output.n82 gnd 0.006397f
C673 output.n83 gnd 0.011243f
C674 output.n84 gnd 0.006041f
C675 output.n85 gnd 0.01428f
C676 output.n86 gnd 0.006397f
C677 output.n87 gnd 0.048111f
C678 output.t17 gnd 0.023274f
C679 output.n88 gnd 0.01071f
C680 output.n89 gnd 0.008435f
C681 output.n90 gnd 0.006041f
C682 output.n91 gnd 0.267512f
C683 output.n92 gnd 0.011243f
C684 output.n93 gnd 0.006041f
C685 output.n94 gnd 0.006397f
C686 output.n95 gnd 0.01428f
C687 output.n96 gnd 0.01428f
C688 output.n97 gnd 0.006397f
C689 output.n98 gnd 0.006041f
C690 output.n99 gnd 0.011243f
C691 output.n100 gnd 0.011243f
C692 output.n101 gnd 0.006041f
C693 output.n102 gnd 0.006397f
C694 output.n103 gnd 0.01428f
C695 output.n104 gnd 0.030913f
C696 output.n105 gnd 0.006397f
C697 output.n106 gnd 0.006041f
C698 output.n107 gnd 0.025987f
C699 output.n108 gnd 0.09306f
C700 output.n109 gnd 0.713089f
C701 output.n110 gnd 0.015803f
C702 output.n111 gnd 0.011243f
C703 output.n112 gnd 0.006041f
C704 output.n113 gnd 0.01428f
C705 output.n114 gnd 0.006397f
C706 output.n115 gnd 0.011243f
C707 output.n116 gnd 0.006041f
C708 output.n117 gnd 0.01428f
C709 output.n118 gnd 0.006397f
C710 output.n119 gnd 0.048111f
C711 output.t18 gnd 0.023274f
C712 output.n120 gnd 0.01071f
C713 output.n121 gnd 0.008435f
C714 output.n122 gnd 0.006041f
C715 output.n123 gnd 0.267512f
C716 output.n124 gnd 0.011243f
C717 output.n125 gnd 0.006041f
C718 output.n126 gnd 0.006397f
C719 output.n127 gnd 0.01428f
C720 output.n128 gnd 0.01428f
C721 output.n129 gnd 0.006397f
C722 output.n130 gnd 0.006041f
C723 output.n131 gnd 0.011243f
C724 output.n132 gnd 0.011243f
C725 output.n133 gnd 0.006041f
C726 output.n134 gnd 0.006397f
C727 output.n135 gnd 0.01428f
C728 output.n136 gnd 0.030913f
C729 output.n137 gnd 0.006397f
C730 output.n138 gnd 0.006041f
C731 output.n139 gnd 0.025987f
C732 output.n140 gnd 0.09306f
C733 output.n141 gnd 1.67353f
C734 a_n9628_8799.n0 gnd 2.75765f
C735 a_n9628_8799.n1 gnd 1.67079f
C736 a_n9628_8799.n2 gnd 3.82259f
C737 a_n9628_8799.n3 gnd 0.208483f
C738 a_n9628_8799.n4 gnd 0.286275f
C739 a_n9628_8799.n5 gnd 0.208483f
C740 a_n9628_8799.n6 gnd 0.208483f
C741 a_n9628_8799.n7 gnd 0.208483f
C742 a_n9628_8799.n8 gnd 0.208483f
C743 a_n9628_8799.n9 gnd 0.208483f
C744 a_n9628_8799.n10 gnd 0.216785f
C745 a_n9628_8799.n11 gnd 0.208483f
C746 a_n9628_8799.n12 gnd 0.286275f
C747 a_n9628_8799.n13 gnd 0.208483f
C748 a_n9628_8799.n14 gnd 0.208483f
C749 a_n9628_8799.n15 gnd 0.208483f
C750 a_n9628_8799.n16 gnd 0.208483f
C751 a_n9628_8799.n17 gnd 0.208483f
C752 a_n9628_8799.n18 gnd 0.216785f
C753 a_n9628_8799.n19 gnd 0.208483f
C754 a_n9628_8799.n20 gnd 0.451874f
C755 a_n9628_8799.n21 gnd 0.208483f
C756 a_n9628_8799.n22 gnd 0.208483f
C757 a_n9628_8799.n23 gnd 0.208483f
C758 a_n9628_8799.n24 gnd 0.208483f
C759 a_n9628_8799.n25 gnd 0.208483f
C760 a_n9628_8799.n26 gnd 0.216785f
C761 a_n9628_8799.n27 gnd 0.208483f
C762 a_n9628_8799.n28 gnd 0.321027f
C763 a_n9628_8799.n29 gnd 0.208483f
C764 a_n9628_8799.n30 gnd 0.208483f
C765 a_n9628_8799.n31 gnd 0.208483f
C766 a_n9628_8799.n32 gnd 0.208483f
C767 a_n9628_8799.n33 gnd 0.208483f
C768 a_n9628_8799.n34 gnd 0.182033f
C769 a_n9628_8799.n35 gnd 0.208483f
C770 a_n9628_8799.n36 gnd 0.321027f
C771 a_n9628_8799.n37 gnd 0.208483f
C772 a_n9628_8799.n38 gnd 0.208483f
C773 a_n9628_8799.n39 gnd 0.208483f
C774 a_n9628_8799.n40 gnd 0.208483f
C775 a_n9628_8799.n41 gnd 0.208483f
C776 a_n9628_8799.n42 gnd 0.182033f
C777 a_n9628_8799.n43 gnd 0.208483f
C778 a_n9628_8799.n44 gnd 0.321027f
C779 a_n9628_8799.n45 gnd 0.208483f
C780 a_n9628_8799.n46 gnd 0.208483f
C781 a_n9628_8799.n47 gnd 0.208483f
C782 a_n9628_8799.n48 gnd 0.208483f
C783 a_n9628_8799.n49 gnd 0.208483f
C784 a_n9628_8799.n50 gnd 0.347632f
C785 a_n9628_8799.n51 gnd 1.02351f
C786 a_n9628_8799.n52 gnd 1.00901f
C787 a_n9628_8799.n53 gnd 3.02795f
C788 a_n9628_8799.n54 gnd 1.52802f
C789 a_n9628_8799.n55 gnd 1.00901f
C790 a_n9628_8799.n56 gnd 0.250994f
C791 a_n9628_8799.n57 gnd 0.003669f
C792 a_n9628_8799.n58 gnd 0.009673f
C793 a_n9628_8799.n59 gnd 0.010568f
C794 a_n9628_8799.n60 gnd 0.005584f
C795 a_n9628_8799.n62 gnd 0.004686f
C796 a_n9628_8799.n63 gnd 0.010134f
C797 a_n9628_8799.n64 gnd 0.010134f
C798 a_n9628_8799.n65 gnd 0.004686f
C799 a_n9628_8799.n67 gnd 0.005584f
C800 a_n9628_8799.n68 gnd 0.010568f
C801 a_n9628_8799.n69 gnd 0.009673f
C802 a_n9628_8799.n70 gnd 0.003669f
C803 a_n9628_8799.n71 gnd 0.250994f
C804 a_n9628_8799.n72 gnd 0.003669f
C805 a_n9628_8799.n73 gnd 0.009673f
C806 a_n9628_8799.n74 gnd 0.010568f
C807 a_n9628_8799.n75 gnd 0.005584f
C808 a_n9628_8799.n77 gnd 0.004686f
C809 a_n9628_8799.n78 gnd 0.010134f
C810 a_n9628_8799.n79 gnd 0.010134f
C811 a_n9628_8799.n80 gnd 0.004686f
C812 a_n9628_8799.n82 gnd 0.005584f
C813 a_n9628_8799.n83 gnd 0.010568f
C814 a_n9628_8799.n84 gnd 0.009673f
C815 a_n9628_8799.n85 gnd 0.003669f
C816 a_n9628_8799.n86 gnd 0.250994f
C817 a_n9628_8799.n87 gnd 0.003669f
C818 a_n9628_8799.n88 gnd 0.009673f
C819 a_n9628_8799.n89 gnd 0.010568f
C820 a_n9628_8799.n90 gnd 0.005584f
C821 a_n9628_8799.n92 gnd 0.004686f
C822 a_n9628_8799.n93 gnd 0.010134f
C823 a_n9628_8799.n94 gnd 0.010134f
C824 a_n9628_8799.n95 gnd 0.004686f
C825 a_n9628_8799.n97 gnd 0.005584f
C826 a_n9628_8799.n98 gnd 0.010568f
C827 a_n9628_8799.n99 gnd 0.009673f
C828 a_n9628_8799.n100 gnd 0.003669f
C829 a_n9628_8799.n101 gnd 0.003669f
C830 a_n9628_8799.n102 gnd 0.009673f
C831 a_n9628_8799.n103 gnd 0.010568f
C832 a_n9628_8799.n104 gnd 0.005584f
C833 a_n9628_8799.n106 gnd 0.004686f
C834 a_n9628_8799.n107 gnd 0.010134f
C835 a_n9628_8799.n108 gnd 0.010134f
C836 a_n9628_8799.n109 gnd 0.004686f
C837 a_n9628_8799.n111 gnd 0.005584f
C838 a_n9628_8799.n112 gnd 0.010568f
C839 a_n9628_8799.n113 gnd 0.009673f
C840 a_n9628_8799.n114 gnd 0.003669f
C841 a_n9628_8799.n115 gnd 0.250994f
C842 a_n9628_8799.n116 gnd 0.003669f
C843 a_n9628_8799.n117 gnd 0.009673f
C844 a_n9628_8799.n118 gnd 0.010568f
C845 a_n9628_8799.n119 gnd 0.005584f
C846 a_n9628_8799.n121 gnd 0.004686f
C847 a_n9628_8799.n122 gnd 0.010134f
C848 a_n9628_8799.n123 gnd 0.010134f
C849 a_n9628_8799.n124 gnd 0.004686f
C850 a_n9628_8799.n126 gnd 0.005584f
C851 a_n9628_8799.n127 gnd 0.010568f
C852 a_n9628_8799.n128 gnd 0.009673f
C853 a_n9628_8799.n129 gnd 0.003669f
C854 a_n9628_8799.n130 gnd 0.250994f
C855 a_n9628_8799.n131 gnd 0.003669f
C856 a_n9628_8799.n132 gnd 0.009673f
C857 a_n9628_8799.n133 gnd 0.010568f
C858 a_n9628_8799.n134 gnd 0.005584f
C859 a_n9628_8799.n136 gnd 0.004686f
C860 a_n9628_8799.n137 gnd 0.010134f
C861 a_n9628_8799.n138 gnd 0.010134f
C862 a_n9628_8799.n139 gnd 0.004686f
C863 a_n9628_8799.n141 gnd 0.005584f
C864 a_n9628_8799.n142 gnd 0.010568f
C865 a_n9628_8799.n143 gnd 0.009673f
C866 a_n9628_8799.n144 gnd 0.003669f
C867 a_n9628_8799.n145 gnd 0.250994f
C868 a_n9628_8799.t23 gnd 0.144606f
C869 a_n9628_8799.t36 gnd 0.144606f
C870 a_n9628_8799.t32 gnd 0.144606f
C871 a_n9628_8799.n146 gnd 1.14053f
C872 a_n9628_8799.t18 gnd 0.144606f
C873 a_n9628_8799.t17 gnd 0.144606f
C874 a_n9628_8799.n147 gnd 1.13865f
C875 a_n9628_8799.t21 gnd 0.144606f
C876 a_n9628_8799.t24 gnd 0.144606f
C877 a_n9628_8799.n148 gnd 1.13865f
C878 a_n9628_8799.t25 gnd 0.144606f
C879 a_n9628_8799.t33 gnd 0.144606f
C880 a_n9628_8799.n149 gnd 1.13865f
C881 a_n9628_8799.t19 gnd 0.144606f
C882 a_n9628_8799.t38 gnd 0.144606f
C883 a_n9628_8799.n150 gnd 1.13865f
C884 a_n9628_8799.t37 gnd 0.144606f
C885 a_n9628_8799.t22 gnd 0.144606f
C886 a_n9628_8799.n151 gnd 1.13865f
C887 a_n9628_8799.t6 gnd 0.112472f
C888 a_n9628_8799.t1 gnd 0.112472f
C889 a_n9628_8799.n152 gnd 0.996769f
C890 a_n9628_8799.t4 gnd 0.112472f
C891 a_n9628_8799.t12 gnd 0.112472f
C892 a_n9628_8799.n153 gnd 0.993839f
C893 a_n9628_8799.t11 gnd 0.112472f
C894 a_n9628_8799.t15 gnd 0.112472f
C895 a_n9628_8799.n154 gnd 0.996768f
C896 a_n9628_8799.t10 gnd 0.112472f
C897 a_n9628_8799.t8 gnd 0.112472f
C898 a_n9628_8799.n155 gnd 0.993838f
C899 a_n9628_8799.t14 gnd 0.112472f
C900 a_n9628_8799.t7 gnd 0.112472f
C901 a_n9628_8799.n156 gnd 0.996768f
C902 a_n9628_8799.t5 gnd 0.112472f
C903 a_n9628_8799.t9 gnd 0.112472f
C904 a_n9628_8799.n157 gnd 0.993838f
C905 a_n9628_8799.t3 gnd 0.112472f
C906 a_n9628_8799.t2 gnd 0.112472f
C907 a_n9628_8799.n158 gnd 0.993839f
C908 a_n9628_8799.t0 gnd 0.112472f
C909 a_n9628_8799.t13 gnd 0.112472f
C910 a_n9628_8799.n159 gnd 0.993839f
C911 a_n9628_8799.t86 gnd 0.599605f
C912 a_n9628_8799.n160 gnd 0.26995f
C913 a_n9628_8799.t122 gnd 0.599605f
C914 a_n9628_8799.t143 gnd 0.599605f
C915 a_n9628_8799.n161 gnd 0.271884f
C916 a_n9628_8799.t144 gnd 0.599605f
C917 a_n9628_8799.t72 gnd 0.599605f
C918 a_n9628_8799.n162 gnd 0.265064f
C919 a_n9628_8799.t112 gnd 0.599605f
C920 a_n9628_8799.t119 gnd 0.599605f
C921 a_n9628_8799.n163 gnd 0.269054f
C922 a_n9628_8799.t48 gnd 0.599605f
C923 a_n9628_8799.t91 gnd 0.599605f
C924 a_n9628_8799.t89 gnd 0.610954f
C925 a_n9628_8799.n164 gnd 0.251359f
C926 a_n9628_8799.n165 gnd 0.272258f
C927 a_n9628_8799.t123 gnd 0.599605f
C928 a_n9628_8799.n166 gnd 0.26995f
C929 a_n9628_8799.n167 gnd 0.265706f
C930 a_n9628_8799.t87 gnd 0.599605f
C931 a_n9628_8799.n168 gnd 0.264421f
C932 a_n9628_8799.t42 gnd 0.599605f
C933 a_n9628_8799.n169 gnd 0.271628f
C934 a_n9628_8799.t74 gnd 0.599605f
C935 a_n9628_8799.n170 gnd 0.271884f
C936 a_n9628_8799.n171 gnd 0.269488f
C937 a_n9628_8799.t147 gnd 0.599605f
C938 a_n9628_8799.n172 gnd 0.265064f
C939 a_n9628_8799.t108 gnd 0.599605f
C940 a_n9628_8799.n173 gnd 0.269488f
C941 a_n9628_8799.n174 gnd 0.271628f
C942 a_n9628_8799.t90 gnd 0.599605f
C943 a_n9628_8799.n175 gnd 0.269054f
C944 a_n9628_8799.n176 gnd 0.264421f
C945 a_n9628_8799.t142 gnd 0.599605f
C946 a_n9628_8799.n177 gnd 0.265706f
C947 a_n9628_8799.t88 gnd 0.599605f
C948 a_n9628_8799.n178 gnd 0.272258f
C949 a_n9628_8799.t120 gnd 0.610943f
C950 a_n9628_8799.t97 gnd 0.599605f
C951 a_n9628_8799.n179 gnd 0.26995f
C952 a_n9628_8799.t136 gnd 0.599605f
C953 a_n9628_8799.t155 gnd 0.599605f
C954 a_n9628_8799.n180 gnd 0.271884f
C955 a_n9628_8799.t157 gnd 0.599605f
C956 a_n9628_8799.t81 gnd 0.599605f
C957 a_n9628_8799.n181 gnd 0.265064f
C958 a_n9628_8799.t125 gnd 0.599605f
C959 a_n9628_8799.t132 gnd 0.599605f
C960 a_n9628_8799.n182 gnd 0.269054f
C961 a_n9628_8799.t60 gnd 0.599605f
C962 a_n9628_8799.t104 gnd 0.599605f
C963 a_n9628_8799.t102 gnd 0.610954f
C964 a_n9628_8799.n183 gnd 0.251359f
C965 a_n9628_8799.n184 gnd 0.272258f
C966 a_n9628_8799.t140 gnd 0.599605f
C967 a_n9628_8799.n185 gnd 0.26995f
C968 a_n9628_8799.n186 gnd 0.265706f
C969 a_n9628_8799.t98 gnd 0.599605f
C970 a_n9628_8799.n187 gnd 0.264421f
C971 a_n9628_8799.t56 gnd 0.599605f
C972 a_n9628_8799.n188 gnd 0.271628f
C973 a_n9628_8799.t84 gnd 0.599605f
C974 a_n9628_8799.n189 gnd 0.271884f
C975 a_n9628_8799.n190 gnd 0.269488f
C976 a_n9628_8799.t159 gnd 0.599605f
C977 a_n9628_8799.n191 gnd 0.265064f
C978 a_n9628_8799.t121 gnd 0.599605f
C979 a_n9628_8799.n192 gnd 0.269488f
C980 a_n9628_8799.n193 gnd 0.271628f
C981 a_n9628_8799.t103 gnd 0.599605f
C982 a_n9628_8799.n194 gnd 0.269054f
C983 a_n9628_8799.n195 gnd 0.264421f
C984 a_n9628_8799.t154 gnd 0.599605f
C985 a_n9628_8799.n196 gnd 0.265706f
C986 a_n9628_8799.t99 gnd 0.599605f
C987 a_n9628_8799.n197 gnd 0.272258f
C988 a_n9628_8799.t133 gnd 0.610943f
C989 a_n9628_8799.n198 gnd 0.901423f
C990 a_n9628_8799.t63 gnd 0.599605f
C991 a_n9628_8799.n199 gnd 0.26995f
C992 a_n9628_8799.t82 gnd 0.599605f
C993 a_n9628_8799.t115 gnd 0.599605f
C994 a_n9628_8799.n200 gnd 0.271884f
C995 a_n9628_8799.t96 gnd 0.599605f
C996 a_n9628_8799.t100 gnd 0.599605f
C997 a_n9628_8799.n201 gnd 0.265064f
C998 a_n9628_8799.t127 gnd 0.599605f
C999 a_n9628_8799.t43 gnd 0.599605f
C1000 a_n9628_8799.n202 gnd 0.269054f
C1001 a_n9628_8799.t69 gnd 0.599605f
C1002 a_n9628_8799.t52 gnd 0.599605f
C1003 a_n9628_8799.t73 gnd 0.610954f
C1004 a_n9628_8799.n203 gnd 0.251359f
C1005 a_n9628_8799.n204 gnd 0.272258f
C1006 a_n9628_8799.t114 gnd 0.599605f
C1007 a_n9628_8799.n205 gnd 0.26995f
C1008 a_n9628_8799.n206 gnd 0.265706f
C1009 a_n9628_8799.t92 gnd 0.599605f
C1010 a_n9628_8799.n207 gnd 0.264421f
C1011 a_n9628_8799.t109 gnd 0.599605f
C1012 a_n9628_8799.n208 gnd 0.271628f
C1013 a_n9628_8799.t61 gnd 0.599605f
C1014 a_n9628_8799.n209 gnd 0.271884f
C1015 a_n9628_8799.n210 gnd 0.269488f
C1016 a_n9628_8799.t77 gnd 0.599605f
C1017 a_n9628_8799.n211 gnd 0.265064f
C1018 a_n9628_8799.t53 gnd 0.599605f
C1019 a_n9628_8799.n212 gnd 0.269488f
C1020 a_n9628_8799.n213 gnd 0.271628f
C1021 a_n9628_8799.t135 gnd 0.599605f
C1022 a_n9628_8799.n214 gnd 0.269054f
C1023 a_n9628_8799.n215 gnd 0.264421f
C1024 a_n9628_8799.t145 gnd 0.599605f
C1025 a_n9628_8799.n216 gnd 0.265706f
C1026 a_n9628_8799.t40 gnd 0.599605f
C1027 a_n9628_8799.n217 gnd 0.272258f
C1028 a_n9628_8799.t105 gnd 0.610943f
C1029 a_n9628_8799.n218 gnd 1.84873f
C1030 a_n9628_8799.t46 gnd 0.610943f
C1031 a_n9628_8799.t45 gnd 0.599605f
C1032 a_n9628_8799.t131 gnd 0.599605f
C1033 a_n9628_8799.n219 gnd 0.26995f
C1034 a_n9628_8799.t67 gnd 0.599605f
C1035 a_n9628_8799.t50 gnd 0.599605f
C1036 a_n9628_8799.t139 gnd 0.599605f
C1037 a_n9628_8799.n220 gnd 0.269054f
C1038 a_n9628_8799.t94 gnd 0.599605f
C1039 a_n9628_8799.t68 gnd 0.599605f
C1040 a_n9628_8799.t156 gnd 0.599605f
C1041 a_n9628_8799.n221 gnd 0.269488f
C1042 a_n9628_8799.t111 gnd 0.599605f
C1043 a_n9628_8799.t71 gnd 0.599605f
C1044 a_n9628_8799.t150 gnd 0.599605f
C1045 a_n9628_8799.n222 gnd 0.269488f
C1046 a_n9628_8799.t113 gnd 0.599605f
C1047 a_n9628_8799.t85 gnd 0.599605f
C1048 a_n9628_8799.t47 gnd 0.599605f
C1049 a_n9628_8799.n223 gnd 0.269054f
C1050 a_n9628_8799.t134 gnd 0.599605f
C1051 a_n9628_8799.t117 gnd 0.599605f
C1052 a_n9628_8799.t51 gnd 0.599605f
C1053 a_n9628_8799.n224 gnd 0.26995f
C1054 a_n9628_8799.t137 gnd 0.610954f
C1055 a_n9628_8799.n225 gnd 0.251359f
C1056 a_n9628_8799.t141 gnd 0.599605f
C1057 a_n9628_8799.n226 gnd 0.272258f
C1058 a_n9628_8799.n227 gnd 0.265706f
C1059 a_n9628_8799.n228 gnd 0.264421f
C1060 a_n9628_8799.n229 gnd 0.271628f
C1061 a_n9628_8799.n230 gnd 0.271884f
C1062 a_n9628_8799.n231 gnd 0.265064f
C1063 a_n9628_8799.n232 gnd 0.265064f
C1064 a_n9628_8799.n233 gnd 0.271884f
C1065 a_n9628_8799.n234 gnd 0.271628f
C1066 a_n9628_8799.n235 gnd 0.264421f
C1067 a_n9628_8799.n236 gnd 0.265706f
C1068 a_n9628_8799.n237 gnd 0.272258f
C1069 a_n9628_8799.t58 gnd 0.610943f
C1070 a_n9628_8799.t57 gnd 0.599605f
C1071 a_n9628_8799.t148 gnd 0.599605f
C1072 a_n9628_8799.n238 gnd 0.26995f
C1073 a_n9628_8799.t76 gnd 0.599605f
C1074 a_n9628_8799.t65 gnd 0.599605f
C1075 a_n9628_8799.t151 gnd 0.599605f
C1076 a_n9628_8799.n239 gnd 0.269054f
C1077 a_n9628_8799.t107 gnd 0.599605f
C1078 a_n9628_8799.t79 gnd 0.599605f
C1079 a_n9628_8799.t49 gnd 0.599605f
C1080 a_n9628_8799.n240 gnd 0.269488f
C1081 a_n9628_8799.t124 gnd 0.599605f
C1082 a_n9628_8799.t80 gnd 0.599605f
C1083 a_n9628_8799.t41 gnd 0.599605f
C1084 a_n9628_8799.n241 gnd 0.269488f
C1085 a_n9628_8799.t129 gnd 0.599605f
C1086 a_n9628_8799.t95 gnd 0.599605f
C1087 a_n9628_8799.t59 gnd 0.599605f
C1088 a_n9628_8799.n242 gnd 0.269054f
C1089 a_n9628_8799.t149 gnd 0.599605f
C1090 a_n9628_8799.t130 gnd 0.599605f
C1091 a_n9628_8799.t66 gnd 0.599605f
C1092 a_n9628_8799.n243 gnd 0.26995f
C1093 a_n9628_8799.t152 gnd 0.610954f
C1094 a_n9628_8799.n244 gnd 0.251359f
C1095 a_n9628_8799.t153 gnd 0.599605f
C1096 a_n9628_8799.n245 gnd 0.272258f
C1097 a_n9628_8799.n246 gnd 0.265706f
C1098 a_n9628_8799.n247 gnd 0.264421f
C1099 a_n9628_8799.n248 gnd 0.271628f
C1100 a_n9628_8799.n249 gnd 0.271884f
C1101 a_n9628_8799.n250 gnd 0.265064f
C1102 a_n9628_8799.n251 gnd 0.265064f
C1103 a_n9628_8799.n252 gnd 0.271884f
C1104 a_n9628_8799.n253 gnd 0.271628f
C1105 a_n9628_8799.n254 gnd 0.264421f
C1106 a_n9628_8799.n255 gnd 0.265706f
C1107 a_n9628_8799.n256 gnd 0.272258f
C1108 a_n9628_8799.n257 gnd 0.901423f
C1109 a_n9628_8799.t106 gnd 0.610943f
C1110 a_n9628_8799.t128 gnd 0.599605f
C1111 a_n9628_8799.t64 gnd 0.599605f
C1112 a_n9628_8799.n258 gnd 0.26995f
C1113 a_n9628_8799.t146 gnd 0.599605f
C1114 a_n9628_8799.t83 gnd 0.599605f
C1115 a_n9628_8799.t138 gnd 0.599605f
C1116 a_n9628_8799.n259 gnd 0.269054f
C1117 a_n9628_8799.t70 gnd 0.599605f
C1118 a_n9628_8799.t118 gnd 0.599605f
C1119 a_n9628_8799.t55 gnd 0.599605f
C1120 a_n9628_8799.n260 gnd 0.269488f
C1121 a_n9628_8799.t101 gnd 0.599605f
C1122 a_n9628_8799.t78 gnd 0.599605f
C1123 a_n9628_8799.t126 gnd 0.599605f
C1124 a_n9628_8799.n261 gnd 0.269488f
C1125 a_n9628_8799.t62 gnd 0.599605f
C1126 a_n9628_8799.t110 gnd 0.599605f
C1127 a_n9628_8799.t44 gnd 0.599605f
C1128 a_n9628_8799.n262 gnd 0.269054f
C1129 a_n9628_8799.t93 gnd 0.599605f
C1130 a_n9628_8799.t158 gnd 0.599605f
C1131 a_n9628_8799.t116 gnd 0.599605f
C1132 a_n9628_8799.n263 gnd 0.26995f
C1133 a_n9628_8799.t75 gnd 0.610954f
C1134 a_n9628_8799.n264 gnd 0.251359f
C1135 a_n9628_8799.t54 gnd 0.599605f
C1136 a_n9628_8799.n265 gnd 0.272258f
C1137 a_n9628_8799.n266 gnd 0.265706f
C1138 a_n9628_8799.n267 gnd 0.264421f
C1139 a_n9628_8799.n268 gnd 0.271628f
C1140 a_n9628_8799.n269 gnd 0.271884f
C1141 a_n9628_8799.n270 gnd 0.265064f
C1142 a_n9628_8799.n271 gnd 0.265064f
C1143 a_n9628_8799.n272 gnd 0.271884f
C1144 a_n9628_8799.n273 gnd 0.271628f
C1145 a_n9628_8799.n274 gnd 0.264421f
C1146 a_n9628_8799.n275 gnd 0.265706f
C1147 a_n9628_8799.n276 gnd 0.272258f
C1148 a_n9628_8799.n277 gnd 1.42258f
C1149 a_n9628_8799.n278 gnd 17.4279f
C1150 a_n9628_8799.n279 gnd 4.38824f
C1151 a_n9628_8799.n280 gnd 7.65255f
C1152 a_n9628_8799.t34 gnd 0.144606f
C1153 a_n9628_8799.t27 gnd 0.144606f
C1154 a_n9628_8799.n281 gnd 1.14053f
C1155 a_n9628_8799.t26 gnd 0.144606f
C1156 a_n9628_8799.t39 gnd 0.144606f
C1157 a_n9628_8799.n282 gnd 1.13865f
C1158 a_n9628_8799.t31 gnd 0.144606f
C1159 a_n9628_8799.t30 gnd 0.144606f
C1160 a_n9628_8799.n283 gnd 1.13865f
C1161 a_n9628_8799.t28 gnd 0.144606f
C1162 a_n9628_8799.t29 gnd 0.144606f
C1163 a_n9628_8799.n284 gnd 1.13865f
C1164 a_n9628_8799.t20 gnd 0.144606f
C1165 a_n9628_8799.t35 gnd 0.144606f
C1166 a_n9628_8799.n285 gnd 1.13865f
C1167 a_n9628_8799.n286 gnd 3.68856f
C1168 a_n9628_8799.n287 gnd 1.13865f
C1169 a_n9628_8799.t16 gnd 0.144606f
C1170 a_n2804_13878.t29 gnd 0.194878f
C1171 a_n2804_13878.t25 gnd 0.194878f
C1172 a_n2804_13878.t31 gnd 0.194878f
C1173 a_n2804_13878.n0 gnd 1.53703f
C1174 a_n2804_13878.t8 gnd 0.194878f
C1175 a_n2804_13878.t20 gnd 0.194878f
C1176 a_n2804_13878.n1 gnd 1.5345f
C1177 a_n2804_13878.n2 gnd 1.37932f
C1178 a_n2804_13878.t12 gnd 0.194878f
C1179 a_n2804_13878.t22 gnd 0.194878f
C1180 a_n2804_13878.n3 gnd 1.53612f
C1181 a_n2804_13878.t27 gnd 0.194878f
C1182 a_n2804_13878.t17 gnd 0.194878f
C1183 a_n2804_13878.n4 gnd 1.5345f
C1184 a_n2804_13878.n5 gnd 2.14416f
C1185 a_n2804_13878.t23 gnd 0.194878f
C1186 a_n2804_13878.t16 gnd 0.194878f
C1187 a_n2804_13878.n6 gnd 1.5345f
C1188 a_n2804_13878.n7 gnd 1.04587f
C1189 a_n2804_13878.t10 gnd 0.194878f
C1190 a_n2804_13878.t13 gnd 0.194878f
C1191 a_n2804_13878.n8 gnd 1.5345f
C1192 a_n2804_13878.n9 gnd 1.04587f
C1193 a_n2804_13878.t26 gnd 0.194878f
C1194 a_n2804_13878.t11 gnd 0.194878f
C1195 a_n2804_13878.n10 gnd 1.5345f
C1196 a_n2804_13878.n11 gnd 1.04587f
C1197 a_n2804_13878.t21 gnd 0.194878f
C1198 a_n2804_13878.t9 gnd 0.194878f
C1199 a_n2804_13878.n12 gnd 1.5345f
C1200 a_n2804_13878.n13 gnd 4.90989f
C1201 a_n2804_13878.t1 gnd 1.82474f
C1202 a_n2804_13878.t4 gnd 0.194878f
C1203 a_n2804_13878.t5 gnd 0.194878f
C1204 a_n2804_13878.n14 gnd 1.37272f
C1205 a_n2804_13878.n15 gnd 1.53381f
C1206 a_n2804_13878.t0 gnd 1.8211f
C1207 a_n2804_13878.n16 gnd 0.771835f
C1208 a_n2804_13878.t3 gnd 1.8211f
C1209 a_n2804_13878.n17 gnd 0.771835f
C1210 a_n2804_13878.t6 gnd 0.194878f
C1211 a_n2804_13878.t7 gnd 0.194878f
C1212 a_n2804_13878.n18 gnd 1.37272f
C1213 a_n2804_13878.n19 gnd 0.77931f
C1214 a_n2804_13878.t2 gnd 1.8211f
C1215 a_n2804_13878.n20 gnd 2.86287f
C1216 a_n2804_13878.n21 gnd 3.75497f
C1217 a_n2804_13878.t15 gnd 0.194878f
C1218 a_n2804_13878.t24 gnd 0.194878f
C1219 a_n2804_13878.n22 gnd 1.53449f
C1220 a_n2804_13878.n23 gnd 2.50654f
C1221 a_n2804_13878.t28 gnd 0.194878f
C1222 a_n2804_13878.t14 gnd 0.194878f
C1223 a_n2804_13878.n24 gnd 1.5345f
C1224 a_n2804_13878.n25 gnd 0.679894f
C1225 a_n2804_13878.t18 gnd 0.194878f
C1226 a_n2804_13878.t19 gnd 0.194878f
C1227 a_n2804_13878.n26 gnd 1.5345f
C1228 a_n2804_13878.n27 gnd 0.679894f
C1229 a_n2804_13878.n28 gnd 0.679892f
C1230 a_n2804_13878.n29 gnd 1.5345f
C1231 a_n2804_13878.t30 gnd 0.194878f
C1232 vdd.t280 gnd 0.036923f
C1233 vdd.t261 gnd 0.036923f
C1234 vdd.n0 gnd 0.291219f
C1235 vdd.t239 gnd 0.036923f
C1236 vdd.t276 gnd 0.036923f
C1237 vdd.n1 gnd 0.290739f
C1238 vdd.n2 gnd 0.268116f
C1239 vdd.t257 gnd 0.036923f
C1240 vdd.t287 gnd 0.036923f
C1241 vdd.n3 gnd 0.290739f
C1242 vdd.n4 gnd 0.135597f
C1243 vdd.t285 gnd 0.036923f
C1244 vdd.t265 gnd 0.036923f
C1245 vdd.n5 gnd 0.290739f
C1246 vdd.n6 gnd 0.127232f
C1247 vdd.t291 gnd 0.036923f
C1248 vdd.t255 gnd 0.036923f
C1249 vdd.n7 gnd 0.291219f
C1250 vdd.t263 gnd 0.036923f
C1251 vdd.t283 gnd 0.036923f
C1252 vdd.n8 gnd 0.290739f
C1253 vdd.n9 gnd 0.268116f
C1254 vdd.t272 gnd 0.036923f
C1255 vdd.t245 gnd 0.036923f
C1256 vdd.n10 gnd 0.290739f
C1257 vdd.n11 gnd 0.135597f
C1258 vdd.t241 gnd 0.036923f
C1259 vdd.t270 gnd 0.036923f
C1260 vdd.n12 gnd 0.290739f
C1261 vdd.n13 gnd 0.127232f
C1262 vdd.n14 gnd 0.089951f
C1263 vdd.t14 gnd 0.020513f
C1264 vdd.t10 gnd 0.020513f
C1265 vdd.n15 gnd 0.188813f
C1266 vdd.t16 gnd 0.020513f
C1267 vdd.t11 gnd 0.020513f
C1268 vdd.n16 gnd 0.18826f
C1269 vdd.n17 gnd 0.327631f
C1270 vdd.t21 gnd 0.020513f
C1271 vdd.t17 gnd 0.020513f
C1272 vdd.n18 gnd 0.18826f
C1273 vdd.n19 gnd 0.135545f
C1274 vdd.t8 gnd 0.020513f
C1275 vdd.t22 gnd 0.020513f
C1276 vdd.n20 gnd 0.188813f
C1277 vdd.t9 gnd 0.020513f
C1278 vdd.t18 gnd 0.020513f
C1279 vdd.n21 gnd 0.18826f
C1280 vdd.n22 gnd 0.327631f
C1281 vdd.t19 gnd 0.020513f
C1282 vdd.t13 gnd 0.020513f
C1283 vdd.n23 gnd 0.18826f
C1284 vdd.n24 gnd 0.135545f
C1285 vdd.t12 gnd 0.020513f
C1286 vdd.t15 gnd 0.020513f
C1287 vdd.n25 gnd 0.18826f
C1288 vdd.t20 gnd 0.020513f
C1289 vdd.t23 gnd 0.020513f
C1290 vdd.n26 gnd 0.18826f
C1291 vdd.n27 gnd 21.743f
C1292 vdd.n28 gnd 8.48534f
C1293 vdd.n29 gnd 0.005595f
C1294 vdd.n30 gnd 0.005192f
C1295 vdd.n31 gnd 0.002872f
C1296 vdd.n32 gnd 0.006594f
C1297 vdd.n33 gnd 0.00279f
C1298 vdd.n34 gnd 0.002954f
C1299 vdd.n35 gnd 0.005192f
C1300 vdd.n36 gnd 0.00279f
C1301 vdd.n37 gnd 0.006594f
C1302 vdd.n38 gnd 0.002954f
C1303 vdd.n39 gnd 0.005192f
C1304 vdd.n40 gnd 0.00279f
C1305 vdd.n41 gnd 0.004945f
C1306 vdd.n42 gnd 0.00496f
C1307 vdd.t32 gnd 0.014167f
C1308 vdd.n43 gnd 0.03152f
C1309 vdd.n44 gnd 0.16404f
C1310 vdd.n45 gnd 0.00279f
C1311 vdd.n46 gnd 0.002954f
C1312 vdd.n47 gnd 0.006594f
C1313 vdd.n48 gnd 0.006594f
C1314 vdd.n49 gnd 0.002954f
C1315 vdd.n50 gnd 0.00279f
C1316 vdd.n51 gnd 0.005192f
C1317 vdd.n52 gnd 0.005192f
C1318 vdd.n53 gnd 0.00279f
C1319 vdd.n54 gnd 0.002954f
C1320 vdd.n55 gnd 0.006594f
C1321 vdd.n56 gnd 0.006594f
C1322 vdd.n57 gnd 0.002954f
C1323 vdd.n58 gnd 0.00279f
C1324 vdd.n59 gnd 0.005192f
C1325 vdd.n60 gnd 0.005192f
C1326 vdd.n61 gnd 0.00279f
C1327 vdd.n62 gnd 0.002954f
C1328 vdd.n63 gnd 0.006594f
C1329 vdd.n64 gnd 0.006594f
C1330 vdd.n65 gnd 0.01559f
C1331 vdd.n66 gnd 0.002872f
C1332 vdd.n67 gnd 0.00279f
C1333 vdd.n68 gnd 0.013419f
C1334 vdd.n69 gnd 0.009368f
C1335 vdd.t28 gnd 0.032821f
C1336 vdd.t294 gnd 0.032821f
C1337 vdd.n70 gnd 0.225566f
C1338 vdd.n71 gnd 0.177373f
C1339 vdd.t197 gnd 0.032821f
C1340 vdd.t223 gnd 0.032821f
C1341 vdd.n72 gnd 0.225566f
C1342 vdd.n73 gnd 0.143139f
C1343 vdd.t25 gnd 0.032821f
C1344 vdd.t226 gnd 0.032821f
C1345 vdd.n74 gnd 0.225566f
C1346 vdd.n75 gnd 0.143139f
C1347 vdd.t302 gnd 0.032821f
C1348 vdd.t231 gnd 0.032821f
C1349 vdd.n76 gnd 0.225566f
C1350 vdd.n77 gnd 0.143139f
C1351 vdd.t171 gnd 0.032821f
C1352 vdd.t199 gnd 0.032821f
C1353 vdd.n78 gnd 0.225566f
C1354 vdd.n79 gnd 0.143139f
C1355 vdd.t188 gnd 0.032821f
C1356 vdd.t292 gnd 0.032821f
C1357 vdd.n80 gnd 0.225566f
C1358 vdd.n81 gnd 0.143139f
C1359 vdd.t190 gnd 0.032821f
C1360 vdd.t234 gnd 0.032821f
C1361 vdd.n82 gnd 0.225566f
C1362 vdd.n83 gnd 0.143139f
C1363 vdd.t7 gnd 0.032821f
C1364 vdd.t195 gnd 0.032821f
C1365 vdd.n84 gnd 0.225566f
C1366 vdd.n85 gnd 0.143139f
C1367 vdd.t1 gnd 0.032821f
C1368 vdd.t230 gnd 0.032821f
C1369 vdd.n86 gnd 0.225566f
C1370 vdd.n87 gnd 0.143139f
C1371 vdd.n88 gnd 0.005595f
C1372 vdd.n89 gnd 0.005192f
C1373 vdd.n90 gnd 0.002872f
C1374 vdd.n91 gnd 0.006594f
C1375 vdd.n92 gnd 0.00279f
C1376 vdd.n93 gnd 0.002954f
C1377 vdd.n94 gnd 0.005192f
C1378 vdd.n95 gnd 0.00279f
C1379 vdd.n96 gnd 0.006594f
C1380 vdd.n97 gnd 0.002954f
C1381 vdd.n98 gnd 0.005192f
C1382 vdd.n99 gnd 0.00279f
C1383 vdd.n100 gnd 0.004945f
C1384 vdd.n101 gnd 0.00496f
C1385 vdd.t202 gnd 0.014167f
C1386 vdd.n102 gnd 0.03152f
C1387 vdd.n103 gnd 0.16404f
C1388 vdd.n104 gnd 0.00279f
C1389 vdd.n105 gnd 0.002954f
C1390 vdd.n106 gnd 0.006594f
C1391 vdd.n107 gnd 0.006594f
C1392 vdd.n108 gnd 0.002954f
C1393 vdd.n109 gnd 0.00279f
C1394 vdd.n110 gnd 0.005192f
C1395 vdd.n111 gnd 0.005192f
C1396 vdd.n112 gnd 0.00279f
C1397 vdd.n113 gnd 0.002954f
C1398 vdd.n114 gnd 0.006594f
C1399 vdd.n115 gnd 0.006594f
C1400 vdd.n116 gnd 0.002954f
C1401 vdd.n117 gnd 0.00279f
C1402 vdd.n118 gnd 0.005192f
C1403 vdd.n119 gnd 0.005192f
C1404 vdd.n120 gnd 0.00279f
C1405 vdd.n121 gnd 0.002954f
C1406 vdd.n122 gnd 0.006594f
C1407 vdd.n123 gnd 0.006594f
C1408 vdd.n124 gnd 0.01559f
C1409 vdd.n125 gnd 0.002872f
C1410 vdd.n126 gnd 0.00279f
C1411 vdd.n127 gnd 0.013419f
C1412 vdd.n128 gnd 0.009074f
C1413 vdd.n129 gnd 0.106496f
C1414 vdd.n130 gnd 0.005595f
C1415 vdd.n131 gnd 0.005192f
C1416 vdd.n132 gnd 0.002872f
C1417 vdd.n133 gnd 0.006594f
C1418 vdd.n134 gnd 0.00279f
C1419 vdd.n135 gnd 0.002954f
C1420 vdd.n136 gnd 0.005192f
C1421 vdd.n137 gnd 0.00279f
C1422 vdd.n138 gnd 0.006594f
C1423 vdd.n139 gnd 0.002954f
C1424 vdd.n140 gnd 0.005192f
C1425 vdd.n141 gnd 0.00279f
C1426 vdd.n142 gnd 0.004945f
C1427 vdd.n143 gnd 0.00496f
C1428 vdd.t81 gnd 0.014167f
C1429 vdd.n144 gnd 0.03152f
C1430 vdd.n145 gnd 0.16404f
C1431 vdd.n146 gnd 0.00279f
C1432 vdd.n147 gnd 0.002954f
C1433 vdd.n148 gnd 0.006594f
C1434 vdd.n149 gnd 0.006594f
C1435 vdd.n150 gnd 0.002954f
C1436 vdd.n151 gnd 0.00279f
C1437 vdd.n152 gnd 0.005192f
C1438 vdd.n153 gnd 0.005192f
C1439 vdd.n154 gnd 0.00279f
C1440 vdd.n155 gnd 0.002954f
C1441 vdd.n156 gnd 0.006594f
C1442 vdd.n157 gnd 0.006594f
C1443 vdd.n158 gnd 0.002954f
C1444 vdd.n159 gnd 0.00279f
C1445 vdd.n160 gnd 0.005192f
C1446 vdd.n161 gnd 0.005192f
C1447 vdd.n162 gnd 0.00279f
C1448 vdd.n163 gnd 0.002954f
C1449 vdd.n164 gnd 0.006594f
C1450 vdd.n165 gnd 0.006594f
C1451 vdd.n166 gnd 0.01559f
C1452 vdd.n167 gnd 0.002872f
C1453 vdd.n168 gnd 0.00279f
C1454 vdd.n169 gnd 0.013419f
C1455 vdd.n170 gnd 0.009368f
C1456 vdd.t205 gnd 0.032821f
C1457 vdd.t63 gnd 0.032821f
C1458 vdd.n171 gnd 0.225566f
C1459 vdd.n172 gnd 0.177373f
C1460 vdd.t74 gnd 0.032821f
C1461 vdd.t295 gnd 0.032821f
C1462 vdd.n173 gnd 0.225566f
C1463 vdd.n174 gnd 0.143139f
C1464 vdd.t41 gnd 0.032821f
C1465 vdd.t34 gnd 0.032821f
C1466 vdd.n175 gnd 0.225566f
C1467 vdd.n176 gnd 0.143139f
C1468 vdd.t200 gnd 0.032821f
C1469 vdd.t218 gnd 0.032821f
C1470 vdd.n177 gnd 0.225566f
C1471 vdd.n178 gnd 0.143139f
C1472 vdd.t300 gnd 0.032821f
C1473 vdd.t71 gnd 0.032821f
C1474 vdd.n179 gnd 0.225566f
C1475 vdd.n180 gnd 0.143139f
C1476 vdd.t69 gnd 0.032821f
C1477 vdd.t30 gnd 0.032821f
C1478 vdd.n181 gnd 0.225566f
C1479 vdd.n182 gnd 0.143139f
C1480 vdd.t173 gnd 0.032821f
C1481 vdd.t82 gnd 0.032821f
C1482 vdd.n183 gnd 0.225566f
C1483 vdd.n184 gnd 0.143139f
C1484 vdd.t64 gnd 0.032821f
C1485 vdd.t177 gnd 0.032821f
C1486 vdd.n185 gnd 0.225566f
C1487 vdd.n186 gnd 0.143139f
C1488 vdd.t53 gnd 0.032821f
C1489 vdd.t187 gnd 0.032821f
C1490 vdd.n187 gnd 0.225566f
C1491 vdd.n188 gnd 0.143139f
C1492 vdd.n189 gnd 0.005595f
C1493 vdd.n190 gnd 0.005192f
C1494 vdd.n191 gnd 0.002872f
C1495 vdd.n192 gnd 0.006594f
C1496 vdd.n193 gnd 0.00279f
C1497 vdd.n194 gnd 0.002954f
C1498 vdd.n195 gnd 0.005192f
C1499 vdd.n196 gnd 0.00279f
C1500 vdd.n197 gnd 0.006594f
C1501 vdd.n198 gnd 0.002954f
C1502 vdd.n199 gnd 0.005192f
C1503 vdd.n200 gnd 0.00279f
C1504 vdd.n201 gnd 0.004945f
C1505 vdd.n202 gnd 0.00496f
C1506 vdd.t185 gnd 0.014167f
C1507 vdd.n203 gnd 0.03152f
C1508 vdd.n204 gnd 0.16404f
C1509 vdd.n205 gnd 0.00279f
C1510 vdd.n206 gnd 0.002954f
C1511 vdd.n207 gnd 0.006594f
C1512 vdd.n208 gnd 0.006594f
C1513 vdd.n209 gnd 0.002954f
C1514 vdd.n210 gnd 0.00279f
C1515 vdd.n211 gnd 0.005192f
C1516 vdd.n212 gnd 0.005192f
C1517 vdd.n213 gnd 0.00279f
C1518 vdd.n214 gnd 0.002954f
C1519 vdd.n215 gnd 0.006594f
C1520 vdd.n216 gnd 0.006594f
C1521 vdd.n217 gnd 0.002954f
C1522 vdd.n218 gnd 0.00279f
C1523 vdd.n219 gnd 0.005192f
C1524 vdd.n220 gnd 0.005192f
C1525 vdd.n221 gnd 0.00279f
C1526 vdd.n222 gnd 0.002954f
C1527 vdd.n223 gnd 0.006594f
C1528 vdd.n224 gnd 0.006594f
C1529 vdd.n225 gnd 0.01559f
C1530 vdd.n226 gnd 0.002872f
C1531 vdd.n227 gnd 0.00279f
C1532 vdd.n228 gnd 0.013419f
C1533 vdd.n229 gnd 0.009074f
C1534 vdd.n230 gnd 0.063354f
C1535 vdd.n231 gnd 0.228283f
C1536 vdd.n232 gnd 0.005595f
C1537 vdd.n233 gnd 0.005192f
C1538 vdd.n234 gnd 0.002872f
C1539 vdd.n235 gnd 0.006594f
C1540 vdd.n236 gnd 0.00279f
C1541 vdd.n237 gnd 0.002954f
C1542 vdd.n238 gnd 0.005192f
C1543 vdd.n239 gnd 0.00279f
C1544 vdd.n240 gnd 0.006594f
C1545 vdd.n241 gnd 0.002954f
C1546 vdd.n242 gnd 0.005192f
C1547 vdd.n243 gnd 0.00279f
C1548 vdd.n244 gnd 0.004945f
C1549 vdd.n245 gnd 0.00496f
C1550 vdd.t65 gnd 0.014167f
C1551 vdd.n246 gnd 0.03152f
C1552 vdd.n247 gnd 0.16404f
C1553 vdd.n248 gnd 0.00279f
C1554 vdd.n249 gnd 0.002954f
C1555 vdd.n250 gnd 0.006594f
C1556 vdd.n251 gnd 0.006594f
C1557 vdd.n252 gnd 0.002954f
C1558 vdd.n253 gnd 0.00279f
C1559 vdd.n254 gnd 0.005192f
C1560 vdd.n255 gnd 0.005192f
C1561 vdd.n256 gnd 0.00279f
C1562 vdd.n257 gnd 0.002954f
C1563 vdd.n258 gnd 0.006594f
C1564 vdd.n259 gnd 0.006594f
C1565 vdd.n260 gnd 0.002954f
C1566 vdd.n261 gnd 0.00279f
C1567 vdd.n262 gnd 0.005192f
C1568 vdd.n263 gnd 0.005192f
C1569 vdd.n264 gnd 0.00279f
C1570 vdd.n265 gnd 0.002954f
C1571 vdd.n266 gnd 0.006594f
C1572 vdd.n267 gnd 0.006594f
C1573 vdd.n268 gnd 0.01559f
C1574 vdd.n269 gnd 0.002872f
C1575 vdd.n270 gnd 0.00279f
C1576 vdd.n271 gnd 0.013419f
C1577 vdd.n272 gnd 0.009368f
C1578 vdd.t235 gnd 0.032821f
C1579 vdd.t178 gnd 0.032821f
C1580 vdd.n273 gnd 0.225566f
C1581 vdd.n274 gnd 0.177373f
C1582 vdd.t55 gnd 0.032821f
C1583 vdd.t232 gnd 0.032821f
C1584 vdd.n275 gnd 0.225566f
C1585 vdd.n276 gnd 0.143139f
C1586 vdd.t26 gnd 0.032821f
C1587 vdd.t172 gnd 0.032821f
C1588 vdd.n277 gnd 0.225566f
C1589 vdd.n278 gnd 0.143139f
C1590 vdd.t78 gnd 0.032821f
C1591 vdd.t160 gnd 0.032821f
C1592 vdd.n279 gnd 0.225566f
C1593 vdd.n280 gnd 0.143139f
C1594 vdd.t191 gnd 0.032821f
C1595 vdd.t227 gnd 0.032821f
C1596 vdd.n281 gnd 0.225566f
C1597 vdd.n282 gnd 0.143139f
C1598 vdd.t40 gnd 0.032821f
C1599 vdd.t181 gnd 0.032821f
C1600 vdd.n283 gnd 0.225566f
C1601 vdd.n284 gnd 0.143139f
C1602 vdd.t52 gnd 0.032821f
C1603 vdd.t67 gnd 0.032821f
C1604 vdd.n285 gnd 0.225566f
C1605 vdd.n286 gnd 0.143139f
C1606 vdd.t42 gnd 0.032821f
C1607 vdd.t3 gnd 0.032821f
C1608 vdd.n287 gnd 0.225566f
C1609 vdd.n288 gnd 0.143139f
C1610 vdd.t233 gnd 0.032821f
C1611 vdd.t297 gnd 0.032821f
C1612 vdd.n289 gnd 0.225566f
C1613 vdd.n290 gnd 0.143139f
C1614 vdd.n291 gnd 0.005595f
C1615 vdd.n292 gnd 0.005192f
C1616 vdd.n293 gnd 0.002872f
C1617 vdd.n294 gnd 0.006594f
C1618 vdd.n295 gnd 0.00279f
C1619 vdd.n296 gnd 0.002954f
C1620 vdd.n297 gnd 0.005192f
C1621 vdd.n298 gnd 0.00279f
C1622 vdd.n299 gnd 0.006594f
C1623 vdd.n300 gnd 0.002954f
C1624 vdd.n301 gnd 0.005192f
C1625 vdd.n302 gnd 0.00279f
C1626 vdd.n303 gnd 0.004945f
C1627 vdd.n304 gnd 0.00496f
C1628 vdd.t210 gnd 0.014167f
C1629 vdd.n305 gnd 0.03152f
C1630 vdd.n306 gnd 0.16404f
C1631 vdd.n307 gnd 0.00279f
C1632 vdd.n308 gnd 0.002954f
C1633 vdd.n309 gnd 0.006594f
C1634 vdd.n310 gnd 0.006594f
C1635 vdd.n311 gnd 0.002954f
C1636 vdd.n312 gnd 0.00279f
C1637 vdd.n313 gnd 0.005192f
C1638 vdd.n314 gnd 0.005192f
C1639 vdd.n315 gnd 0.00279f
C1640 vdd.n316 gnd 0.002954f
C1641 vdd.n317 gnd 0.006594f
C1642 vdd.n318 gnd 0.006594f
C1643 vdd.n319 gnd 0.002954f
C1644 vdd.n320 gnd 0.00279f
C1645 vdd.n321 gnd 0.005192f
C1646 vdd.n322 gnd 0.005192f
C1647 vdd.n323 gnd 0.00279f
C1648 vdd.n324 gnd 0.002954f
C1649 vdd.n325 gnd 0.006594f
C1650 vdd.n326 gnd 0.006594f
C1651 vdd.n327 gnd 0.01559f
C1652 vdd.n328 gnd 0.002872f
C1653 vdd.n329 gnd 0.00279f
C1654 vdd.n330 gnd 0.013419f
C1655 vdd.n331 gnd 0.009074f
C1656 vdd.n332 gnd 0.063354f
C1657 vdd.n333 gnd 0.261334f
C1658 vdd.n334 gnd 0.007835f
C1659 vdd.n335 gnd 0.010194f
C1660 vdd.n336 gnd 0.008205f
C1661 vdd.n337 gnd 0.008205f
C1662 vdd.n338 gnd 0.010194f
C1663 vdd.n339 gnd 0.010194f
C1664 vdd.n340 gnd 0.744892f
C1665 vdd.n341 gnd 0.010194f
C1666 vdd.n342 gnd 0.010194f
C1667 vdd.n343 gnd 0.010194f
C1668 vdd.n344 gnd 0.8074f
C1669 vdd.n345 gnd 0.010194f
C1670 vdd.n346 gnd 0.010194f
C1671 vdd.n347 gnd 0.010194f
C1672 vdd.n348 gnd 0.010194f
C1673 vdd.n349 gnd 0.008205f
C1674 vdd.n350 gnd 0.010194f
C1675 vdd.t29 gnd 0.520903f
C1676 vdd.n351 gnd 0.010194f
C1677 vdd.n352 gnd 0.010194f
C1678 vdd.n353 gnd 0.010194f
C1679 vdd.t66 gnd 0.520903f
C1680 vdd.n354 gnd 0.010194f
C1681 vdd.n355 gnd 0.010194f
C1682 vdd.n356 gnd 0.010194f
C1683 vdd.n357 gnd 0.010194f
C1684 vdd.n358 gnd 0.010194f
C1685 vdd.n359 gnd 0.008205f
C1686 vdd.n360 gnd 0.010194f
C1687 vdd.n361 gnd 0.588621f
C1688 vdd.n362 gnd 0.010194f
C1689 vdd.n363 gnd 0.010194f
C1690 vdd.n364 gnd 0.010194f
C1691 vdd.t2 gnd 0.520903f
C1692 vdd.n365 gnd 0.010194f
C1693 vdd.n366 gnd 0.010194f
C1694 vdd.n367 gnd 0.010194f
C1695 vdd.n368 gnd 0.010194f
C1696 vdd.n369 gnd 0.010194f
C1697 vdd.n370 gnd 0.008205f
C1698 vdd.n371 gnd 0.010194f
C1699 vdd.t0 gnd 0.520903f
C1700 vdd.n372 gnd 0.010194f
C1701 vdd.n373 gnd 0.010194f
C1702 vdd.n374 gnd 0.010194f
C1703 vdd.n375 gnd 0.609457f
C1704 vdd.n376 gnd 0.010194f
C1705 vdd.n377 gnd 0.010194f
C1706 vdd.n378 gnd 0.010194f
C1707 vdd.n379 gnd 0.010194f
C1708 vdd.n380 gnd 0.010194f
C1709 vdd.n381 gnd 0.008205f
C1710 vdd.n382 gnd 0.010194f
C1711 vdd.t184 gnd 0.520903f
C1712 vdd.n383 gnd 0.010194f
C1713 vdd.n384 gnd 0.010194f
C1714 vdd.n385 gnd 0.010194f
C1715 vdd.n386 gnd 0.526112f
C1716 vdd.n387 gnd 0.010194f
C1717 vdd.n388 gnd 0.010194f
C1718 vdd.n389 gnd 0.010194f
C1719 vdd.n390 gnd 0.010194f
C1720 vdd.n391 gnd 0.024661f
C1721 vdd.n392 gnd 0.025189f
C1722 vdd.t96 gnd 0.520903f
C1723 vdd.n393 gnd 0.024661f
C1724 vdd.n425 gnd 0.010194f
C1725 vdd.t124 gnd 0.125416f
C1726 vdd.t123 gnd 0.134036f
C1727 vdd.t122 gnd 0.163792f
C1728 vdd.n426 gnd 0.209958f
C1729 vdd.n427 gnd 0.177224f
C1730 vdd.n428 gnd 0.013457f
C1731 vdd.n429 gnd 0.010194f
C1732 vdd.n430 gnd 0.008205f
C1733 vdd.n431 gnd 0.010194f
C1734 vdd.n432 gnd 0.008205f
C1735 vdd.n433 gnd 0.010194f
C1736 vdd.n434 gnd 0.008205f
C1737 vdd.n435 gnd 0.010194f
C1738 vdd.n436 gnd 0.008205f
C1739 vdd.n437 gnd 0.010194f
C1740 vdd.n438 gnd 0.008205f
C1741 vdd.n439 gnd 0.010194f
C1742 vdd.t98 gnd 0.125416f
C1743 vdd.t97 gnd 0.134036f
C1744 vdd.t95 gnd 0.163792f
C1745 vdd.n440 gnd 0.209958f
C1746 vdd.n441 gnd 0.177224f
C1747 vdd.n442 gnd 0.008205f
C1748 vdd.n443 gnd 0.010194f
C1749 vdd.n444 gnd 0.008205f
C1750 vdd.n445 gnd 0.010194f
C1751 vdd.n446 gnd 0.008205f
C1752 vdd.n447 gnd 0.010194f
C1753 vdd.n448 gnd 0.008205f
C1754 vdd.n449 gnd 0.010194f
C1755 vdd.n450 gnd 0.008205f
C1756 vdd.n451 gnd 0.010194f
C1757 vdd.t104 gnd 0.125416f
C1758 vdd.t103 gnd 0.134036f
C1759 vdd.t102 gnd 0.163792f
C1760 vdd.n452 gnd 0.209958f
C1761 vdd.n453 gnd 0.177224f
C1762 vdd.n454 gnd 0.017559f
C1763 vdd.n455 gnd 0.010194f
C1764 vdd.n456 gnd 0.008205f
C1765 vdd.n457 gnd 0.010194f
C1766 vdd.n458 gnd 0.008205f
C1767 vdd.n459 gnd 0.010194f
C1768 vdd.n460 gnd 0.008205f
C1769 vdd.n461 gnd 0.010194f
C1770 vdd.n462 gnd 0.008205f
C1771 vdd.n463 gnd 0.010194f
C1772 vdd.n464 gnd 0.025189f
C1773 vdd.n465 gnd 0.00681f
C1774 vdd.n466 gnd 0.008205f
C1775 vdd.n467 gnd 0.010194f
C1776 vdd.n468 gnd 0.010194f
C1777 vdd.n469 gnd 0.008205f
C1778 vdd.n470 gnd 0.010194f
C1779 vdd.n471 gnd 0.010194f
C1780 vdd.n472 gnd 0.010194f
C1781 vdd.n473 gnd 0.010194f
C1782 vdd.n474 gnd 0.010194f
C1783 vdd.n475 gnd 0.008205f
C1784 vdd.n476 gnd 0.008205f
C1785 vdd.n477 gnd 0.010194f
C1786 vdd.n478 gnd 0.010194f
C1787 vdd.n479 gnd 0.008205f
C1788 vdd.n480 gnd 0.010194f
C1789 vdd.n481 gnd 0.010194f
C1790 vdd.n482 gnd 0.010194f
C1791 vdd.n483 gnd 0.010194f
C1792 vdd.n484 gnd 0.010194f
C1793 vdd.n485 gnd 0.008205f
C1794 vdd.n486 gnd 0.008205f
C1795 vdd.n487 gnd 0.010194f
C1796 vdd.n488 gnd 0.010194f
C1797 vdd.n489 gnd 0.008205f
C1798 vdd.n490 gnd 0.010194f
C1799 vdd.n491 gnd 0.010194f
C1800 vdd.n492 gnd 0.010194f
C1801 vdd.n493 gnd 0.010194f
C1802 vdd.n494 gnd 0.010194f
C1803 vdd.n495 gnd 0.008205f
C1804 vdd.n496 gnd 0.008205f
C1805 vdd.n497 gnd 0.010194f
C1806 vdd.n498 gnd 0.010194f
C1807 vdd.n499 gnd 0.008205f
C1808 vdd.n500 gnd 0.010194f
C1809 vdd.n501 gnd 0.010194f
C1810 vdd.n502 gnd 0.010194f
C1811 vdd.n503 gnd 0.010194f
C1812 vdd.n504 gnd 0.010194f
C1813 vdd.n505 gnd 0.008205f
C1814 vdd.n506 gnd 0.008205f
C1815 vdd.n507 gnd 0.010194f
C1816 vdd.n508 gnd 0.010194f
C1817 vdd.n509 gnd 0.006851f
C1818 vdd.n510 gnd 0.010194f
C1819 vdd.n511 gnd 0.010194f
C1820 vdd.n512 gnd 0.010194f
C1821 vdd.n513 gnd 0.010194f
C1822 vdd.n514 gnd 0.010194f
C1823 vdd.n515 gnd 0.006851f
C1824 vdd.n516 gnd 0.008205f
C1825 vdd.n517 gnd 0.010194f
C1826 vdd.n518 gnd 0.010194f
C1827 vdd.n519 gnd 0.008205f
C1828 vdd.n520 gnd 0.010194f
C1829 vdd.n521 gnd 0.010194f
C1830 vdd.n522 gnd 0.010194f
C1831 vdd.n523 gnd 0.010194f
C1832 vdd.n524 gnd 0.010194f
C1833 vdd.n525 gnd 0.008205f
C1834 vdd.n526 gnd 0.008205f
C1835 vdd.n527 gnd 0.010194f
C1836 vdd.n528 gnd 0.010194f
C1837 vdd.n529 gnd 0.008205f
C1838 vdd.n530 gnd 0.010194f
C1839 vdd.n531 gnd 0.010194f
C1840 vdd.n532 gnd 0.010194f
C1841 vdd.n533 gnd 0.010194f
C1842 vdd.n534 gnd 0.010194f
C1843 vdd.n535 gnd 0.008205f
C1844 vdd.n536 gnd 0.008205f
C1845 vdd.n537 gnd 0.010194f
C1846 vdd.n538 gnd 0.010194f
C1847 vdd.n539 gnd 0.008205f
C1848 vdd.n540 gnd 0.010194f
C1849 vdd.n541 gnd 0.010194f
C1850 vdd.n542 gnd 0.010194f
C1851 vdd.n543 gnd 0.010194f
C1852 vdd.n544 gnd 0.010194f
C1853 vdd.n545 gnd 0.008205f
C1854 vdd.n546 gnd 0.008205f
C1855 vdd.n547 gnd 0.010194f
C1856 vdd.n548 gnd 0.010194f
C1857 vdd.n549 gnd 0.008205f
C1858 vdd.n550 gnd 0.010194f
C1859 vdd.n551 gnd 0.010194f
C1860 vdd.n552 gnd 0.010194f
C1861 vdd.n553 gnd 0.010194f
C1862 vdd.n554 gnd 0.010194f
C1863 vdd.n555 gnd 0.008205f
C1864 vdd.n556 gnd 0.008205f
C1865 vdd.n557 gnd 0.010194f
C1866 vdd.n558 gnd 0.010194f
C1867 vdd.n559 gnd 0.008205f
C1868 vdd.n560 gnd 0.010194f
C1869 vdd.n561 gnd 0.010194f
C1870 vdd.n562 gnd 0.010194f
C1871 vdd.n563 gnd 0.010194f
C1872 vdd.n564 gnd 0.010194f
C1873 vdd.n565 gnd 0.00558f
C1874 vdd.n566 gnd 0.017559f
C1875 vdd.n567 gnd 0.010194f
C1876 vdd.n568 gnd 0.010194f
C1877 vdd.n569 gnd 0.008123f
C1878 vdd.n570 gnd 0.010194f
C1879 vdd.n571 gnd 0.010194f
C1880 vdd.n572 gnd 0.010194f
C1881 vdd.n573 gnd 0.010194f
C1882 vdd.n574 gnd 0.010194f
C1883 vdd.n575 gnd 0.008205f
C1884 vdd.n576 gnd 0.008205f
C1885 vdd.n577 gnd 0.010194f
C1886 vdd.n578 gnd 0.010194f
C1887 vdd.n579 gnd 0.008205f
C1888 vdd.n580 gnd 0.010194f
C1889 vdd.n581 gnd 0.010194f
C1890 vdd.n582 gnd 0.010194f
C1891 vdd.n583 gnd 0.010194f
C1892 vdd.n584 gnd 0.010194f
C1893 vdd.n585 gnd 0.008205f
C1894 vdd.n586 gnd 0.008205f
C1895 vdd.n587 gnd 0.010194f
C1896 vdd.n588 gnd 0.010194f
C1897 vdd.n589 gnd 0.008205f
C1898 vdd.n590 gnd 0.010194f
C1899 vdd.n591 gnd 0.010194f
C1900 vdd.n592 gnd 0.010194f
C1901 vdd.n593 gnd 0.010194f
C1902 vdd.n594 gnd 0.010194f
C1903 vdd.n595 gnd 0.008205f
C1904 vdd.n596 gnd 0.008205f
C1905 vdd.n597 gnd 0.010194f
C1906 vdd.n598 gnd 0.010194f
C1907 vdd.n599 gnd 0.008205f
C1908 vdd.n600 gnd 0.010194f
C1909 vdd.n601 gnd 0.010194f
C1910 vdd.n602 gnd 0.010194f
C1911 vdd.n603 gnd 0.010194f
C1912 vdd.n604 gnd 0.010194f
C1913 vdd.n605 gnd 0.008205f
C1914 vdd.n606 gnd 0.008205f
C1915 vdd.n607 gnd 0.010194f
C1916 vdd.n608 gnd 0.010194f
C1917 vdd.n609 gnd 0.008205f
C1918 vdd.n610 gnd 0.010194f
C1919 vdd.n611 gnd 0.010194f
C1920 vdd.n612 gnd 0.010194f
C1921 vdd.n613 gnd 0.010194f
C1922 vdd.n614 gnd 0.010194f
C1923 vdd.n615 gnd 0.008205f
C1924 vdd.n616 gnd 0.010194f
C1925 vdd.n617 gnd 0.008205f
C1926 vdd.n618 gnd 0.004308f
C1927 vdd.n619 gnd 0.010194f
C1928 vdd.n620 gnd 0.010194f
C1929 vdd.n621 gnd 0.008205f
C1930 vdd.n622 gnd 0.010194f
C1931 vdd.n623 gnd 0.008205f
C1932 vdd.n624 gnd 0.010194f
C1933 vdd.n625 gnd 0.008205f
C1934 vdd.n626 gnd 0.010194f
C1935 vdd.n627 gnd 0.008205f
C1936 vdd.n628 gnd 0.010194f
C1937 vdd.n629 gnd 0.008205f
C1938 vdd.n630 gnd 0.010194f
C1939 vdd.n631 gnd 0.008205f
C1940 vdd.n632 gnd 0.010194f
C1941 vdd.n633 gnd 0.567785f
C1942 vdd.t170 gnd 0.520903f
C1943 vdd.n634 gnd 0.010194f
C1944 vdd.n635 gnd 0.008205f
C1945 vdd.n636 gnd 0.010194f
C1946 vdd.n637 gnd 0.008205f
C1947 vdd.n638 gnd 0.010194f
C1948 vdd.t77 gnd 0.520903f
C1949 vdd.n639 gnd 0.010194f
C1950 vdd.n640 gnd 0.008205f
C1951 vdd.n641 gnd 0.010194f
C1952 vdd.n642 gnd 0.008205f
C1953 vdd.n643 gnd 0.010194f
C1954 vdd.t33 gnd 0.520903f
C1955 vdd.n644 gnd 0.651129f
C1956 vdd.n645 gnd 0.010194f
C1957 vdd.n646 gnd 0.008205f
C1958 vdd.n647 gnd 0.010194f
C1959 vdd.n648 gnd 0.008205f
C1960 vdd.n649 gnd 0.010194f
C1961 vdd.t24 gnd 0.520903f
C1962 vdd.n650 gnd 0.010194f
C1963 vdd.n651 gnd 0.008205f
C1964 vdd.n652 gnd 0.010194f
C1965 vdd.n653 gnd 0.008205f
C1966 vdd.n654 gnd 0.010194f
C1967 vdd.n655 gnd 0.724056f
C1968 vdd.n656 gnd 0.864699f
C1969 vdd.t222 gnd 0.520903f
C1970 vdd.n657 gnd 0.010194f
C1971 vdd.n658 gnd 0.008205f
C1972 vdd.n659 gnd 0.010194f
C1973 vdd.n660 gnd 0.008205f
C1974 vdd.n661 gnd 0.010194f
C1975 vdd.n662 gnd 0.546948f
C1976 vdd.n663 gnd 0.010194f
C1977 vdd.n664 gnd 0.008205f
C1978 vdd.n665 gnd 0.010194f
C1979 vdd.n666 gnd 0.008205f
C1980 vdd.n667 gnd 0.010194f
C1981 vdd.t27 gnd 0.520903f
C1982 vdd.t62 gnd 0.520903f
C1983 vdd.n668 gnd 0.010194f
C1984 vdd.n669 gnd 0.008205f
C1985 vdd.n670 gnd 0.010194f
C1986 vdd.n671 gnd 0.008205f
C1987 vdd.n672 gnd 0.010194f
C1988 vdd.t31 gnd 0.520903f
C1989 vdd.n673 gnd 0.010194f
C1990 vdd.n674 gnd 0.008205f
C1991 vdd.n675 gnd 0.010194f
C1992 vdd.n676 gnd 0.008205f
C1993 vdd.n677 gnd 0.010194f
C1994 vdd.n678 gnd 1.04181f
C1995 vdd.n679 gnd 0.849072f
C1996 vdd.n680 gnd 0.010194f
C1997 vdd.n681 gnd 0.008205f
C1998 vdd.n682 gnd 0.024661f
C1999 vdd.n683 gnd 0.00681f
C2000 vdd.n684 gnd 0.024661f
C2001 vdd.t109 gnd 0.520903f
C2002 vdd.n685 gnd 0.024661f
C2003 vdd.n686 gnd 0.00681f
C2004 vdd.n687 gnd 0.008767f
C2005 vdd.t110 gnd 0.125416f
C2006 vdd.t111 gnd 0.134036f
C2007 vdd.t108 gnd 0.163792f
C2008 vdd.n688 gnd 0.209958f
C2009 vdd.n689 gnd 0.176403f
C2010 vdd.n690 gnd 0.012636f
C2011 vdd.n691 gnd 0.010194f
C2012 vdd.n692 gnd 12.303699f
C2013 vdd.n723 gnd 1.43248f
C2014 vdd.n724 gnd 0.010194f
C2015 vdd.n725 gnd 0.010194f
C2016 vdd.n726 gnd 0.025189f
C2017 vdd.n727 gnd 0.008767f
C2018 vdd.n728 gnd 0.010194f
C2019 vdd.n729 gnd 0.008205f
C2020 vdd.n730 gnd 0.006524f
C2021 vdd.n731 gnd 0.042805f
C2022 vdd.n732 gnd 0.008205f
C2023 vdd.n733 gnd 0.010194f
C2024 vdd.n734 gnd 0.010194f
C2025 vdd.n735 gnd 0.010194f
C2026 vdd.n736 gnd 0.010194f
C2027 vdd.n737 gnd 0.010194f
C2028 vdd.n738 gnd 0.010194f
C2029 vdd.n739 gnd 0.010194f
C2030 vdd.n740 gnd 0.010194f
C2031 vdd.n741 gnd 0.010194f
C2032 vdd.n742 gnd 0.010194f
C2033 vdd.n743 gnd 0.010194f
C2034 vdd.n744 gnd 0.010194f
C2035 vdd.n745 gnd 0.010194f
C2036 vdd.n746 gnd 0.010194f
C2037 vdd.n747 gnd 0.006851f
C2038 vdd.n748 gnd 0.010194f
C2039 vdd.n749 gnd 0.010194f
C2040 vdd.n750 gnd 0.010194f
C2041 vdd.n751 gnd 0.010194f
C2042 vdd.n752 gnd 0.010194f
C2043 vdd.n753 gnd 0.010194f
C2044 vdd.n754 gnd 0.010194f
C2045 vdd.n755 gnd 0.010194f
C2046 vdd.n756 gnd 0.010194f
C2047 vdd.n757 gnd 0.010194f
C2048 vdd.n758 gnd 0.010194f
C2049 vdd.n759 gnd 0.010194f
C2050 vdd.n760 gnd 0.010194f
C2051 vdd.n761 gnd 0.010194f
C2052 vdd.n762 gnd 0.010194f
C2053 vdd.n763 gnd 0.010194f
C2054 vdd.n764 gnd 0.010194f
C2055 vdd.n765 gnd 0.010194f
C2056 vdd.n766 gnd 0.010194f
C2057 vdd.n767 gnd 0.008123f
C2058 vdd.t120 gnd 0.125416f
C2059 vdd.t121 gnd 0.134036f
C2060 vdd.t119 gnd 0.163792f
C2061 vdd.n768 gnd 0.209958f
C2062 vdd.n769 gnd 0.176403f
C2063 vdd.n770 gnd 0.010194f
C2064 vdd.n771 gnd 0.010194f
C2065 vdd.n772 gnd 0.010194f
C2066 vdd.n773 gnd 0.010194f
C2067 vdd.n774 gnd 0.010194f
C2068 vdd.n775 gnd 0.010194f
C2069 vdd.n776 gnd 0.010194f
C2070 vdd.n777 gnd 0.010194f
C2071 vdd.n778 gnd 0.010194f
C2072 vdd.n779 gnd 0.010194f
C2073 vdd.n780 gnd 0.010194f
C2074 vdd.n781 gnd 0.010194f
C2075 vdd.n782 gnd 0.010194f
C2076 vdd.n783 gnd 0.006524f
C2077 vdd.n785 gnd 0.006932f
C2078 vdd.n786 gnd 0.006932f
C2079 vdd.n787 gnd 0.006932f
C2080 vdd.n788 gnd 0.006932f
C2081 vdd.n789 gnd 0.006932f
C2082 vdd.n790 gnd 0.006932f
C2083 vdd.n792 gnd 0.006932f
C2084 vdd.n793 gnd 0.006932f
C2085 vdd.n795 gnd 0.006932f
C2086 vdd.n796 gnd 0.005046f
C2087 vdd.n798 gnd 0.006932f
C2088 vdd.t86 gnd 0.280125f
C2089 vdd.t85 gnd 0.286743f
C2090 vdd.t83 gnd 0.182877f
C2091 vdd.n799 gnd 0.098835f
C2092 vdd.n800 gnd 0.056062f
C2093 vdd.n801 gnd 0.009907f
C2094 vdd.n802 gnd 0.01574f
C2095 vdd.n804 gnd 0.006932f
C2096 vdd.n805 gnd 0.708428f
C2097 vdd.n806 gnd 0.014843f
C2098 vdd.n807 gnd 0.014843f
C2099 vdd.n808 gnd 0.006932f
C2100 vdd.n809 gnd 0.01574f
C2101 vdd.n810 gnd 0.006932f
C2102 vdd.n811 gnd 0.006932f
C2103 vdd.n812 gnd 0.006932f
C2104 vdd.n813 gnd 0.006932f
C2105 vdd.n814 gnd 0.006932f
C2106 vdd.n816 gnd 0.006932f
C2107 vdd.n817 gnd 0.006932f
C2108 vdd.n819 gnd 0.006932f
C2109 vdd.n820 gnd 0.006932f
C2110 vdd.n822 gnd 0.006932f
C2111 vdd.n823 gnd 0.006932f
C2112 vdd.n825 gnd 0.006932f
C2113 vdd.n826 gnd 0.006932f
C2114 vdd.n828 gnd 0.006932f
C2115 vdd.n829 gnd 0.006932f
C2116 vdd.n831 gnd 0.006932f
C2117 vdd.t107 gnd 0.280125f
C2118 vdd.t106 gnd 0.286743f
C2119 vdd.t105 gnd 0.182877f
C2120 vdd.n832 gnd 0.098835f
C2121 vdd.n833 gnd 0.056062f
C2122 vdd.n834 gnd 0.006932f
C2123 vdd.n836 gnd 0.006932f
C2124 vdd.n837 gnd 0.006932f
C2125 vdd.t84 gnd 0.354214f
C2126 vdd.n838 gnd 0.006932f
C2127 vdd.n839 gnd 0.006932f
C2128 vdd.n840 gnd 0.006932f
C2129 vdd.n841 gnd 0.006932f
C2130 vdd.n842 gnd 0.006932f
C2131 vdd.n843 gnd 0.708428f
C2132 vdd.n844 gnd 0.006932f
C2133 vdd.n845 gnd 0.006932f
C2134 vdd.n846 gnd 0.557367f
C2135 vdd.n847 gnd 0.006932f
C2136 vdd.n848 gnd 0.006932f
C2137 vdd.n849 gnd 0.006932f
C2138 vdd.n850 gnd 0.006932f
C2139 vdd.n851 gnd 0.708428f
C2140 vdd.n852 gnd 0.006932f
C2141 vdd.n853 gnd 0.006932f
C2142 vdd.n854 gnd 0.006932f
C2143 vdd.n855 gnd 0.006932f
C2144 vdd.n856 gnd 0.006932f
C2145 vdd.t252 gnd 0.354214f
C2146 vdd.n857 gnd 0.006932f
C2147 vdd.n858 gnd 0.006932f
C2148 vdd.n859 gnd 0.006932f
C2149 vdd.n860 gnd 0.006932f
C2150 vdd.n861 gnd 0.006932f
C2151 vdd.t267 gnd 0.354214f
C2152 vdd.n862 gnd 0.006932f
C2153 vdd.n863 gnd 0.006932f
C2154 vdd.n864 gnd 0.682383f
C2155 vdd.n865 gnd 0.006932f
C2156 vdd.n866 gnd 0.006932f
C2157 vdd.n867 gnd 0.006932f
C2158 vdd.t266 gnd 0.354214f
C2159 vdd.n868 gnd 0.006932f
C2160 vdd.n869 gnd 0.006932f
C2161 vdd.n870 gnd 0.526112f
C2162 vdd.n871 gnd 0.006932f
C2163 vdd.n872 gnd 0.006932f
C2164 vdd.n873 gnd 0.006932f
C2165 vdd.n874 gnd 0.494858f
C2166 vdd.n875 gnd 0.006932f
C2167 vdd.n876 gnd 0.006932f
C2168 vdd.n877 gnd 0.369841f
C2169 vdd.n878 gnd 0.006932f
C2170 vdd.n879 gnd 0.006932f
C2171 vdd.n880 gnd 0.006932f
C2172 vdd.n881 gnd 0.651129f
C2173 vdd.n882 gnd 0.006932f
C2174 vdd.n883 gnd 0.006932f
C2175 vdd.t273 gnd 0.354214f
C2176 vdd.n884 gnd 0.006932f
C2177 vdd.n885 gnd 0.006932f
C2178 vdd.n886 gnd 0.006932f
C2179 vdd.n887 gnd 0.708428f
C2180 vdd.n888 gnd 0.006932f
C2181 vdd.n889 gnd 0.006932f
C2182 vdd.t274 gnd 0.354214f
C2183 vdd.n890 gnd 0.006932f
C2184 vdd.n891 gnd 0.006932f
C2185 vdd.n892 gnd 0.006932f
C2186 vdd.t246 gnd 0.354214f
C2187 vdd.n893 gnd 0.006932f
C2188 vdd.n894 gnd 0.006932f
C2189 vdd.n895 gnd 0.006932f
C2190 vdd.t114 gnd 0.286743f
C2191 vdd.t112 gnd 0.182877f
C2192 vdd.t115 gnd 0.286743f
C2193 vdd.n896 gnd 0.161161f
C2194 vdd.n897 gnd 0.020081f
C2195 vdd.n898 gnd 0.006932f
C2196 vdd.t113 gnd 0.255243f
C2197 vdd.n899 gnd 0.006932f
C2198 vdd.n900 gnd 0.006932f
C2199 vdd.n901 gnd 0.609457f
C2200 vdd.n902 gnd 0.006932f
C2201 vdd.n903 gnd 0.006932f
C2202 vdd.n904 gnd 0.006932f
C2203 vdd.n905 gnd 0.411514f
C2204 vdd.n906 gnd 0.006932f
C2205 vdd.n907 gnd 0.006932f
C2206 vdd.t247 gnd 0.145853f
C2207 vdd.n908 gnd 0.453186f
C2208 vdd.n909 gnd 0.006932f
C2209 vdd.n910 gnd 0.006932f
C2210 vdd.n911 gnd 0.006932f
C2211 vdd.n912 gnd 0.567785f
C2212 vdd.n913 gnd 0.006932f
C2213 vdd.n914 gnd 0.006932f
C2214 vdd.t258 gnd 0.354214f
C2215 vdd.n915 gnd 0.006932f
C2216 vdd.n916 gnd 0.006932f
C2217 vdd.n917 gnd 0.006932f
C2218 vdd.t254 gnd 0.354214f
C2219 vdd.n918 gnd 0.006932f
C2220 vdd.n919 gnd 0.006932f
C2221 vdd.t277 gnd 0.354214f
C2222 vdd.n920 gnd 0.006932f
C2223 vdd.n921 gnd 0.006932f
C2224 vdd.n922 gnd 0.006932f
C2225 vdd.t236 gnd 0.239616f
C2226 vdd.n923 gnd 0.006932f
C2227 vdd.n924 gnd 0.006932f
C2228 vdd.n925 gnd 0.625084f
C2229 vdd.n926 gnd 0.006932f
C2230 vdd.n927 gnd 0.006932f
C2231 vdd.n928 gnd 0.006932f
C2232 vdd.t278 gnd 0.354214f
C2233 vdd.n929 gnd 0.006932f
C2234 vdd.n930 gnd 0.006932f
C2235 vdd.t290 gnd 0.338587f
C2236 vdd.n931 gnd 0.468813f
C2237 vdd.n932 gnd 0.006932f
C2238 vdd.n933 gnd 0.006932f
C2239 vdd.n934 gnd 0.006932f
C2240 vdd.t242 gnd 0.354214f
C2241 vdd.n935 gnd 0.006932f
C2242 vdd.n936 gnd 0.006932f
C2243 vdd.t282 gnd 0.354214f
C2244 vdd.n937 gnd 0.006932f
C2245 vdd.n938 gnd 0.006932f
C2246 vdd.n939 gnd 0.006932f
C2247 vdd.n940 gnd 0.708428f
C2248 vdd.n941 gnd 0.006932f
C2249 vdd.n942 gnd 0.006932f
C2250 vdd.t262 gnd 0.354214f
C2251 vdd.n943 gnd 0.006932f
C2252 vdd.n944 gnd 0.006932f
C2253 vdd.n945 gnd 0.006932f
C2254 vdd.n946 gnd 0.489649f
C2255 vdd.n947 gnd 0.006932f
C2256 vdd.n948 gnd 0.006932f
C2257 vdd.n949 gnd 0.006932f
C2258 vdd.n950 gnd 0.006932f
C2259 vdd.n951 gnd 0.006932f
C2260 vdd.t136 gnd 0.354214f
C2261 vdd.n952 gnd 0.006932f
C2262 vdd.n953 gnd 0.006932f
C2263 vdd.t244 gnd 0.354214f
C2264 vdd.n954 gnd 0.006932f
C2265 vdd.n955 gnd 0.014843f
C2266 vdd.n956 gnd 0.014843f
C2267 vdd.n957 gnd 0.802191f
C2268 vdd.n958 gnd 0.006932f
C2269 vdd.n959 gnd 0.006932f
C2270 vdd.t271 gnd 0.354214f
C2271 vdd.n960 gnd 0.014843f
C2272 vdd.n961 gnd 0.006932f
C2273 vdd.n962 gnd 0.006932f
C2274 vdd.t284 gnd 0.604248f
C2275 vdd.n980 gnd 0.01574f
C2276 vdd.n998 gnd 0.014843f
C2277 vdd.n999 gnd 0.006932f
C2278 vdd.n1000 gnd 0.014843f
C2279 vdd.t152 gnd 0.280125f
C2280 vdd.t151 gnd 0.286743f
C2281 vdd.t150 gnd 0.182877f
C2282 vdd.n1001 gnd 0.098835f
C2283 vdd.n1002 gnd 0.056062f
C2284 vdd.n1003 gnd 0.01574f
C2285 vdd.n1004 gnd 0.006932f
C2286 vdd.n1005 gnd 0.416723f
C2287 vdd.n1006 gnd 0.014843f
C2288 vdd.n1007 gnd 0.006932f
C2289 vdd.n1008 gnd 0.01574f
C2290 vdd.n1009 gnd 0.006932f
C2291 vdd.t131 gnd 0.280125f
C2292 vdd.t130 gnd 0.286743f
C2293 vdd.t128 gnd 0.182877f
C2294 vdd.n1010 gnd 0.098835f
C2295 vdd.n1011 gnd 0.056062f
C2296 vdd.n1012 gnd 0.009907f
C2297 vdd.n1013 gnd 0.006932f
C2298 vdd.n1014 gnd 0.006932f
C2299 vdd.t129 gnd 0.354214f
C2300 vdd.n1015 gnd 0.006932f
C2301 vdd.t286 gnd 0.354214f
C2302 vdd.n1016 gnd 0.006932f
C2303 vdd.n1017 gnd 0.006932f
C2304 vdd.n1018 gnd 0.006932f
C2305 vdd.n1019 gnd 0.006932f
C2306 vdd.n1020 gnd 0.006932f
C2307 vdd.n1021 gnd 0.708428f
C2308 vdd.n1022 gnd 0.006932f
C2309 vdd.n1023 gnd 0.006932f
C2310 vdd.t256 gnd 0.354214f
C2311 vdd.n1024 gnd 0.006932f
C2312 vdd.n1025 gnd 0.006932f
C2313 vdd.n1026 gnd 0.006932f
C2314 vdd.n1027 gnd 0.006932f
C2315 vdd.n1028 gnd 0.510485f
C2316 vdd.n1029 gnd 0.006932f
C2317 vdd.n1030 gnd 0.006932f
C2318 vdd.n1031 gnd 0.006932f
C2319 vdd.n1032 gnd 0.006932f
C2320 vdd.n1033 gnd 0.006932f
C2321 vdd.t237 gnd 0.354214f
C2322 vdd.n1034 gnd 0.006932f
C2323 vdd.n1035 gnd 0.006932f
C2324 vdd.t275 gnd 0.354214f
C2325 vdd.n1036 gnd 0.006932f
C2326 vdd.n1037 gnd 0.006932f
C2327 vdd.n1038 gnd 0.006932f
C2328 vdd.t259 gnd 0.354214f
C2329 vdd.n1039 gnd 0.006932f
C2330 vdd.n1040 gnd 0.006932f
C2331 vdd.t238 gnd 0.354214f
C2332 vdd.n1041 gnd 0.006932f
C2333 vdd.n1042 gnd 0.006932f
C2334 vdd.n1043 gnd 0.006932f
C2335 vdd.t260 gnd 0.338587f
C2336 vdd.n1044 gnd 0.006932f
C2337 vdd.n1045 gnd 0.006932f
C2338 vdd.n1046 gnd 0.526112f
C2339 vdd.n1047 gnd 0.006932f
C2340 vdd.n1048 gnd 0.006932f
C2341 vdd.n1049 gnd 0.006932f
C2342 vdd.t279 gnd 0.354214f
C2343 vdd.n1050 gnd 0.006932f
C2344 vdd.n1051 gnd 0.006932f
C2345 vdd.t249 gnd 0.239616f
C2346 vdd.n1052 gnd 0.369841f
C2347 vdd.n1053 gnd 0.006932f
C2348 vdd.n1054 gnd 0.006932f
C2349 vdd.n1055 gnd 0.006932f
C2350 vdd.n1056 gnd 0.651129f
C2351 vdd.n1057 gnd 0.006932f
C2352 vdd.n1058 gnd 0.006932f
C2353 vdd.t288 gnd 0.354214f
C2354 vdd.n1059 gnd 0.006932f
C2355 vdd.n1060 gnd 0.006932f
C2356 vdd.n1061 gnd 0.006932f
C2357 vdd.n1062 gnd 0.708428f
C2358 vdd.n1063 gnd 0.006932f
C2359 vdd.n1064 gnd 0.006932f
C2360 vdd.t253 gnd 0.354214f
C2361 vdd.n1065 gnd 0.006932f
C2362 vdd.n1066 gnd 0.006932f
C2363 vdd.n1067 gnd 0.006932f
C2364 vdd.t248 gnd 0.145853f
C2365 vdd.n1068 gnd 0.006932f
C2366 vdd.n1069 gnd 0.006932f
C2367 vdd.n1070 gnd 0.006932f
C2368 vdd.t141 gnd 0.286743f
C2369 vdd.t139 gnd 0.182877f
C2370 vdd.t142 gnd 0.286743f
C2371 vdd.n1071 gnd 0.161161f
C2372 vdd.n1072 gnd 0.006932f
C2373 vdd.n1073 gnd 0.006932f
C2374 vdd.t268 gnd 0.354214f
C2375 vdd.n1074 gnd 0.006932f
C2376 vdd.n1075 gnd 0.006932f
C2377 vdd.t140 gnd 0.255243f
C2378 vdd.n1076 gnd 0.562576f
C2379 vdd.n1077 gnd 0.006932f
C2380 vdd.n1078 gnd 0.006932f
C2381 vdd.n1079 gnd 0.006932f
C2382 vdd.n1080 gnd 0.411514f
C2383 vdd.n1081 gnd 0.006932f
C2384 vdd.n1082 gnd 0.006932f
C2385 vdd.n1083 gnd 0.453186f
C2386 vdd.n1084 gnd 0.006932f
C2387 vdd.n1085 gnd 0.006932f
C2388 vdd.n1086 gnd 0.006932f
C2389 vdd.n1087 gnd 0.567785f
C2390 vdd.n1088 gnd 0.006932f
C2391 vdd.n1089 gnd 0.006932f
C2392 vdd.t250 gnd 0.354214f
C2393 vdd.n1090 gnd 0.006932f
C2394 vdd.n1091 gnd 0.006932f
C2395 vdd.n1092 gnd 0.006932f
C2396 vdd.n1093 gnd 0.708428f
C2397 vdd.n1094 gnd 0.006932f
C2398 vdd.n1095 gnd 0.006932f
C2399 vdd.t251 gnd 0.354214f
C2400 vdd.n1096 gnd 0.006932f
C2401 vdd.n1097 gnd 0.006932f
C2402 vdd.n1098 gnd 0.006932f
C2403 vdd.t289 gnd 0.354214f
C2404 vdd.n1099 gnd 0.006932f
C2405 vdd.n1100 gnd 0.006932f
C2406 vdd.n1101 gnd 0.006932f
C2407 vdd.n1102 gnd 0.006932f
C2408 vdd.n1103 gnd 0.006932f
C2409 vdd.t281 gnd 0.354214f
C2410 vdd.n1104 gnd 0.006932f
C2411 vdd.n1105 gnd 0.006932f
C2412 vdd.n1106 gnd 0.692801f
C2413 vdd.n1107 gnd 0.006932f
C2414 vdd.n1108 gnd 0.006932f
C2415 vdd.n1109 gnd 0.006932f
C2416 vdd.t243 gnd 0.354214f
C2417 vdd.n1110 gnd 0.006932f
C2418 vdd.n1111 gnd 0.006932f
C2419 vdd.n1112 gnd 0.53653f
C2420 vdd.n1113 gnd 0.006932f
C2421 vdd.n1114 gnd 0.006932f
C2422 vdd.n1115 gnd 0.006932f
C2423 vdd.n1116 gnd 0.708428f
C2424 vdd.n1117 gnd 0.006932f
C2425 vdd.n1118 gnd 0.006932f
C2426 vdd.n1119 gnd 0.380259f
C2427 vdd.n1120 gnd 0.006932f
C2428 vdd.n1121 gnd 0.006932f
C2429 vdd.n1122 gnd 0.006932f
C2430 vdd.n1123 gnd 0.708428f
C2431 vdd.n1124 gnd 0.006932f
C2432 vdd.n1125 gnd 0.006932f
C2433 vdd.n1126 gnd 0.006932f
C2434 vdd.n1127 gnd 0.006932f
C2435 vdd.n1128 gnd 0.006932f
C2436 vdd.t88 gnd 0.354214f
C2437 vdd.n1129 gnd 0.006932f
C2438 vdd.n1130 gnd 0.006932f
C2439 vdd.n1131 gnd 0.006932f
C2440 vdd.n1132 gnd 0.014843f
C2441 vdd.n1133 gnd 0.014843f
C2442 vdd.n1134 gnd 0.958462f
C2443 vdd.n1135 gnd 0.006932f
C2444 vdd.n1136 gnd 0.006932f
C2445 vdd.n1137 gnd 0.505276f
C2446 vdd.n1138 gnd 0.014843f
C2447 vdd.n1139 gnd 0.006932f
C2448 vdd.n1140 gnd 0.006932f
C2449 vdd.n1141 gnd 12.7205f
C2450 vdd.n1175 gnd 0.01574f
C2451 vdd.n1176 gnd 0.006932f
C2452 vdd.n1177 gnd 0.006932f
C2453 vdd.n1178 gnd 0.006524f
C2454 vdd.n1181 gnd 0.025189f
C2455 vdd.n1182 gnd 0.00681f
C2456 vdd.n1183 gnd 0.008205f
C2457 vdd.n1185 gnd 0.010194f
C2458 vdd.n1186 gnd 0.010194f
C2459 vdd.n1187 gnd 0.008205f
C2460 vdd.n1189 gnd 0.010194f
C2461 vdd.n1190 gnd 0.010194f
C2462 vdd.n1191 gnd 0.010194f
C2463 vdd.n1192 gnd 0.010194f
C2464 vdd.n1193 gnd 0.010194f
C2465 vdd.n1194 gnd 0.008205f
C2466 vdd.n1196 gnd 0.010194f
C2467 vdd.n1197 gnd 0.010194f
C2468 vdd.n1198 gnd 0.010194f
C2469 vdd.n1199 gnd 0.010194f
C2470 vdd.n1200 gnd 0.010194f
C2471 vdd.n1201 gnd 0.008205f
C2472 vdd.n1203 gnd 0.010194f
C2473 vdd.n1204 gnd 0.010194f
C2474 vdd.n1205 gnd 0.010194f
C2475 vdd.n1206 gnd 0.010194f
C2476 vdd.n1207 gnd 0.006851f
C2477 vdd.t101 gnd 0.125416f
C2478 vdd.t100 gnd 0.134036f
C2479 vdd.t99 gnd 0.163792f
C2480 vdd.n1208 gnd 0.209958f
C2481 vdd.n1209 gnd 0.176403f
C2482 vdd.n1211 gnd 0.010194f
C2483 vdd.n1212 gnd 0.010194f
C2484 vdd.n1213 gnd 0.008205f
C2485 vdd.n1214 gnd 0.010194f
C2486 vdd.n1216 gnd 0.010194f
C2487 vdd.n1217 gnd 0.010194f
C2488 vdd.n1218 gnd 0.010194f
C2489 vdd.n1219 gnd 0.010194f
C2490 vdd.n1220 gnd 0.008205f
C2491 vdd.n1222 gnd 0.010194f
C2492 vdd.n1223 gnd 0.010194f
C2493 vdd.n1224 gnd 0.010194f
C2494 vdd.n1225 gnd 0.010194f
C2495 vdd.n1226 gnd 0.010194f
C2496 vdd.n1227 gnd 0.008205f
C2497 vdd.n1229 gnd 0.010194f
C2498 vdd.n1230 gnd 0.010194f
C2499 vdd.n1231 gnd 0.010194f
C2500 vdd.n1232 gnd 0.010194f
C2501 vdd.n1233 gnd 0.010194f
C2502 vdd.n1234 gnd 0.008205f
C2503 vdd.n1236 gnd 0.010194f
C2504 vdd.n1237 gnd 0.010194f
C2505 vdd.n1238 gnd 0.010194f
C2506 vdd.n1239 gnd 0.010194f
C2507 vdd.n1240 gnd 0.010194f
C2508 vdd.n1241 gnd 0.008205f
C2509 vdd.n1243 gnd 0.010194f
C2510 vdd.n1244 gnd 0.010194f
C2511 vdd.n1245 gnd 0.010194f
C2512 vdd.n1246 gnd 0.010194f
C2513 vdd.n1247 gnd 0.008123f
C2514 vdd.t94 gnd 0.125416f
C2515 vdd.t93 gnd 0.134036f
C2516 vdd.t91 gnd 0.163792f
C2517 vdd.n1248 gnd 0.209958f
C2518 vdd.n1249 gnd 0.176403f
C2519 vdd.n1251 gnd 0.010194f
C2520 vdd.n1252 gnd 0.010194f
C2521 vdd.n1253 gnd 0.008205f
C2522 vdd.n1254 gnd 0.010194f
C2523 vdd.n1256 gnd 0.010194f
C2524 vdd.n1257 gnd 0.010194f
C2525 vdd.n1258 gnd 0.010194f
C2526 vdd.n1259 gnd 0.010194f
C2527 vdd.n1260 gnd 0.008205f
C2528 vdd.n1262 gnd 0.010194f
C2529 vdd.n1263 gnd 0.010194f
C2530 vdd.n1264 gnd 0.010194f
C2531 vdd.n1265 gnd 0.010194f
C2532 vdd.n1266 gnd 0.010194f
C2533 vdd.n1267 gnd 0.008205f
C2534 vdd.n1269 gnd 0.010194f
C2535 vdd.n1270 gnd 0.010194f
C2536 vdd.n1271 gnd 0.010194f
C2537 vdd.n1272 gnd 0.010194f
C2538 vdd.n1273 gnd 0.010194f
C2539 vdd.n1274 gnd 0.008205f
C2540 vdd.n1276 gnd 0.010194f
C2541 vdd.n1277 gnd 0.010194f
C2542 vdd.n1278 gnd 0.006524f
C2543 vdd.n1279 gnd 0.008205f
C2544 vdd.n1280 gnd 0.01574f
C2545 vdd.n1281 gnd 0.01574f
C2546 vdd.n1282 gnd 0.006932f
C2547 vdd.n1283 gnd 0.006932f
C2548 vdd.n1284 gnd 0.006932f
C2549 vdd.n1285 gnd 0.006932f
C2550 vdd.n1286 gnd 0.006932f
C2551 vdd.n1287 gnd 0.006932f
C2552 vdd.n1288 gnd 0.006932f
C2553 vdd.n1289 gnd 0.006932f
C2554 vdd.n1290 gnd 0.006932f
C2555 vdd.n1291 gnd 0.006932f
C2556 vdd.n1292 gnd 0.006932f
C2557 vdd.n1293 gnd 0.006932f
C2558 vdd.n1294 gnd 0.006932f
C2559 vdd.n1295 gnd 0.006932f
C2560 vdd.n1296 gnd 0.006932f
C2561 vdd.n1297 gnd 0.006932f
C2562 vdd.n1298 gnd 0.006932f
C2563 vdd.n1299 gnd 0.006932f
C2564 vdd.n1300 gnd 0.006932f
C2565 vdd.n1301 gnd 0.006932f
C2566 vdd.n1302 gnd 0.006932f
C2567 vdd.n1303 gnd 0.006932f
C2568 vdd.n1304 gnd 0.006932f
C2569 vdd.n1305 gnd 0.006932f
C2570 vdd.n1306 gnd 0.006932f
C2571 vdd.n1307 gnd 0.006932f
C2572 vdd.n1308 gnd 0.006932f
C2573 vdd.n1309 gnd 0.006932f
C2574 vdd.n1310 gnd 0.006932f
C2575 vdd.n1311 gnd 0.006932f
C2576 vdd.n1312 gnd 0.006932f
C2577 vdd.n1313 gnd 0.006932f
C2578 vdd.n1314 gnd 0.006932f
C2579 vdd.t89 gnd 0.280125f
C2580 vdd.t90 gnd 0.286743f
C2581 vdd.t87 gnd 0.182877f
C2582 vdd.n1315 gnd 0.098835f
C2583 vdd.n1316 gnd 0.056062f
C2584 vdd.n1317 gnd 0.009907f
C2585 vdd.n1318 gnd 0.006932f
C2586 vdd.t126 gnd 0.280125f
C2587 vdd.t127 gnd 0.286743f
C2588 vdd.t125 gnd 0.182877f
C2589 vdd.n1319 gnd 0.098835f
C2590 vdd.n1320 gnd 0.056062f
C2591 vdd.n1321 gnd 0.006932f
C2592 vdd.n1322 gnd 0.006932f
C2593 vdd.n1323 gnd 0.006932f
C2594 vdd.n1324 gnd 0.006932f
C2595 vdd.n1325 gnd 0.006932f
C2596 vdd.n1326 gnd 0.006932f
C2597 vdd.n1327 gnd 0.006932f
C2598 vdd.n1328 gnd 0.006932f
C2599 vdd.n1329 gnd 0.006932f
C2600 vdd.n1330 gnd 0.006932f
C2601 vdd.n1331 gnd 0.006932f
C2602 vdd.n1332 gnd 0.006932f
C2603 vdd.n1333 gnd 0.006932f
C2604 vdd.n1334 gnd 0.006932f
C2605 vdd.n1335 gnd 0.006932f
C2606 vdd.n1336 gnd 0.006932f
C2607 vdd.n1337 gnd 0.006932f
C2608 vdd.n1338 gnd 0.006932f
C2609 vdd.n1339 gnd 0.006932f
C2610 vdd.n1340 gnd 0.006932f
C2611 vdd.n1341 gnd 0.006932f
C2612 vdd.n1342 gnd 0.006932f
C2613 vdd.n1343 gnd 0.006932f
C2614 vdd.n1344 gnd 0.006932f
C2615 vdd.n1345 gnd 0.006932f
C2616 vdd.n1346 gnd 0.006932f
C2617 vdd.n1347 gnd 0.005046f
C2618 vdd.n1348 gnd 0.009907f
C2619 vdd.n1349 gnd 0.005352f
C2620 vdd.n1350 gnd 0.006932f
C2621 vdd.n1351 gnd 0.006932f
C2622 vdd.n1352 gnd 0.006932f
C2623 vdd.n1353 gnd 0.01574f
C2624 vdd.n1354 gnd 0.01574f
C2625 vdd.n1355 gnd 0.014843f
C2626 vdd.n1356 gnd 0.014843f
C2627 vdd.n1357 gnd 0.006932f
C2628 vdd.n1358 gnd 0.006932f
C2629 vdd.n1359 gnd 0.006932f
C2630 vdd.n1360 gnd 0.006932f
C2631 vdd.n1361 gnd 0.006932f
C2632 vdd.n1362 gnd 0.006932f
C2633 vdd.n1363 gnd 0.006932f
C2634 vdd.n1364 gnd 0.006932f
C2635 vdd.n1365 gnd 0.006932f
C2636 vdd.n1366 gnd 0.006932f
C2637 vdd.n1367 gnd 0.006932f
C2638 vdd.n1368 gnd 0.006932f
C2639 vdd.n1369 gnd 0.006932f
C2640 vdd.n1370 gnd 0.006932f
C2641 vdd.n1371 gnd 0.006932f
C2642 vdd.n1372 gnd 0.006932f
C2643 vdd.n1373 gnd 0.006932f
C2644 vdd.n1374 gnd 0.006932f
C2645 vdd.n1375 gnd 0.006932f
C2646 vdd.n1376 gnd 0.006932f
C2647 vdd.n1377 gnd 0.006932f
C2648 vdd.n1378 gnd 0.006932f
C2649 vdd.n1379 gnd 0.006932f
C2650 vdd.n1380 gnd 0.006932f
C2651 vdd.n1381 gnd 0.006932f
C2652 vdd.n1382 gnd 0.006932f
C2653 vdd.n1383 gnd 0.006932f
C2654 vdd.n1384 gnd 0.006932f
C2655 vdd.n1385 gnd 0.006932f
C2656 vdd.n1386 gnd 0.006932f
C2657 vdd.n1387 gnd 0.006932f
C2658 vdd.n1388 gnd 0.006932f
C2659 vdd.n1389 gnd 0.006932f
C2660 vdd.n1390 gnd 0.006932f
C2661 vdd.n1391 gnd 0.006932f
C2662 vdd.n1392 gnd 0.006932f
C2663 vdd.n1393 gnd 0.006932f
C2664 vdd.n1394 gnd 0.006932f
C2665 vdd.n1395 gnd 0.006932f
C2666 vdd.n1396 gnd 0.006932f
C2667 vdd.n1397 gnd 0.006932f
C2668 vdd.n1398 gnd 0.006932f
C2669 vdd.n1399 gnd 0.421932f
C2670 vdd.n1400 gnd 0.006932f
C2671 vdd.n1401 gnd 0.006932f
C2672 vdd.n1402 gnd 0.006932f
C2673 vdd.n1403 gnd 0.006932f
C2674 vdd.n1404 gnd 0.006932f
C2675 vdd.n1405 gnd 0.006932f
C2676 vdd.n1406 gnd 0.006932f
C2677 vdd.n1407 gnd 0.006932f
C2678 vdd.n1408 gnd 0.006932f
C2679 vdd.n1409 gnd 0.006932f
C2680 vdd.n1410 gnd 0.006932f
C2681 vdd.n1411 gnd 0.006932f
C2682 vdd.n1412 gnd 0.006932f
C2683 vdd.n1413 gnd 0.006932f
C2684 vdd.n1414 gnd 0.006932f
C2685 vdd.n1415 gnd 0.006932f
C2686 vdd.n1416 gnd 0.006932f
C2687 vdd.n1417 gnd 0.006932f
C2688 vdd.n1418 gnd 0.006932f
C2689 vdd.n1419 gnd 0.006932f
C2690 vdd.n1420 gnd 0.006932f
C2691 vdd.n1421 gnd 0.006932f
C2692 vdd.n1422 gnd 0.006932f
C2693 vdd.n1423 gnd 0.006932f
C2694 vdd.n1424 gnd 0.006932f
C2695 vdd.n1425 gnd 0.640711f
C2696 vdd.n1426 gnd 0.006932f
C2697 vdd.n1427 gnd 0.006932f
C2698 vdd.n1428 gnd 0.006932f
C2699 vdd.n1429 gnd 0.006932f
C2700 vdd.n1430 gnd 0.006932f
C2701 vdd.n1431 gnd 0.006932f
C2702 vdd.n1432 gnd 0.006932f
C2703 vdd.n1433 gnd 0.006932f
C2704 vdd.n1434 gnd 0.006932f
C2705 vdd.n1435 gnd 0.006932f
C2706 vdd.n1436 gnd 0.006932f
C2707 vdd.n1437 gnd 0.223988f
C2708 vdd.n1438 gnd 0.006932f
C2709 vdd.n1439 gnd 0.006932f
C2710 vdd.n1440 gnd 0.006932f
C2711 vdd.n1441 gnd 0.006932f
C2712 vdd.n1442 gnd 0.006932f
C2713 vdd.n1443 gnd 0.006932f
C2714 vdd.n1444 gnd 0.006932f
C2715 vdd.n1445 gnd 0.006932f
C2716 vdd.n1446 gnd 0.006932f
C2717 vdd.n1447 gnd 0.006932f
C2718 vdd.n1448 gnd 0.006932f
C2719 vdd.n1449 gnd 0.006932f
C2720 vdd.n1450 gnd 0.006932f
C2721 vdd.n1451 gnd 0.006932f
C2722 vdd.n1452 gnd 0.006932f
C2723 vdd.n1453 gnd 0.006932f
C2724 vdd.n1454 gnd 0.006932f
C2725 vdd.n1455 gnd 0.006932f
C2726 vdd.n1456 gnd 0.006932f
C2727 vdd.n1457 gnd 0.006932f
C2728 vdd.n1458 gnd 0.006932f
C2729 vdd.n1459 gnd 0.006932f
C2730 vdd.n1460 gnd 0.006932f
C2731 vdd.n1461 gnd 0.006932f
C2732 vdd.n1462 gnd 0.006932f
C2733 vdd.n1463 gnd 0.006932f
C2734 vdd.n1464 gnd 0.006932f
C2735 vdd.n1465 gnd 0.006932f
C2736 vdd.n1466 gnd 0.006932f
C2737 vdd.n1467 gnd 0.006932f
C2738 vdd.n1468 gnd 0.006932f
C2739 vdd.n1469 gnd 0.006932f
C2740 vdd.n1470 gnd 0.006932f
C2741 vdd.n1471 gnd 0.006932f
C2742 vdd.n1472 gnd 0.006932f
C2743 vdd.n1473 gnd 0.006932f
C2744 vdd.n1474 gnd 0.006932f
C2745 vdd.n1475 gnd 0.006932f
C2746 vdd.n1476 gnd 0.006932f
C2747 vdd.n1477 gnd 0.006932f
C2748 vdd.n1478 gnd 0.006932f
C2749 vdd.n1479 gnd 0.006932f
C2750 vdd.n1480 gnd 0.014843f
C2751 vdd.n1481 gnd 0.014843f
C2752 vdd.n1482 gnd 0.01574f
C2753 vdd.n1483 gnd 0.006932f
C2754 vdd.n1484 gnd 0.006932f
C2755 vdd.n1485 gnd 0.005352f
C2756 vdd.n1486 gnd 0.006932f
C2757 vdd.n1487 gnd 0.006932f
C2758 vdd.n1488 gnd 0.005046f
C2759 vdd.n1489 gnd 0.006932f
C2760 vdd.n1490 gnd 0.006932f
C2761 vdd.n1491 gnd 0.006932f
C2762 vdd.n1492 gnd 0.006932f
C2763 vdd.n1493 gnd 0.006932f
C2764 vdd.n1494 gnd 0.006932f
C2765 vdd.n1495 gnd 0.006932f
C2766 vdd.n1496 gnd 0.006932f
C2767 vdd.n1497 gnd 0.006932f
C2768 vdd.n1498 gnd 0.006932f
C2769 vdd.n1499 gnd 0.006932f
C2770 vdd.n1500 gnd 0.006932f
C2771 vdd.n1501 gnd 0.006932f
C2772 vdd.n1502 gnd 0.006932f
C2773 vdd.n1503 gnd 0.006932f
C2774 vdd.n1504 gnd 0.006932f
C2775 vdd.n1505 gnd 0.006932f
C2776 vdd.n1506 gnd 0.006932f
C2777 vdd.n1507 gnd 0.006932f
C2778 vdd.n1508 gnd 0.006932f
C2779 vdd.n1509 gnd 0.006932f
C2780 vdd.n1510 gnd 0.006932f
C2781 vdd.n1511 gnd 0.006932f
C2782 vdd.n1512 gnd 0.006932f
C2783 vdd.n1513 gnd 0.006932f
C2784 vdd.n1514 gnd 0.006932f
C2785 vdd.n1515 gnd 0.046698f
C2786 vdd.n1517 gnd 0.025189f
C2787 vdd.n1518 gnd 0.008205f
C2788 vdd.n1520 gnd 0.010194f
C2789 vdd.n1521 gnd 0.008205f
C2790 vdd.n1522 gnd 0.010194f
C2791 vdd.n1524 gnd 0.010194f
C2792 vdd.n1525 gnd 0.010194f
C2793 vdd.n1527 gnd 0.010194f
C2794 vdd.n1528 gnd 0.00681f
C2795 vdd.t92 gnd 0.520903f
C2796 vdd.n1529 gnd 0.010194f
C2797 vdd.n1530 gnd 0.025189f
C2798 vdd.n1531 gnd 0.008205f
C2799 vdd.n1532 gnd 0.010194f
C2800 vdd.n1533 gnd 0.008205f
C2801 vdd.n1534 gnd 0.010194f
C2802 vdd.n1535 gnd 1.04181f
C2803 vdd.n1536 gnd 0.010194f
C2804 vdd.n1537 gnd 0.008205f
C2805 vdd.n1538 gnd 0.008205f
C2806 vdd.n1539 gnd 0.010194f
C2807 vdd.n1540 gnd 0.008205f
C2808 vdd.n1541 gnd 0.010194f
C2809 vdd.t47 gnd 0.520903f
C2810 vdd.n1542 gnd 0.010194f
C2811 vdd.n1543 gnd 0.008205f
C2812 vdd.n1544 gnd 0.010194f
C2813 vdd.n1545 gnd 0.008205f
C2814 vdd.n1546 gnd 0.010194f
C2815 vdd.t35 gnd 0.520903f
C2816 vdd.n1547 gnd 0.010194f
C2817 vdd.n1548 gnd 0.008205f
C2818 vdd.n1549 gnd 0.010194f
C2819 vdd.n1550 gnd 0.008205f
C2820 vdd.n1551 gnd 0.010194f
C2821 vdd.n1552 gnd 0.838654f
C2822 vdd.n1553 gnd 0.864699f
C2823 vdd.t193 gnd 0.520903f
C2824 vdd.n1554 gnd 0.010194f
C2825 vdd.n1555 gnd 0.008205f
C2826 vdd.n1556 gnd 0.010194f
C2827 vdd.n1557 gnd 0.008205f
C2828 vdd.n1558 gnd 0.010194f
C2829 vdd.n1559 gnd 0.661547f
C2830 vdd.n1560 gnd 0.010194f
C2831 vdd.n1561 gnd 0.008205f
C2832 vdd.n1562 gnd 0.010194f
C2833 vdd.n1563 gnd 0.008205f
C2834 vdd.n1564 gnd 0.010194f
C2835 vdd.t43 gnd 0.520903f
C2836 vdd.t56 gnd 0.520903f
C2837 vdd.n1565 gnd 0.010194f
C2838 vdd.n1566 gnd 0.008205f
C2839 vdd.n1567 gnd 0.010194f
C2840 vdd.n1568 gnd 0.008205f
C2841 vdd.n1569 gnd 0.010194f
C2842 vdd.t161 gnd 0.520903f
C2843 vdd.n1570 gnd 0.010194f
C2844 vdd.n1571 gnd 0.008205f
C2845 vdd.n1572 gnd 0.010194f
C2846 vdd.n1573 gnd 0.008205f
C2847 vdd.n1574 gnd 0.010194f
C2848 vdd.t167 gnd 0.520903f
C2849 vdd.n1575 gnd 0.734474f
C2850 vdd.n1576 gnd 0.010194f
C2851 vdd.n1577 gnd 0.008205f
C2852 vdd.n1578 gnd 0.010194f
C2853 vdd.n1579 gnd 0.008205f
C2854 vdd.n1580 gnd 0.010194f
C2855 vdd.n1581 gnd 0.817818f
C2856 vdd.n1582 gnd 0.010194f
C2857 vdd.n1583 gnd 0.008205f
C2858 vdd.n1584 gnd 0.010194f
C2859 vdd.n1585 gnd 0.008205f
C2860 vdd.n1586 gnd 0.010194f
C2861 vdd.n1587 gnd 0.640711f
C2862 vdd.t72 gnd 0.520903f
C2863 vdd.n1588 gnd 0.010194f
C2864 vdd.n1589 gnd 0.008205f
C2865 vdd.n1590 gnd 0.010194f
C2866 vdd.n1591 gnd 0.008205f
C2867 vdd.n1592 gnd 0.010194f
C2868 vdd.t179 gnd 0.520903f
C2869 vdd.n1593 gnd 0.010194f
C2870 vdd.n1594 gnd 0.008205f
C2871 vdd.n1595 gnd 0.010194f
C2872 vdd.n1596 gnd 0.008205f
C2873 vdd.n1597 gnd 0.010194f
C2874 vdd.t49 gnd 0.520903f
C2875 vdd.n1598 gnd 0.578203f
C2876 vdd.n1599 gnd 0.010194f
C2877 vdd.n1600 gnd 0.008205f
C2878 vdd.n1601 gnd 0.010194f
C2879 vdd.n1602 gnd 0.008205f
C2880 vdd.n1603 gnd 0.010194f
C2881 vdd.t203 gnd 0.520903f
C2882 vdd.n1604 gnd 0.010194f
C2883 vdd.n1605 gnd 0.008205f
C2884 vdd.n1606 gnd 0.010194f
C2885 vdd.n1607 gnd 0.008205f
C2886 vdd.n1608 gnd 0.010194f
C2887 vdd.n1609 gnd 0.796982f
C2888 vdd.n1610 gnd 0.864699f
C2889 vdd.t163 gnd 0.520903f
C2890 vdd.n1611 gnd 0.010194f
C2891 vdd.n1612 gnd 0.008205f
C2892 vdd.n1613 gnd 0.010194f
C2893 vdd.n1614 gnd 0.008205f
C2894 vdd.n1615 gnd 0.010194f
C2895 vdd.n1616 gnd 0.619875f
C2896 vdd.n1617 gnd 0.010194f
C2897 vdd.n1618 gnd 0.008205f
C2898 vdd.n1619 gnd 0.010194f
C2899 vdd.n1620 gnd 0.008205f
C2900 vdd.n1621 gnd 0.010194f
C2901 vdd.t58 gnd 0.520903f
C2902 vdd.t79 gnd 0.520903f
C2903 vdd.n1622 gnd 0.010194f
C2904 vdd.n1623 gnd 0.008205f
C2905 vdd.n1624 gnd 0.010194f
C2906 vdd.n1625 gnd 0.008205f
C2907 vdd.n1626 gnd 0.010194f
C2908 vdd.t45 gnd 0.520903f
C2909 vdd.n1627 gnd 0.010194f
C2910 vdd.n1628 gnd 0.008205f
C2911 vdd.n1629 gnd 0.010194f
C2912 vdd.n1630 gnd 0.008205f
C2913 vdd.n1631 gnd 0.010194f
C2914 vdd.t37 gnd 0.520903f
C2915 vdd.n1632 gnd 0.776146f
C2916 vdd.n1633 gnd 0.010194f
C2917 vdd.n1634 gnd 0.008205f
C2918 vdd.n1635 gnd 0.010194f
C2919 vdd.n1636 gnd 0.008205f
C2920 vdd.n1637 gnd 0.010194f
C2921 vdd.n1638 gnd 1.04181f
C2922 vdd.n1639 gnd 0.010194f
C2923 vdd.n1640 gnd 0.008205f
C2924 vdd.n1641 gnd 0.024661f
C2925 vdd.n1642 gnd 0.00681f
C2926 vdd.n1643 gnd 0.024661f
C2927 vdd.t147 gnd 0.520903f
C2928 vdd.n1644 gnd 0.024661f
C2929 vdd.n1645 gnd 0.00681f
C2930 vdd.n1646 gnd 0.010194f
C2931 vdd.n1647 gnd 0.008205f
C2932 vdd.n1648 gnd 0.010194f
C2933 vdd.n1679 gnd 0.025189f
C2934 vdd.n1680 gnd 1.53666f
C2935 vdd.n1681 gnd 0.010194f
C2936 vdd.n1682 gnd 0.008205f
C2937 vdd.n1683 gnd 0.010194f
C2938 vdd.n1684 gnd 0.010194f
C2939 vdd.n1685 gnd 0.010194f
C2940 vdd.n1686 gnd 0.010194f
C2941 vdd.n1687 gnd 0.010194f
C2942 vdd.n1688 gnd 0.008205f
C2943 vdd.n1689 gnd 0.010194f
C2944 vdd.n1690 gnd 0.010194f
C2945 vdd.n1691 gnd 0.010194f
C2946 vdd.n1692 gnd 0.010194f
C2947 vdd.n1693 gnd 0.010194f
C2948 vdd.n1694 gnd 0.008205f
C2949 vdd.n1695 gnd 0.010194f
C2950 vdd.n1696 gnd 0.010194f
C2951 vdd.n1697 gnd 0.010194f
C2952 vdd.n1698 gnd 0.010194f
C2953 vdd.n1699 gnd 0.010194f
C2954 vdd.n1700 gnd 0.008205f
C2955 vdd.n1701 gnd 0.010194f
C2956 vdd.n1702 gnd 0.010194f
C2957 vdd.n1703 gnd 0.010194f
C2958 vdd.n1704 gnd 0.010194f
C2959 vdd.n1705 gnd 0.010194f
C2960 vdd.t157 gnd 0.125416f
C2961 vdd.t158 gnd 0.134036f
C2962 vdd.t156 gnd 0.163792f
C2963 vdd.n1706 gnd 0.209958f
C2964 vdd.n1707 gnd 0.177224f
C2965 vdd.n1708 gnd 0.017559f
C2966 vdd.n1709 gnd 0.010194f
C2967 vdd.n1710 gnd 0.010194f
C2968 vdd.n1711 gnd 0.010194f
C2969 vdd.n1712 gnd 0.010194f
C2970 vdd.n1713 gnd 0.010194f
C2971 vdd.n1714 gnd 0.008205f
C2972 vdd.n1715 gnd 0.010194f
C2973 vdd.n1716 gnd 0.010194f
C2974 vdd.n1717 gnd 0.010194f
C2975 vdd.n1718 gnd 0.010194f
C2976 vdd.n1719 gnd 0.010194f
C2977 vdd.n1720 gnd 0.008205f
C2978 vdd.n1721 gnd 0.010194f
C2979 vdd.n1722 gnd 0.010194f
C2980 vdd.n1723 gnd 0.010194f
C2981 vdd.n1724 gnd 0.010194f
C2982 vdd.n1725 gnd 0.010194f
C2983 vdd.n1726 gnd 0.008205f
C2984 vdd.n1727 gnd 0.010194f
C2985 vdd.n1728 gnd 0.010194f
C2986 vdd.n1729 gnd 0.010194f
C2987 vdd.n1730 gnd 0.010194f
C2988 vdd.n1731 gnd 0.010194f
C2989 vdd.n1732 gnd 0.008205f
C2990 vdd.n1733 gnd 0.010194f
C2991 vdd.n1734 gnd 0.010194f
C2992 vdd.n1735 gnd 0.010194f
C2993 vdd.n1736 gnd 0.010194f
C2994 vdd.n1737 gnd 0.010194f
C2995 vdd.n1738 gnd 0.008205f
C2996 vdd.n1739 gnd 0.010194f
C2997 vdd.n1740 gnd 0.010194f
C2998 vdd.n1741 gnd 0.010194f
C2999 vdd.n1742 gnd 0.010194f
C3000 vdd.n1743 gnd 0.008205f
C3001 vdd.n1744 gnd 0.010194f
C3002 vdd.n1745 gnd 0.010194f
C3003 vdd.n1746 gnd 0.010194f
C3004 vdd.n1747 gnd 0.010194f
C3005 vdd.n1748 gnd 0.010194f
C3006 vdd.n1749 gnd 0.008205f
C3007 vdd.n1750 gnd 0.010194f
C3008 vdd.n1751 gnd 0.010194f
C3009 vdd.n1752 gnd 0.010194f
C3010 vdd.n1753 gnd 0.010194f
C3011 vdd.n1754 gnd 0.010194f
C3012 vdd.n1755 gnd 0.008205f
C3013 vdd.n1756 gnd 0.010194f
C3014 vdd.n1757 gnd 0.010194f
C3015 vdd.n1758 gnd 0.010194f
C3016 vdd.n1759 gnd 0.010194f
C3017 vdd.n1760 gnd 0.010194f
C3018 vdd.n1761 gnd 0.008205f
C3019 vdd.n1762 gnd 0.010194f
C3020 vdd.n1763 gnd 0.010194f
C3021 vdd.n1764 gnd 0.010194f
C3022 vdd.n1765 gnd 0.010194f
C3023 vdd.n1766 gnd 0.010194f
C3024 vdd.n1767 gnd 0.008205f
C3025 vdd.n1768 gnd 0.010194f
C3026 vdd.n1769 gnd 0.010194f
C3027 vdd.n1770 gnd 0.010194f
C3028 vdd.n1771 gnd 0.010194f
C3029 vdd.t154 gnd 0.125416f
C3030 vdd.t155 gnd 0.134036f
C3031 vdd.t153 gnd 0.163792f
C3032 vdd.n1772 gnd 0.209958f
C3033 vdd.n1773 gnd 0.177224f
C3034 vdd.n1774 gnd 0.013457f
C3035 vdd.n1775 gnd 0.003897f
C3036 vdd.n1776 gnd 0.025189f
C3037 vdd.n1777 gnd 0.010194f
C3038 vdd.n1778 gnd 0.004308f
C3039 vdd.n1779 gnd 0.008205f
C3040 vdd.n1780 gnd 0.008205f
C3041 vdd.n1781 gnd 0.010194f
C3042 vdd.n1782 gnd 0.010194f
C3043 vdd.n1783 gnd 0.010194f
C3044 vdd.n1784 gnd 0.008205f
C3045 vdd.n1785 gnd 0.008205f
C3046 vdd.n1786 gnd 0.008205f
C3047 vdd.n1787 gnd 0.010194f
C3048 vdd.n1788 gnd 0.010194f
C3049 vdd.n1789 gnd 0.010194f
C3050 vdd.n1790 gnd 0.008205f
C3051 vdd.n1791 gnd 0.008205f
C3052 vdd.n1792 gnd 0.008205f
C3053 vdd.n1793 gnd 0.010194f
C3054 vdd.n1794 gnd 0.010194f
C3055 vdd.n1795 gnd 0.010194f
C3056 vdd.n1796 gnd 0.008205f
C3057 vdd.n1797 gnd 0.008205f
C3058 vdd.n1798 gnd 0.008205f
C3059 vdd.n1799 gnd 0.010194f
C3060 vdd.n1800 gnd 0.010194f
C3061 vdd.n1801 gnd 0.010194f
C3062 vdd.n1802 gnd 0.008205f
C3063 vdd.n1803 gnd 0.008205f
C3064 vdd.n1804 gnd 0.008205f
C3065 vdd.n1805 gnd 0.010194f
C3066 vdd.n1806 gnd 0.010194f
C3067 vdd.n1807 gnd 0.010194f
C3068 vdd.n1808 gnd 0.008123f
C3069 vdd.n1809 gnd 0.010194f
C3070 vdd.t148 gnd 0.125416f
C3071 vdd.t149 gnd 0.134036f
C3072 vdd.t146 gnd 0.163792f
C3073 vdd.n1810 gnd 0.209958f
C3074 vdd.n1811 gnd 0.177224f
C3075 vdd.n1812 gnd 0.017559f
C3076 vdd.n1813 gnd 0.00558f
C3077 vdd.n1814 gnd 0.010194f
C3078 vdd.n1815 gnd 0.010194f
C3079 vdd.n1816 gnd 0.010194f
C3080 vdd.n1817 gnd 0.008205f
C3081 vdd.n1818 gnd 0.008205f
C3082 vdd.n1819 gnd 0.008205f
C3083 vdd.n1820 gnd 0.010194f
C3084 vdd.n1821 gnd 0.010194f
C3085 vdd.n1822 gnd 0.010194f
C3086 vdd.n1823 gnd 0.008205f
C3087 vdd.n1824 gnd 0.008205f
C3088 vdd.n1825 gnd 0.008205f
C3089 vdd.n1826 gnd 0.010194f
C3090 vdd.n1827 gnd 0.010194f
C3091 vdd.n1828 gnd 0.010194f
C3092 vdd.n1829 gnd 0.008205f
C3093 vdd.n1830 gnd 0.008205f
C3094 vdd.n1831 gnd 0.008205f
C3095 vdd.n1832 gnd 0.010194f
C3096 vdd.n1833 gnd 0.010194f
C3097 vdd.n1834 gnd 0.010194f
C3098 vdd.n1835 gnd 0.008205f
C3099 vdd.n1836 gnd 0.008205f
C3100 vdd.n1837 gnd 0.008205f
C3101 vdd.n1838 gnd 0.010194f
C3102 vdd.n1839 gnd 0.010194f
C3103 vdd.n1840 gnd 0.010194f
C3104 vdd.n1841 gnd 0.008205f
C3105 vdd.n1842 gnd 0.008205f
C3106 vdd.n1843 gnd 0.006851f
C3107 vdd.n1844 gnd 0.010194f
C3108 vdd.n1845 gnd 0.010194f
C3109 vdd.n1846 gnd 0.010194f
C3110 vdd.n1847 gnd 0.006851f
C3111 vdd.n1848 gnd 0.008205f
C3112 vdd.n1849 gnd 0.008205f
C3113 vdd.n1850 gnd 0.010194f
C3114 vdd.n1851 gnd 0.010194f
C3115 vdd.n1852 gnd 0.010194f
C3116 vdd.n1853 gnd 0.008205f
C3117 vdd.n1854 gnd 0.008205f
C3118 vdd.n1855 gnd 0.008205f
C3119 vdd.n1856 gnd 0.010194f
C3120 vdd.n1857 gnd 0.010194f
C3121 vdd.n1858 gnd 0.010194f
C3122 vdd.n1859 gnd 0.008205f
C3123 vdd.n1860 gnd 0.008205f
C3124 vdd.n1861 gnd 0.008205f
C3125 vdd.n1862 gnd 0.010194f
C3126 vdd.n1863 gnd 0.010194f
C3127 vdd.n1864 gnd 0.010194f
C3128 vdd.n1865 gnd 0.008205f
C3129 vdd.n1866 gnd 0.008205f
C3130 vdd.n1867 gnd 0.008205f
C3131 vdd.n1868 gnd 0.010194f
C3132 vdd.n1869 gnd 0.010194f
C3133 vdd.n1870 gnd 0.010194f
C3134 vdd.n1871 gnd 0.008205f
C3135 vdd.n1872 gnd 0.010194f
C3136 vdd.n1873 gnd 2.46908f
C3137 vdd.n1875 gnd 0.025189f
C3138 vdd.n1876 gnd 0.00681f
C3139 vdd.n1877 gnd 0.025189f
C3140 vdd.n1878 gnd 0.024661f
C3141 vdd.n1879 gnd 0.010194f
C3142 vdd.n1880 gnd 0.008205f
C3143 vdd.n1881 gnd 0.010194f
C3144 vdd.n1882 gnd 0.526112f
C3145 vdd.n1883 gnd 0.010194f
C3146 vdd.n1884 gnd 0.008205f
C3147 vdd.n1885 gnd 0.010194f
C3148 vdd.n1886 gnd 0.010194f
C3149 vdd.n1887 gnd 0.010194f
C3150 vdd.n1888 gnd 0.008205f
C3151 vdd.n1889 gnd 0.010194f
C3152 vdd.n1890 gnd 0.953253f
C3153 vdd.n1891 gnd 1.04181f
C3154 vdd.n1892 gnd 0.010194f
C3155 vdd.n1893 gnd 0.008205f
C3156 vdd.n1894 gnd 0.010194f
C3157 vdd.n1895 gnd 0.010194f
C3158 vdd.n1896 gnd 0.010194f
C3159 vdd.n1897 gnd 0.008205f
C3160 vdd.n1898 gnd 0.010194f
C3161 vdd.n1899 gnd 0.609457f
C3162 vdd.n1900 gnd 0.010194f
C3163 vdd.n1901 gnd 0.008205f
C3164 vdd.n1902 gnd 0.010194f
C3165 vdd.n1903 gnd 0.010194f
C3166 vdd.n1904 gnd 0.010194f
C3167 vdd.n1905 gnd 0.008205f
C3168 vdd.n1906 gnd 0.010194f
C3169 vdd.n1907 gnd 0.599039f
C3170 vdd.n1908 gnd 0.786564f
C3171 vdd.n1909 gnd 0.010194f
C3172 vdd.n1910 gnd 0.008205f
C3173 vdd.n1911 gnd 0.010194f
C3174 vdd.n1912 gnd 0.010194f
C3175 vdd.n1913 gnd 0.010194f
C3176 vdd.n1914 gnd 0.008205f
C3177 vdd.n1915 gnd 0.010194f
C3178 vdd.n1916 gnd 0.864699f
C3179 vdd.n1917 gnd 0.010194f
C3180 vdd.n1918 gnd 0.008205f
C3181 vdd.n1919 gnd 0.010194f
C3182 vdd.n1920 gnd 0.010194f
C3183 vdd.n1921 gnd 0.010194f
C3184 vdd.n1922 gnd 0.008205f
C3185 vdd.n1923 gnd 0.010194f
C3186 vdd.t4 gnd 0.520903f
C3187 vdd.n1924 gnd 0.765728f
C3188 vdd.n1925 gnd 0.010194f
C3189 vdd.n1926 gnd 0.008205f
C3190 vdd.n1927 gnd 0.010194f
C3191 vdd.n1928 gnd 0.010194f
C3192 vdd.n1929 gnd 0.010194f
C3193 vdd.n1930 gnd 0.008205f
C3194 vdd.n1931 gnd 0.010194f
C3195 vdd.n1932 gnd 0.588621f
C3196 vdd.n1933 gnd 0.010194f
C3197 vdd.n1934 gnd 0.008205f
C3198 vdd.n1935 gnd 0.010194f
C3199 vdd.n1936 gnd 0.010194f
C3200 vdd.n1937 gnd 0.010194f
C3201 vdd.n1938 gnd 0.008205f
C3202 vdd.n1939 gnd 0.010194f
C3203 vdd.n1940 gnd 0.75531f
C3204 vdd.n1941 gnd 0.630293f
C3205 vdd.n1942 gnd 0.010194f
C3206 vdd.n1943 gnd 0.008205f
C3207 vdd.n1944 gnd 0.010194f
C3208 vdd.n1945 gnd 0.010194f
C3209 vdd.n1946 gnd 0.010194f
C3210 vdd.n1947 gnd 0.008205f
C3211 vdd.n1948 gnd 0.010194f
C3212 vdd.n1949 gnd 0.8074f
C3213 vdd.n1950 gnd 0.010194f
C3214 vdd.n1951 gnd 0.008205f
C3215 vdd.n1952 gnd 0.010194f
C3216 vdd.n1953 gnd 0.010194f
C3217 vdd.n1954 gnd 0.010194f
C3218 vdd.n1955 gnd 0.008205f
C3219 vdd.n1956 gnd 0.010194f
C3220 vdd.t75 gnd 0.520903f
C3221 vdd.n1957 gnd 0.864699f
C3222 vdd.n1958 gnd 0.010194f
C3223 vdd.n1959 gnd 0.008205f
C3224 vdd.n1960 gnd 0.010194f
C3225 vdd.n1961 gnd 0.007835f
C3226 vdd.n1962 gnd 0.005595f
C3227 vdd.n1963 gnd 0.005192f
C3228 vdd.n1964 gnd 0.002872f
C3229 vdd.n1965 gnd 0.006594f
C3230 vdd.n1966 gnd 0.00279f
C3231 vdd.n1967 gnd 0.002954f
C3232 vdd.n1968 gnd 0.005192f
C3233 vdd.n1969 gnd 0.00279f
C3234 vdd.n1970 gnd 0.006594f
C3235 vdd.n1971 gnd 0.002954f
C3236 vdd.n1972 gnd 0.005192f
C3237 vdd.n1973 gnd 0.00279f
C3238 vdd.n1974 gnd 0.004945f
C3239 vdd.n1975 gnd 0.00496f
C3240 vdd.t48 gnd 0.014167f
C3241 vdd.n1976 gnd 0.03152f
C3242 vdd.n1977 gnd 0.16404f
C3243 vdd.n1978 gnd 0.00279f
C3244 vdd.n1979 gnd 0.002954f
C3245 vdd.n1980 gnd 0.006594f
C3246 vdd.n1981 gnd 0.006594f
C3247 vdd.n1982 gnd 0.002954f
C3248 vdd.n1983 gnd 0.00279f
C3249 vdd.n1984 gnd 0.005192f
C3250 vdd.n1985 gnd 0.005192f
C3251 vdd.n1986 gnd 0.00279f
C3252 vdd.n1987 gnd 0.002954f
C3253 vdd.n1988 gnd 0.006594f
C3254 vdd.n1989 gnd 0.006594f
C3255 vdd.n1990 gnd 0.002954f
C3256 vdd.n1991 gnd 0.00279f
C3257 vdd.n1992 gnd 0.005192f
C3258 vdd.n1993 gnd 0.005192f
C3259 vdd.n1994 gnd 0.00279f
C3260 vdd.n1995 gnd 0.002954f
C3261 vdd.n1996 gnd 0.006594f
C3262 vdd.n1997 gnd 0.006594f
C3263 vdd.n1998 gnd 0.01559f
C3264 vdd.n1999 gnd 0.002872f
C3265 vdd.n2000 gnd 0.00279f
C3266 vdd.n2001 gnd 0.013419f
C3267 vdd.n2002 gnd 0.009368f
C3268 vdd.t293 gnd 0.032821f
C3269 vdd.t68 gnd 0.032821f
C3270 vdd.n2003 gnd 0.225566f
C3271 vdd.n2004 gnd 0.177373f
C3272 vdd.t221 gnd 0.032821f
C3273 vdd.t214 gnd 0.032821f
C3274 vdd.n2005 gnd 0.225566f
C3275 vdd.n2006 gnd 0.143139f
C3276 vdd.t192 gnd 0.032821f
C3277 vdd.t44 gnd 0.032821f
C3278 vdd.n2007 gnd 0.225566f
C3279 vdd.n2008 gnd 0.143139f
C3280 vdd.t208 gnd 0.032821f
C3281 vdd.t168 gnd 0.032821f
C3282 vdd.n2009 gnd 0.225566f
C3283 vdd.n2010 gnd 0.143139f
C3284 vdd.t76 gnd 0.032821f
C3285 vdd.t169 gnd 0.032821f
C3286 vdd.n2011 gnd 0.225566f
C3287 vdd.n2012 gnd 0.143139f
C3288 vdd.t229 gnd 0.032821f
C3289 vdd.t189 gnd 0.032821f
C3290 vdd.n2013 gnd 0.225566f
C3291 vdd.n2014 gnd 0.143139f
C3292 vdd.t220 gnd 0.032821f
C3293 vdd.t305 gnd 0.032821f
C3294 vdd.n2015 gnd 0.225566f
C3295 vdd.n2016 gnd 0.143139f
C3296 vdd.t80 gnd 0.032821f
C3297 vdd.t5 gnd 0.032821f
C3298 vdd.n2017 gnd 0.225566f
C3299 vdd.n2018 gnd 0.143139f
C3300 vdd.t206 gnd 0.032821f
C3301 vdd.t166 gnd 0.032821f
C3302 vdd.n2019 gnd 0.225566f
C3303 vdd.n2020 gnd 0.143139f
C3304 vdd.n2021 gnd 0.005595f
C3305 vdd.n2022 gnd 0.005192f
C3306 vdd.n2023 gnd 0.002872f
C3307 vdd.n2024 gnd 0.006594f
C3308 vdd.n2025 gnd 0.00279f
C3309 vdd.n2026 gnd 0.002954f
C3310 vdd.n2027 gnd 0.005192f
C3311 vdd.n2028 gnd 0.00279f
C3312 vdd.n2029 gnd 0.006594f
C3313 vdd.n2030 gnd 0.002954f
C3314 vdd.n2031 gnd 0.005192f
C3315 vdd.n2032 gnd 0.00279f
C3316 vdd.n2033 gnd 0.004945f
C3317 vdd.n2034 gnd 0.00496f
C3318 vdd.t225 gnd 0.014167f
C3319 vdd.n2035 gnd 0.03152f
C3320 vdd.n2036 gnd 0.16404f
C3321 vdd.n2037 gnd 0.00279f
C3322 vdd.n2038 gnd 0.002954f
C3323 vdd.n2039 gnd 0.006594f
C3324 vdd.n2040 gnd 0.006594f
C3325 vdd.n2041 gnd 0.002954f
C3326 vdd.n2042 gnd 0.00279f
C3327 vdd.n2043 gnd 0.005192f
C3328 vdd.n2044 gnd 0.005192f
C3329 vdd.n2045 gnd 0.00279f
C3330 vdd.n2046 gnd 0.002954f
C3331 vdd.n2047 gnd 0.006594f
C3332 vdd.n2048 gnd 0.006594f
C3333 vdd.n2049 gnd 0.002954f
C3334 vdd.n2050 gnd 0.00279f
C3335 vdd.n2051 gnd 0.005192f
C3336 vdd.n2052 gnd 0.005192f
C3337 vdd.n2053 gnd 0.00279f
C3338 vdd.n2054 gnd 0.002954f
C3339 vdd.n2055 gnd 0.006594f
C3340 vdd.n2056 gnd 0.006594f
C3341 vdd.n2057 gnd 0.01559f
C3342 vdd.n2058 gnd 0.002872f
C3343 vdd.n2059 gnd 0.00279f
C3344 vdd.n2060 gnd 0.013419f
C3345 vdd.n2061 gnd 0.009074f
C3346 vdd.n2062 gnd 0.106496f
C3347 vdd.n2063 gnd 0.005595f
C3348 vdd.n2064 gnd 0.005192f
C3349 vdd.n2065 gnd 0.002872f
C3350 vdd.n2066 gnd 0.006594f
C3351 vdd.n2067 gnd 0.00279f
C3352 vdd.n2068 gnd 0.002954f
C3353 vdd.n2069 gnd 0.005192f
C3354 vdd.n2070 gnd 0.00279f
C3355 vdd.n2071 gnd 0.006594f
C3356 vdd.n2072 gnd 0.002954f
C3357 vdd.n2073 gnd 0.005192f
C3358 vdd.n2074 gnd 0.00279f
C3359 vdd.n2075 gnd 0.004945f
C3360 vdd.n2076 gnd 0.00496f
C3361 vdd.t165 gnd 0.014167f
C3362 vdd.n2077 gnd 0.03152f
C3363 vdd.n2078 gnd 0.16404f
C3364 vdd.n2079 gnd 0.00279f
C3365 vdd.n2080 gnd 0.002954f
C3366 vdd.n2081 gnd 0.006594f
C3367 vdd.n2082 gnd 0.006594f
C3368 vdd.n2083 gnd 0.002954f
C3369 vdd.n2084 gnd 0.00279f
C3370 vdd.n2085 gnd 0.005192f
C3371 vdd.n2086 gnd 0.005192f
C3372 vdd.n2087 gnd 0.00279f
C3373 vdd.n2088 gnd 0.002954f
C3374 vdd.n2089 gnd 0.006594f
C3375 vdd.n2090 gnd 0.006594f
C3376 vdd.n2091 gnd 0.002954f
C3377 vdd.n2092 gnd 0.00279f
C3378 vdd.n2093 gnd 0.005192f
C3379 vdd.n2094 gnd 0.005192f
C3380 vdd.n2095 gnd 0.00279f
C3381 vdd.n2096 gnd 0.002954f
C3382 vdd.n2097 gnd 0.006594f
C3383 vdd.n2098 gnd 0.006594f
C3384 vdd.n2099 gnd 0.01559f
C3385 vdd.n2100 gnd 0.002872f
C3386 vdd.n2101 gnd 0.00279f
C3387 vdd.n2102 gnd 0.013419f
C3388 vdd.n2103 gnd 0.009368f
C3389 vdd.t194 gnd 0.032821f
C3390 vdd.t183 gnd 0.032821f
C3391 vdd.n2104 gnd 0.225566f
C3392 vdd.n2105 gnd 0.177373f
C3393 vdd.t209 gnd 0.032821f
C3394 vdd.t175 gnd 0.032821f
C3395 vdd.n2106 gnd 0.225566f
C3396 vdd.n2107 gnd 0.143139f
C3397 vdd.t162 gnd 0.032821f
C3398 vdd.t61 gnd 0.032821f
C3399 vdd.n2108 gnd 0.225566f
C3400 vdd.n2109 gnd 0.143139f
C3401 vdd.t212 gnd 0.032821f
C3402 vdd.t176 gnd 0.032821f
C3403 vdd.n2110 gnd 0.225566f
C3404 vdd.n2111 gnd 0.143139f
C3405 vdd.t196 gnd 0.032821f
C3406 vdd.t73 gnd 0.032821f
C3407 vdd.n2112 gnd 0.225566f
C3408 vdd.n2113 gnd 0.143139f
C3409 vdd.t50 gnd 0.032821f
C3410 vdd.t301 gnd 0.032821f
C3411 vdd.n2114 gnd 0.225566f
C3412 vdd.n2115 gnd 0.143139f
C3413 vdd.t164 gnd 0.032821f
C3414 vdd.t204 gnd 0.032821f
C3415 vdd.n2116 gnd 0.225566f
C3416 vdd.n2117 gnd 0.143139f
C3417 vdd.t228 gnd 0.032821f
C3418 vdd.t182 gnd 0.032821f
C3419 vdd.n2118 gnd 0.225566f
C3420 vdd.n2119 gnd 0.143139f
C3421 vdd.t46 gnd 0.032821f
C3422 vdd.t296 gnd 0.032821f
C3423 vdd.n2120 gnd 0.225566f
C3424 vdd.n2121 gnd 0.143139f
C3425 vdd.n2122 gnd 0.005595f
C3426 vdd.n2123 gnd 0.005192f
C3427 vdd.n2124 gnd 0.002872f
C3428 vdd.n2125 gnd 0.006594f
C3429 vdd.n2126 gnd 0.00279f
C3430 vdd.n2127 gnd 0.002954f
C3431 vdd.n2128 gnd 0.005192f
C3432 vdd.n2129 gnd 0.00279f
C3433 vdd.n2130 gnd 0.006594f
C3434 vdd.n2131 gnd 0.002954f
C3435 vdd.n2132 gnd 0.005192f
C3436 vdd.n2133 gnd 0.00279f
C3437 vdd.n2134 gnd 0.004945f
C3438 vdd.n2135 gnd 0.00496f
C3439 vdd.t60 gnd 0.014167f
C3440 vdd.n2136 gnd 0.03152f
C3441 vdd.n2137 gnd 0.16404f
C3442 vdd.n2138 gnd 0.00279f
C3443 vdd.n2139 gnd 0.002954f
C3444 vdd.n2140 gnd 0.006594f
C3445 vdd.n2141 gnd 0.006594f
C3446 vdd.n2142 gnd 0.002954f
C3447 vdd.n2143 gnd 0.00279f
C3448 vdd.n2144 gnd 0.005192f
C3449 vdd.n2145 gnd 0.005192f
C3450 vdd.n2146 gnd 0.00279f
C3451 vdd.n2147 gnd 0.002954f
C3452 vdd.n2148 gnd 0.006594f
C3453 vdd.n2149 gnd 0.006594f
C3454 vdd.n2150 gnd 0.002954f
C3455 vdd.n2151 gnd 0.00279f
C3456 vdd.n2152 gnd 0.005192f
C3457 vdd.n2153 gnd 0.005192f
C3458 vdd.n2154 gnd 0.00279f
C3459 vdd.n2155 gnd 0.002954f
C3460 vdd.n2156 gnd 0.006594f
C3461 vdd.n2157 gnd 0.006594f
C3462 vdd.n2158 gnd 0.01559f
C3463 vdd.n2159 gnd 0.002872f
C3464 vdd.n2160 gnd 0.00279f
C3465 vdd.n2161 gnd 0.013419f
C3466 vdd.n2162 gnd 0.009074f
C3467 vdd.n2163 gnd 0.063354f
C3468 vdd.n2164 gnd 0.228283f
C3469 vdd.n2165 gnd 0.005595f
C3470 vdd.n2166 gnd 0.005192f
C3471 vdd.n2167 gnd 0.002872f
C3472 vdd.n2168 gnd 0.006594f
C3473 vdd.n2169 gnd 0.00279f
C3474 vdd.n2170 gnd 0.002954f
C3475 vdd.n2171 gnd 0.005192f
C3476 vdd.n2172 gnd 0.00279f
C3477 vdd.n2173 gnd 0.006594f
C3478 vdd.n2174 gnd 0.002954f
C3479 vdd.n2175 gnd 0.005192f
C3480 vdd.n2176 gnd 0.00279f
C3481 vdd.n2177 gnd 0.004945f
C3482 vdd.n2178 gnd 0.00496f
C3483 vdd.t211 gnd 0.014167f
C3484 vdd.n2179 gnd 0.03152f
C3485 vdd.n2180 gnd 0.16404f
C3486 vdd.n2181 gnd 0.00279f
C3487 vdd.n2182 gnd 0.002954f
C3488 vdd.n2183 gnd 0.006594f
C3489 vdd.n2184 gnd 0.006594f
C3490 vdd.n2185 gnd 0.002954f
C3491 vdd.n2186 gnd 0.00279f
C3492 vdd.n2187 gnd 0.005192f
C3493 vdd.n2188 gnd 0.005192f
C3494 vdd.n2189 gnd 0.00279f
C3495 vdd.n2190 gnd 0.002954f
C3496 vdd.n2191 gnd 0.006594f
C3497 vdd.n2192 gnd 0.006594f
C3498 vdd.n2193 gnd 0.002954f
C3499 vdd.n2194 gnd 0.00279f
C3500 vdd.n2195 gnd 0.005192f
C3501 vdd.n2196 gnd 0.005192f
C3502 vdd.n2197 gnd 0.00279f
C3503 vdd.n2198 gnd 0.002954f
C3504 vdd.n2199 gnd 0.006594f
C3505 vdd.n2200 gnd 0.006594f
C3506 vdd.n2201 gnd 0.01559f
C3507 vdd.n2202 gnd 0.002872f
C3508 vdd.n2203 gnd 0.00279f
C3509 vdd.n2204 gnd 0.013419f
C3510 vdd.n2205 gnd 0.009368f
C3511 vdd.t298 gnd 0.032821f
C3512 vdd.t36 gnd 0.032821f
C3513 vdd.n2206 gnd 0.225566f
C3514 vdd.n2207 gnd 0.177373f
C3515 vdd.t57 gnd 0.032821f
C3516 vdd.t306 gnd 0.032821f
C3517 vdd.n2208 gnd 0.225566f
C3518 vdd.n2209 gnd 0.143139f
C3519 vdd.t213 gnd 0.032821f
C3520 vdd.t215 gnd 0.032821f
C3521 vdd.n2210 gnd 0.225566f
C3522 vdd.n2211 gnd 0.143139f
C3523 vdd.t304 gnd 0.032821f
C3524 vdd.t307 gnd 0.032821f
C3525 vdd.n2212 gnd 0.225566f
C3526 vdd.n2213 gnd 0.143139f
C3527 vdd.t198 gnd 0.032821f
C3528 vdd.t224 gnd 0.032821f
C3529 vdd.n2214 gnd 0.225566f
C3530 vdd.n2215 gnd 0.143139f
C3531 vdd.t201 gnd 0.032821f
C3532 vdd.t180 gnd 0.032821f
C3533 vdd.n2216 gnd 0.225566f
C3534 vdd.n2217 gnd 0.143139f
C3535 vdd.t303 gnd 0.032821f
C3536 vdd.t219 gnd 0.032821f
C3537 vdd.n2218 gnd 0.225566f
C3538 vdd.n2219 gnd 0.143139f
C3539 vdd.t217 gnd 0.032821f
C3540 vdd.t299 gnd 0.032821f
C3541 vdd.n2220 gnd 0.225566f
C3542 vdd.n2221 gnd 0.143139f
C3543 vdd.t216 gnd 0.032821f
C3544 vdd.t59 gnd 0.032821f
C3545 vdd.n2222 gnd 0.225566f
C3546 vdd.n2223 gnd 0.143139f
C3547 vdd.n2224 gnd 0.005595f
C3548 vdd.n2225 gnd 0.005192f
C3549 vdd.n2226 gnd 0.002872f
C3550 vdd.n2227 gnd 0.006594f
C3551 vdd.n2228 gnd 0.00279f
C3552 vdd.n2229 gnd 0.002954f
C3553 vdd.n2230 gnd 0.005192f
C3554 vdd.n2231 gnd 0.00279f
C3555 vdd.n2232 gnd 0.006594f
C3556 vdd.n2233 gnd 0.002954f
C3557 vdd.n2234 gnd 0.005192f
C3558 vdd.n2235 gnd 0.00279f
C3559 vdd.n2236 gnd 0.004945f
C3560 vdd.n2237 gnd 0.00496f
C3561 vdd.t38 gnd 0.014167f
C3562 vdd.n2238 gnd 0.03152f
C3563 vdd.n2239 gnd 0.16404f
C3564 vdd.n2240 gnd 0.00279f
C3565 vdd.n2241 gnd 0.002954f
C3566 vdd.n2242 gnd 0.006594f
C3567 vdd.n2243 gnd 0.006594f
C3568 vdd.n2244 gnd 0.002954f
C3569 vdd.n2245 gnd 0.00279f
C3570 vdd.n2246 gnd 0.005192f
C3571 vdd.n2247 gnd 0.005192f
C3572 vdd.n2248 gnd 0.00279f
C3573 vdd.n2249 gnd 0.002954f
C3574 vdd.n2250 gnd 0.006594f
C3575 vdd.n2251 gnd 0.006594f
C3576 vdd.n2252 gnd 0.002954f
C3577 vdd.n2253 gnd 0.00279f
C3578 vdd.n2254 gnd 0.005192f
C3579 vdd.n2255 gnd 0.005192f
C3580 vdd.n2256 gnd 0.00279f
C3581 vdd.n2257 gnd 0.002954f
C3582 vdd.n2258 gnd 0.006594f
C3583 vdd.n2259 gnd 0.006594f
C3584 vdd.n2260 gnd 0.01559f
C3585 vdd.n2261 gnd 0.002872f
C3586 vdd.n2262 gnd 0.00279f
C3587 vdd.n2263 gnd 0.013419f
C3588 vdd.n2264 gnd 0.009074f
C3589 vdd.n2265 gnd 0.063354f
C3590 vdd.n2266 gnd 0.261334f
C3591 vdd.n2267 gnd 2.98821f
C3592 vdd.n2268 gnd 0.601297f
C3593 vdd.n2269 gnd 0.007835f
C3594 vdd.n2270 gnd 0.008205f
C3595 vdd.n2271 gnd 0.010194f
C3596 vdd.n2272 gnd 0.744892f
C3597 vdd.n2273 gnd 0.010194f
C3598 vdd.n2274 gnd 0.008205f
C3599 vdd.n2275 gnd 0.010194f
C3600 vdd.n2276 gnd 0.010194f
C3601 vdd.n2277 gnd 0.010194f
C3602 vdd.n2278 gnd 0.008205f
C3603 vdd.n2279 gnd 0.010194f
C3604 vdd.n2280 gnd 0.864699f
C3605 vdd.t207 gnd 0.520903f
C3606 vdd.n2281 gnd 0.567785f
C3607 vdd.n2282 gnd 0.010194f
C3608 vdd.n2283 gnd 0.008205f
C3609 vdd.n2284 gnd 0.010194f
C3610 vdd.n2285 gnd 0.010194f
C3611 vdd.n2286 gnd 0.010194f
C3612 vdd.n2287 gnd 0.008205f
C3613 vdd.n2288 gnd 0.010194f
C3614 vdd.n2289 gnd 0.651129f
C3615 vdd.n2290 gnd 0.010194f
C3616 vdd.n2291 gnd 0.008205f
C3617 vdd.n2292 gnd 0.010194f
C3618 vdd.n2293 gnd 0.010194f
C3619 vdd.n2294 gnd 0.010194f
C3620 vdd.n2295 gnd 0.008205f
C3621 vdd.n2296 gnd 0.010194f
C3622 vdd.n2297 gnd 0.557367f
C3623 vdd.n2298 gnd 0.828236f
C3624 vdd.n2299 gnd 0.010194f
C3625 vdd.n2300 gnd 0.008205f
C3626 vdd.n2301 gnd 0.010194f
C3627 vdd.n2302 gnd 0.010194f
C3628 vdd.n2303 gnd 0.010194f
C3629 vdd.n2304 gnd 0.008205f
C3630 vdd.n2305 gnd 0.010194f
C3631 vdd.n2306 gnd 0.864699f
C3632 vdd.n2307 gnd 0.010194f
C3633 vdd.n2308 gnd 0.008205f
C3634 vdd.n2309 gnd 0.010194f
C3635 vdd.n2310 gnd 0.010194f
C3636 vdd.n2311 gnd 0.010194f
C3637 vdd.n2312 gnd 0.008205f
C3638 vdd.n2313 gnd 0.010194f
C3639 vdd.t174 gnd 0.520903f
C3640 vdd.n2314 gnd 0.724056f
C3641 vdd.n2315 gnd 0.010194f
C3642 vdd.n2316 gnd 0.008205f
C3643 vdd.n2317 gnd 0.010194f
C3644 vdd.n2318 gnd 0.010194f
C3645 vdd.n2319 gnd 0.010194f
C3646 vdd.n2320 gnd 0.008205f
C3647 vdd.n2321 gnd 0.010194f
C3648 vdd.n2322 gnd 0.546948f
C3649 vdd.n2323 gnd 0.010194f
C3650 vdd.n2324 gnd 0.008205f
C3651 vdd.n2325 gnd 0.010194f
C3652 vdd.n2326 gnd 0.010194f
C3653 vdd.n2327 gnd 0.010194f
C3654 vdd.n2328 gnd 0.008205f
C3655 vdd.n2329 gnd 0.010194f
C3656 vdd.n2330 gnd 0.713638f
C3657 vdd.n2331 gnd 0.671965f
C3658 vdd.n2332 gnd 0.010194f
C3659 vdd.n2333 gnd 0.008205f
C3660 vdd.n2334 gnd 0.010194f
C3661 vdd.n2335 gnd 0.010194f
C3662 vdd.n2336 gnd 0.010194f
C3663 vdd.n2337 gnd 0.008205f
C3664 vdd.n2338 gnd 0.010194f
C3665 vdd.n2339 gnd 0.849072f
C3666 vdd.n2340 gnd 0.010194f
C3667 vdd.n2341 gnd 0.008205f
C3668 vdd.n2342 gnd 0.010194f
C3669 vdd.n2343 gnd 0.010194f
C3670 vdd.n2344 gnd 0.024661f
C3671 vdd.n2345 gnd 0.010194f
C3672 vdd.n2346 gnd 0.010194f
C3673 vdd.n2347 gnd 0.008205f
C3674 vdd.n2348 gnd 0.010194f
C3675 vdd.n2349 gnd 0.630293f
C3676 vdd.n2350 gnd 1.04181f
C3677 vdd.n2351 gnd 0.010194f
C3678 vdd.n2352 gnd 0.008205f
C3679 vdd.n2353 gnd 0.010194f
C3680 vdd.n2354 gnd 0.010194f
C3681 vdd.n2355 gnd 0.024661f
C3682 vdd.n2356 gnd 0.00681f
C3683 vdd.n2357 gnd 0.024661f
C3684 vdd.n2358 gnd 1.43248f
C3685 vdd.n2359 gnd 0.024661f
C3686 vdd.n2360 gnd 0.025189f
C3687 vdd.n2361 gnd 0.003897f
C3688 vdd.t118 gnd 0.125416f
C3689 vdd.t117 gnd 0.134036f
C3690 vdd.t116 gnd 0.163792f
C3691 vdd.n2362 gnd 0.209958f
C3692 vdd.n2363 gnd 0.176403f
C3693 vdd.n2364 gnd 0.012636f
C3694 vdd.n2365 gnd 0.004308f
C3695 vdd.n2366 gnd 0.008767f
C3696 vdd.n2367 gnd 1.08223f
C3697 vdd.n2369 gnd 0.008205f
C3698 vdd.n2370 gnd 0.008205f
C3699 vdd.n2371 gnd 0.010194f
C3700 vdd.n2373 gnd 0.010194f
C3701 vdd.n2374 gnd 0.010194f
C3702 vdd.n2375 gnd 0.008205f
C3703 vdd.n2376 gnd 0.008205f
C3704 vdd.n2377 gnd 0.008205f
C3705 vdd.n2378 gnd 0.010194f
C3706 vdd.n2380 gnd 0.010194f
C3707 vdd.n2381 gnd 0.010194f
C3708 vdd.n2382 gnd 0.008205f
C3709 vdd.n2383 gnd 0.008205f
C3710 vdd.n2384 gnd 0.008205f
C3711 vdd.n2385 gnd 0.010194f
C3712 vdd.n2387 gnd 0.010194f
C3713 vdd.n2388 gnd 0.010194f
C3714 vdd.n2389 gnd 0.008205f
C3715 vdd.n2390 gnd 0.008205f
C3716 vdd.n2391 gnd 0.008205f
C3717 vdd.n2392 gnd 0.010194f
C3718 vdd.n2394 gnd 0.010194f
C3719 vdd.n2395 gnd 0.010194f
C3720 vdd.n2396 gnd 0.008205f
C3721 vdd.n2397 gnd 0.010194f
C3722 vdd.n2398 gnd 0.010194f
C3723 vdd.n2399 gnd 0.010194f
C3724 vdd.n2400 gnd 0.016739f
C3725 vdd.n2401 gnd 0.00558f
C3726 vdd.n2402 gnd 0.008205f
C3727 vdd.n2403 gnd 0.010194f
C3728 vdd.n2405 gnd 0.010194f
C3729 vdd.n2406 gnd 0.010194f
C3730 vdd.n2407 gnd 0.008205f
C3731 vdd.n2408 gnd 0.008205f
C3732 vdd.n2409 gnd 0.008205f
C3733 vdd.n2410 gnd 0.010194f
C3734 vdd.n2412 gnd 0.010194f
C3735 vdd.n2413 gnd 0.010194f
C3736 vdd.n2414 gnd 0.008205f
C3737 vdd.n2415 gnd 0.008205f
C3738 vdd.n2416 gnd 0.008205f
C3739 vdd.n2417 gnd 0.010194f
C3740 vdd.n2419 gnd 0.010194f
C3741 vdd.n2420 gnd 0.010194f
C3742 vdd.n2421 gnd 0.008205f
C3743 vdd.n2422 gnd 0.008205f
C3744 vdd.n2423 gnd 0.008205f
C3745 vdd.n2424 gnd 0.010194f
C3746 vdd.n2426 gnd 0.010194f
C3747 vdd.n2427 gnd 0.010194f
C3748 vdd.n2428 gnd 0.008205f
C3749 vdd.n2429 gnd 0.008205f
C3750 vdd.n2430 gnd 0.008205f
C3751 vdd.n2431 gnd 0.010194f
C3752 vdd.n2433 gnd 0.010194f
C3753 vdd.n2434 gnd 0.010194f
C3754 vdd.n2435 gnd 0.008205f
C3755 vdd.n2436 gnd 0.010194f
C3756 vdd.n2437 gnd 0.010194f
C3757 vdd.n2438 gnd 0.010194f
C3758 vdd.n2439 gnd 0.016739f
C3759 vdd.n2440 gnd 0.006851f
C3760 vdd.n2441 gnd 0.008205f
C3761 vdd.n2442 gnd 0.010194f
C3762 vdd.n2444 gnd 0.010194f
C3763 vdd.n2445 gnd 0.010194f
C3764 vdd.n2446 gnd 0.008205f
C3765 vdd.n2447 gnd 0.008205f
C3766 vdd.n2448 gnd 0.008205f
C3767 vdd.n2449 gnd 0.010194f
C3768 vdd.n2451 gnd 0.010194f
C3769 vdd.n2452 gnd 0.010194f
C3770 vdd.n2453 gnd 0.008205f
C3771 vdd.n2454 gnd 0.008205f
C3772 vdd.n2455 gnd 0.008205f
C3773 vdd.n2456 gnd 0.010194f
C3774 vdd.n2458 gnd 0.010194f
C3775 vdd.n2459 gnd 0.010194f
C3776 vdd.n2460 gnd 0.008205f
C3777 vdd.n2461 gnd 0.008205f
C3778 vdd.n2462 gnd 0.008205f
C3779 vdd.n2463 gnd 0.010194f
C3780 vdd.n2465 gnd 0.010194f
C3781 vdd.n2466 gnd 0.008205f
C3782 vdd.n2467 gnd 0.008205f
C3783 vdd.n2468 gnd 0.010194f
C3784 vdd.n2470 gnd 0.010194f
C3785 vdd.n2471 gnd 0.010194f
C3786 vdd.n2472 gnd 0.008205f
C3787 vdd.n2473 gnd 0.008767f
C3788 vdd.n2474 gnd 1.08223f
C3789 vdd.n2475 gnd 0.046698f
C3790 vdd.n2476 gnd 0.006932f
C3791 vdd.n2477 gnd 0.006932f
C3792 vdd.n2478 gnd 0.006932f
C3793 vdd.n2479 gnd 0.006932f
C3794 vdd.n2480 gnd 0.006932f
C3795 vdd.n2481 gnd 0.006932f
C3796 vdd.n2482 gnd 0.006932f
C3797 vdd.n2483 gnd 0.006932f
C3798 vdd.n2484 gnd 0.006932f
C3799 vdd.n2485 gnd 0.006932f
C3800 vdd.n2486 gnd 0.006932f
C3801 vdd.n2487 gnd 0.006932f
C3802 vdd.n2488 gnd 0.006932f
C3803 vdd.n2489 gnd 0.006932f
C3804 vdd.n2490 gnd 0.006932f
C3805 vdd.n2491 gnd 0.006932f
C3806 vdd.n2492 gnd 0.006932f
C3807 vdd.n2493 gnd 0.006932f
C3808 vdd.n2494 gnd 0.006932f
C3809 vdd.n2495 gnd 0.006932f
C3810 vdd.n2496 gnd 0.006932f
C3811 vdd.n2497 gnd 0.006932f
C3812 vdd.n2498 gnd 0.006932f
C3813 vdd.n2499 gnd 0.006932f
C3814 vdd.n2500 gnd 0.006932f
C3815 vdd.n2501 gnd 0.006932f
C3816 vdd.n2502 gnd 0.006932f
C3817 vdd.n2503 gnd 0.006932f
C3818 vdd.n2504 gnd 0.006932f
C3819 vdd.n2505 gnd 0.006932f
C3820 vdd.n2506 gnd 12.303699f
C3821 vdd.n2508 gnd 0.01574f
C3822 vdd.n2509 gnd 0.01574f
C3823 vdd.n2510 gnd 0.014843f
C3824 vdd.n2511 gnd 0.006932f
C3825 vdd.n2512 gnd 0.006932f
C3826 vdd.n2513 gnd 0.708428f
C3827 vdd.n2514 gnd 0.006932f
C3828 vdd.n2515 gnd 0.006932f
C3829 vdd.n2516 gnd 0.006932f
C3830 vdd.n2517 gnd 0.006932f
C3831 vdd.n2518 gnd 0.006932f
C3832 vdd.n2519 gnd 0.557367f
C3833 vdd.n2520 gnd 0.006932f
C3834 vdd.n2521 gnd 0.006932f
C3835 vdd.n2522 gnd 0.006932f
C3836 vdd.n2523 gnd 0.006932f
C3837 vdd.n2524 gnd 0.006932f
C3838 vdd.n2525 gnd 0.708428f
C3839 vdd.n2526 gnd 0.006932f
C3840 vdd.n2527 gnd 0.006932f
C3841 vdd.n2528 gnd 0.006932f
C3842 vdd.n2529 gnd 0.006932f
C3843 vdd.n2530 gnd 0.006932f
C3844 vdd.n2531 gnd 0.708428f
C3845 vdd.n2532 gnd 0.006932f
C3846 vdd.n2533 gnd 0.006932f
C3847 vdd.n2534 gnd 0.006932f
C3848 vdd.n2535 gnd 0.006932f
C3849 vdd.n2536 gnd 0.006932f
C3850 vdd.n2537 gnd 0.682383f
C3851 vdd.n2538 gnd 0.006932f
C3852 vdd.n2539 gnd 0.006932f
C3853 vdd.n2540 gnd 0.006932f
C3854 vdd.n2541 gnd 0.006932f
C3855 vdd.n2542 gnd 0.006932f
C3856 vdd.n2543 gnd 0.526112f
C3857 vdd.n2544 gnd 0.006932f
C3858 vdd.n2545 gnd 0.006932f
C3859 vdd.n2546 gnd 0.006932f
C3860 vdd.n2547 gnd 0.006932f
C3861 vdd.n2548 gnd 0.006932f
C3862 vdd.n2549 gnd 0.369841f
C3863 vdd.n2550 gnd 0.006932f
C3864 vdd.n2551 gnd 0.006932f
C3865 vdd.n2552 gnd 0.006932f
C3866 vdd.n2553 gnd 0.006932f
C3867 vdd.n2554 gnd 0.006932f
C3868 vdd.n2555 gnd 0.494858f
C3869 vdd.n2556 gnd 0.006932f
C3870 vdd.n2557 gnd 0.006932f
C3871 vdd.n2558 gnd 0.006932f
C3872 vdd.n2559 gnd 0.006932f
C3873 vdd.n2560 gnd 0.006932f
C3874 vdd.n2561 gnd 0.651129f
C3875 vdd.n2562 gnd 0.006932f
C3876 vdd.n2563 gnd 0.006932f
C3877 vdd.n2564 gnd 0.006932f
C3878 vdd.n2565 gnd 0.006932f
C3879 vdd.n2566 gnd 0.006932f
C3880 vdd.n2567 gnd 0.708428f
C3881 vdd.n2568 gnd 0.006932f
C3882 vdd.n2569 gnd 0.006932f
C3883 vdd.n2570 gnd 0.006932f
C3884 vdd.n2571 gnd 0.006932f
C3885 vdd.n2572 gnd 0.006932f
C3886 vdd.n2573 gnd 0.609457f
C3887 vdd.n2574 gnd 0.006932f
C3888 vdd.n2575 gnd 0.006932f
C3889 vdd.n2576 gnd 0.005505f
C3890 vdd.n2577 gnd 0.020081f
C3891 vdd.n2578 gnd 0.004893f
C3892 vdd.n2579 gnd 0.006932f
C3893 vdd.n2580 gnd 0.453186f
C3894 vdd.n2581 gnd 0.006932f
C3895 vdd.n2582 gnd 0.006932f
C3896 vdd.n2583 gnd 0.006932f
C3897 vdd.n2584 gnd 0.006932f
C3898 vdd.n2585 gnd 0.006932f
C3899 vdd.n2586 gnd 0.411514f
C3900 vdd.n2587 gnd 0.006932f
C3901 vdd.n2588 gnd 0.006932f
C3902 vdd.n2589 gnd 0.006932f
C3903 vdd.n2590 gnd 0.006932f
C3904 vdd.n2591 gnd 0.006932f
C3905 vdd.n2592 gnd 0.567785f
C3906 vdd.n2593 gnd 0.006932f
C3907 vdd.n2594 gnd 0.006932f
C3908 vdd.n2595 gnd 0.006932f
C3909 vdd.n2596 gnd 0.006932f
C3910 vdd.n2597 gnd 0.006932f
C3911 vdd.n2598 gnd 0.625084f
C3912 vdd.n2599 gnd 0.006932f
C3913 vdd.n2600 gnd 0.006932f
C3914 vdd.n2601 gnd 0.006932f
C3915 vdd.n2602 gnd 0.006932f
C3916 vdd.n2603 gnd 0.006932f
C3917 vdd.n2604 gnd 0.468813f
C3918 vdd.n2605 gnd 0.006932f
C3919 vdd.n2606 gnd 0.006932f
C3920 vdd.n2607 gnd 0.006932f
C3921 vdd.n2608 gnd 0.006932f
C3922 vdd.n2609 gnd 0.006932f
C3923 vdd.n2610 gnd 0.223988f
C3924 vdd.n2611 gnd 0.006932f
C3925 vdd.n2612 gnd 0.006932f
C3926 vdd.n2613 gnd 0.006932f
C3927 vdd.n2614 gnd 0.006932f
C3928 vdd.n2615 gnd 0.006932f
C3929 vdd.n2616 gnd 0.223988f
C3930 vdd.n2617 gnd 0.006932f
C3931 vdd.n2618 gnd 0.006932f
C3932 vdd.n2619 gnd 0.006932f
C3933 vdd.n2620 gnd 0.006932f
C3934 vdd.n2621 gnd 0.006932f
C3935 vdd.n2622 gnd 0.708428f
C3936 vdd.n2623 gnd 0.006932f
C3937 vdd.n2624 gnd 0.006932f
C3938 vdd.n2625 gnd 0.006932f
C3939 vdd.n2626 gnd 0.006932f
C3940 vdd.n2627 gnd 0.006932f
C3941 vdd.n2628 gnd 0.006932f
C3942 vdd.n2629 gnd 0.006932f
C3943 vdd.n2630 gnd 0.489649f
C3944 vdd.n2631 gnd 0.006932f
C3945 vdd.n2632 gnd 0.006932f
C3946 vdd.n2633 gnd 0.006932f
C3947 vdd.n2634 gnd 0.006932f
C3948 vdd.n2635 gnd 0.006932f
C3949 vdd.n2636 gnd 0.006932f
C3950 vdd.n2637 gnd 0.442768f
C3951 vdd.n2638 gnd 0.006932f
C3952 vdd.n2639 gnd 0.006932f
C3953 vdd.n2640 gnd 0.006932f
C3954 vdd.n2641 gnd 0.01574f
C3955 vdd.n2642 gnd 0.014843f
C3956 vdd.n2643 gnd 0.006932f
C3957 vdd.n2644 gnd 0.006932f
C3958 vdd.n2645 gnd 0.005352f
C3959 vdd.n2646 gnd 0.006932f
C3960 vdd.n2647 gnd 0.006932f
C3961 vdd.n2648 gnd 0.005046f
C3962 vdd.n2649 gnd 0.006932f
C3963 vdd.n2650 gnd 0.006932f
C3964 vdd.n2651 gnd 0.006932f
C3965 vdd.n2652 gnd 0.006932f
C3966 vdd.n2653 gnd 0.006932f
C3967 vdd.n2654 gnd 0.006932f
C3968 vdd.n2655 gnd 0.006932f
C3969 vdd.n2656 gnd 0.006932f
C3970 vdd.n2657 gnd 0.006932f
C3971 vdd.n2658 gnd 0.006932f
C3972 vdd.n2659 gnd 0.006932f
C3973 vdd.n2660 gnd 0.006932f
C3974 vdd.n2661 gnd 0.006932f
C3975 vdd.n2662 gnd 0.006932f
C3976 vdd.n2663 gnd 0.006932f
C3977 vdd.n2664 gnd 0.006932f
C3978 vdd.n2665 gnd 0.006932f
C3979 vdd.n2666 gnd 0.006932f
C3980 vdd.n2667 gnd 0.006932f
C3981 vdd.n2668 gnd 0.006932f
C3982 vdd.n2669 gnd 0.006932f
C3983 vdd.n2670 gnd 0.006932f
C3984 vdd.n2671 gnd 0.006932f
C3985 vdd.n2672 gnd 0.006932f
C3986 vdd.n2673 gnd 0.006932f
C3987 vdd.n2674 gnd 0.006932f
C3988 vdd.n2675 gnd 0.006932f
C3989 vdd.n2676 gnd 0.006932f
C3990 vdd.n2677 gnd 0.006932f
C3991 vdd.n2678 gnd 0.006932f
C3992 vdd.n2679 gnd 0.006932f
C3993 vdd.n2680 gnd 0.006932f
C3994 vdd.n2681 gnd 0.006932f
C3995 vdd.n2682 gnd 0.006932f
C3996 vdd.n2683 gnd 0.006932f
C3997 vdd.n2684 gnd 0.006932f
C3998 vdd.n2685 gnd 0.006932f
C3999 vdd.n2686 gnd 0.006932f
C4000 vdd.n2687 gnd 0.006932f
C4001 vdd.n2688 gnd 0.006932f
C4002 vdd.n2689 gnd 0.006932f
C4003 vdd.n2690 gnd 0.006932f
C4004 vdd.n2691 gnd 0.006932f
C4005 vdd.n2692 gnd 0.006932f
C4006 vdd.n2693 gnd 0.006932f
C4007 vdd.n2694 gnd 0.006932f
C4008 vdd.n2695 gnd 0.006932f
C4009 vdd.n2696 gnd 0.006932f
C4010 vdd.n2697 gnd 0.006932f
C4011 vdd.n2698 gnd 0.006932f
C4012 vdd.n2699 gnd 0.006932f
C4013 vdd.n2700 gnd 0.006932f
C4014 vdd.n2701 gnd 0.006932f
C4015 vdd.n2702 gnd 0.006932f
C4016 vdd.n2703 gnd 0.006932f
C4017 vdd.n2704 gnd 0.006932f
C4018 vdd.n2705 gnd 0.006932f
C4019 vdd.n2706 gnd 0.006932f
C4020 vdd.n2707 gnd 0.006932f
C4021 vdd.n2708 gnd 0.006932f
C4022 vdd.n2709 gnd 0.01574f
C4023 vdd.n2710 gnd 0.014843f
C4024 vdd.n2711 gnd 0.014843f
C4025 vdd.n2712 gnd 0.802191f
C4026 vdd.n2713 gnd 0.014843f
C4027 vdd.n2714 gnd 0.01574f
C4028 vdd.n2715 gnd 0.014843f
C4029 vdd.n2716 gnd 0.006932f
C4030 vdd.n2717 gnd 0.006932f
C4031 vdd.n2718 gnd 0.006932f
C4032 vdd.n2719 gnd 0.005352f
C4033 vdd.n2720 gnd 0.009907f
C4034 vdd.n2721 gnd 0.005046f
C4035 vdd.n2722 gnd 0.006932f
C4036 vdd.n2723 gnd 0.006932f
C4037 vdd.n2724 gnd 0.006932f
C4038 vdd.n2725 gnd 0.006932f
C4039 vdd.n2726 gnd 0.006932f
C4040 vdd.n2727 gnd 0.006932f
C4041 vdd.n2728 gnd 0.006932f
C4042 vdd.n2729 gnd 0.006932f
C4043 vdd.n2730 gnd 0.006932f
C4044 vdd.n2731 gnd 0.006932f
C4045 vdd.n2732 gnd 0.006932f
C4046 vdd.n2733 gnd 0.006932f
C4047 vdd.n2734 gnd 0.006932f
C4048 vdd.n2735 gnd 0.006932f
C4049 vdd.n2736 gnd 0.006932f
C4050 vdd.n2737 gnd 0.006932f
C4051 vdd.n2738 gnd 0.006932f
C4052 vdd.n2739 gnd 0.006932f
C4053 vdd.n2740 gnd 0.006932f
C4054 vdd.n2741 gnd 0.006932f
C4055 vdd.n2742 gnd 0.006932f
C4056 vdd.n2743 gnd 0.006932f
C4057 vdd.n2744 gnd 0.006932f
C4058 vdd.n2745 gnd 0.006932f
C4059 vdd.n2746 gnd 0.006932f
C4060 vdd.n2747 gnd 0.006932f
C4061 vdd.n2748 gnd 0.006932f
C4062 vdd.n2749 gnd 0.006932f
C4063 vdd.n2750 gnd 0.006932f
C4064 vdd.n2751 gnd 0.006932f
C4065 vdd.n2752 gnd 0.006932f
C4066 vdd.n2753 gnd 0.006932f
C4067 vdd.n2754 gnd 0.006932f
C4068 vdd.n2755 gnd 0.006932f
C4069 vdd.n2756 gnd 0.006932f
C4070 vdd.n2757 gnd 0.006932f
C4071 vdd.n2758 gnd 0.006932f
C4072 vdd.n2759 gnd 0.006932f
C4073 vdd.n2760 gnd 0.006932f
C4074 vdd.n2761 gnd 0.006932f
C4075 vdd.n2762 gnd 0.006932f
C4076 vdd.n2763 gnd 0.006932f
C4077 vdd.n2764 gnd 0.006932f
C4078 vdd.n2765 gnd 0.006932f
C4079 vdd.n2766 gnd 0.006932f
C4080 vdd.n2767 gnd 0.006932f
C4081 vdd.n2768 gnd 0.006932f
C4082 vdd.n2769 gnd 0.006932f
C4083 vdd.n2770 gnd 0.006932f
C4084 vdd.n2771 gnd 0.006932f
C4085 vdd.n2772 gnd 0.006932f
C4086 vdd.n2773 gnd 0.006932f
C4087 vdd.n2774 gnd 0.006932f
C4088 vdd.n2775 gnd 0.006932f
C4089 vdd.n2776 gnd 0.006932f
C4090 vdd.n2777 gnd 0.006932f
C4091 vdd.n2778 gnd 0.006932f
C4092 vdd.n2779 gnd 0.006932f
C4093 vdd.n2780 gnd 0.006932f
C4094 vdd.n2781 gnd 0.006932f
C4095 vdd.n2782 gnd 0.01574f
C4096 vdd.n2783 gnd 0.01574f
C4097 vdd.n2784 gnd 0.864699f
C4098 vdd.t264 gnd 3.07333f
C4099 vdd.t240 gnd 3.07333f
C4100 vdd.n2818 gnd 0.01574f
C4101 vdd.t269 gnd 0.604248f
C4102 vdd.n2819 gnd 0.006932f
C4103 vdd.t137 gnd 0.280125f
C4104 vdd.t138 gnd 0.286743f
C4105 vdd.t135 gnd 0.182877f
C4106 vdd.n2820 gnd 0.098835f
C4107 vdd.n2821 gnd 0.056062f
C4108 vdd.n2822 gnd 0.006932f
C4109 vdd.t144 gnd 0.280125f
C4110 vdd.t145 gnd 0.286743f
C4111 vdd.t143 gnd 0.182877f
C4112 vdd.n2823 gnd 0.098835f
C4113 vdd.n2824 gnd 0.056062f
C4114 vdd.n2825 gnd 0.009907f
C4115 vdd.n2826 gnd 0.01574f
C4116 vdd.n2827 gnd 0.01574f
C4117 vdd.n2828 gnd 0.006932f
C4118 vdd.n2829 gnd 0.006932f
C4119 vdd.n2830 gnd 0.006932f
C4120 vdd.n2831 gnd 0.006932f
C4121 vdd.n2832 gnd 0.006932f
C4122 vdd.n2833 gnd 0.006932f
C4123 vdd.n2834 gnd 0.006932f
C4124 vdd.n2835 gnd 0.006932f
C4125 vdd.n2836 gnd 0.006932f
C4126 vdd.n2837 gnd 0.006932f
C4127 vdd.n2838 gnd 0.006932f
C4128 vdd.n2839 gnd 0.006932f
C4129 vdd.n2840 gnd 0.006932f
C4130 vdd.n2841 gnd 0.006932f
C4131 vdd.n2842 gnd 0.006932f
C4132 vdd.n2843 gnd 0.006932f
C4133 vdd.n2844 gnd 0.006932f
C4134 vdd.n2845 gnd 0.006932f
C4135 vdd.n2846 gnd 0.006932f
C4136 vdd.n2847 gnd 0.006932f
C4137 vdd.n2848 gnd 0.006932f
C4138 vdd.n2849 gnd 0.006932f
C4139 vdd.n2850 gnd 0.006932f
C4140 vdd.n2851 gnd 0.006932f
C4141 vdd.n2852 gnd 0.006932f
C4142 vdd.n2853 gnd 0.006932f
C4143 vdd.n2854 gnd 0.006932f
C4144 vdd.n2855 gnd 0.006932f
C4145 vdd.n2856 gnd 0.006932f
C4146 vdd.n2857 gnd 0.006932f
C4147 vdd.n2858 gnd 0.006932f
C4148 vdd.n2859 gnd 0.006932f
C4149 vdd.n2860 gnd 0.006932f
C4150 vdd.n2861 gnd 0.006932f
C4151 vdd.n2862 gnd 0.006932f
C4152 vdd.n2863 gnd 0.006932f
C4153 vdd.n2864 gnd 0.006932f
C4154 vdd.n2865 gnd 0.006932f
C4155 vdd.n2866 gnd 0.006932f
C4156 vdd.n2867 gnd 0.006932f
C4157 vdd.n2868 gnd 0.006932f
C4158 vdd.n2869 gnd 0.006932f
C4159 vdd.n2870 gnd 0.006932f
C4160 vdd.n2871 gnd 0.006932f
C4161 vdd.n2872 gnd 0.006932f
C4162 vdd.n2873 gnd 0.006932f
C4163 vdd.n2874 gnd 0.006932f
C4164 vdd.n2875 gnd 0.006932f
C4165 vdd.n2876 gnd 0.006932f
C4166 vdd.n2877 gnd 0.006932f
C4167 vdd.n2878 gnd 0.006932f
C4168 vdd.n2879 gnd 0.006932f
C4169 vdd.n2880 gnd 0.006932f
C4170 vdd.n2881 gnd 0.006932f
C4171 vdd.n2882 gnd 0.006932f
C4172 vdd.n2883 gnd 0.006932f
C4173 vdd.n2884 gnd 0.006932f
C4174 vdd.n2885 gnd 0.006932f
C4175 vdd.n2886 gnd 0.006932f
C4176 vdd.n2887 gnd 0.006932f
C4177 vdd.n2888 gnd 0.005046f
C4178 vdd.n2889 gnd 0.006932f
C4179 vdd.n2890 gnd 0.006932f
C4180 vdd.n2891 gnd 0.005352f
C4181 vdd.n2892 gnd 0.006932f
C4182 vdd.n2893 gnd 0.006932f
C4183 vdd.n2894 gnd 0.01574f
C4184 vdd.n2895 gnd 0.014843f
C4185 vdd.n2896 gnd 0.014843f
C4186 vdd.n2897 gnd 0.006932f
C4187 vdd.n2898 gnd 0.006932f
C4188 vdd.n2899 gnd 0.006932f
C4189 vdd.n2900 gnd 0.006932f
C4190 vdd.n2901 gnd 0.006932f
C4191 vdd.n2902 gnd 0.006932f
C4192 vdd.n2903 gnd 0.006932f
C4193 vdd.n2904 gnd 0.006932f
C4194 vdd.n2905 gnd 0.006932f
C4195 vdd.n2906 gnd 0.006932f
C4196 vdd.n2907 gnd 0.006932f
C4197 vdd.n2908 gnd 0.006932f
C4198 vdd.n2909 gnd 0.006932f
C4199 vdd.n2910 gnd 0.006932f
C4200 vdd.n2911 gnd 0.006932f
C4201 vdd.n2912 gnd 0.006932f
C4202 vdd.n2913 gnd 0.006932f
C4203 vdd.n2914 gnd 0.006932f
C4204 vdd.n2915 gnd 0.006932f
C4205 vdd.n2916 gnd 0.006932f
C4206 vdd.n2917 gnd 0.006932f
C4207 vdd.n2918 gnd 0.006932f
C4208 vdd.n2919 gnd 0.006932f
C4209 vdd.n2920 gnd 0.006932f
C4210 vdd.n2921 gnd 0.006932f
C4211 vdd.n2922 gnd 0.006932f
C4212 vdd.n2923 gnd 0.006932f
C4213 vdd.n2924 gnd 0.006932f
C4214 vdd.n2925 gnd 0.006932f
C4215 vdd.n2926 gnd 0.006932f
C4216 vdd.n2927 gnd 0.006932f
C4217 vdd.n2928 gnd 0.006932f
C4218 vdd.n2929 gnd 0.006932f
C4219 vdd.n2930 gnd 0.006932f
C4220 vdd.n2931 gnd 0.006932f
C4221 vdd.n2932 gnd 0.006932f
C4222 vdd.n2933 gnd 0.006932f
C4223 vdd.n2934 gnd 0.006932f
C4224 vdd.n2935 gnd 0.006932f
C4225 vdd.n2936 gnd 0.006932f
C4226 vdd.n2937 gnd 0.006932f
C4227 vdd.n2938 gnd 0.006932f
C4228 vdd.n2939 gnd 0.006932f
C4229 vdd.n2940 gnd 0.006932f
C4230 vdd.n2941 gnd 0.006932f
C4231 vdd.n2942 gnd 0.006932f
C4232 vdd.n2943 gnd 0.006932f
C4233 vdd.n2944 gnd 0.006932f
C4234 vdd.n2945 gnd 0.006932f
C4235 vdd.n2946 gnd 0.006932f
C4236 vdd.n2947 gnd 0.006932f
C4237 vdd.n2948 gnd 0.006932f
C4238 vdd.n2949 gnd 0.006932f
C4239 vdd.n2950 gnd 0.006932f
C4240 vdd.n2951 gnd 0.006932f
C4241 vdd.n2952 gnd 0.006932f
C4242 vdd.n2953 gnd 0.006932f
C4243 vdd.n2954 gnd 0.006932f
C4244 vdd.n2955 gnd 0.006932f
C4245 vdd.n2956 gnd 0.006932f
C4246 vdd.n2957 gnd 0.006932f
C4247 vdd.n2958 gnd 0.006932f
C4248 vdd.n2959 gnd 0.006932f
C4249 vdd.n2960 gnd 0.006932f
C4250 vdd.n2961 gnd 0.006932f
C4251 vdd.n2962 gnd 0.006932f
C4252 vdd.n2963 gnd 0.006932f
C4253 vdd.n2964 gnd 0.006932f
C4254 vdd.n2965 gnd 0.006932f
C4255 vdd.n2966 gnd 0.006932f
C4256 vdd.n2967 gnd 0.006932f
C4257 vdd.n2968 gnd 0.006932f
C4258 vdd.n2969 gnd 0.006932f
C4259 vdd.n2970 gnd 0.006932f
C4260 vdd.n2971 gnd 0.006932f
C4261 vdd.n2972 gnd 0.006932f
C4262 vdd.n2973 gnd 0.006932f
C4263 vdd.n2974 gnd 0.006932f
C4264 vdd.n2975 gnd 0.006932f
C4265 vdd.n2976 gnd 0.006932f
C4266 vdd.n2977 gnd 0.006932f
C4267 vdd.n2978 gnd 0.006932f
C4268 vdd.n2979 gnd 0.006932f
C4269 vdd.n2980 gnd 0.006932f
C4270 vdd.n2981 gnd 0.006932f
C4271 vdd.n2982 gnd 0.006932f
C4272 vdd.n2983 gnd 0.006932f
C4273 vdd.n2984 gnd 0.006932f
C4274 vdd.n2985 gnd 0.006932f
C4275 vdd.n2986 gnd 0.006932f
C4276 vdd.n2987 gnd 0.006932f
C4277 vdd.n2988 gnd 0.006932f
C4278 vdd.n2989 gnd 0.006932f
C4279 vdd.n2990 gnd 0.006932f
C4280 vdd.n2991 gnd 0.006932f
C4281 vdd.n2992 gnd 0.006932f
C4282 vdd.n2993 gnd 0.006932f
C4283 vdd.n2994 gnd 0.006932f
C4284 vdd.n2995 gnd 0.006932f
C4285 vdd.n2996 gnd 0.006932f
C4286 vdd.n2997 gnd 0.006932f
C4287 vdd.n2998 gnd 0.223988f
C4288 vdd.n2999 gnd 0.006932f
C4289 vdd.n3000 gnd 0.006932f
C4290 vdd.n3001 gnd 0.006932f
C4291 vdd.n3002 gnd 0.006932f
C4292 vdd.n3003 gnd 0.006932f
C4293 vdd.n3004 gnd 0.223988f
C4294 vdd.n3005 gnd 0.006932f
C4295 vdd.n3006 gnd 0.006932f
C4296 vdd.n3007 gnd 0.006932f
C4297 vdd.n3008 gnd 0.006932f
C4298 vdd.n3009 gnd 0.006932f
C4299 vdd.n3010 gnd 0.006932f
C4300 vdd.n3011 gnd 0.006932f
C4301 vdd.n3012 gnd 0.006932f
C4302 vdd.n3013 gnd 0.006932f
C4303 vdd.n3014 gnd 0.006932f
C4304 vdd.n3015 gnd 0.006932f
C4305 vdd.n3016 gnd 0.442768f
C4306 vdd.n3017 gnd 0.006932f
C4307 vdd.n3018 gnd 0.006932f
C4308 vdd.n3019 gnd 0.006932f
C4309 vdd.n3020 gnd 0.014843f
C4310 vdd.n3021 gnd 0.014843f
C4311 vdd.n3022 gnd 0.01574f
C4312 vdd.n3023 gnd 0.01574f
C4313 vdd.n3024 gnd 0.006932f
C4314 vdd.n3025 gnd 0.006932f
C4315 vdd.n3026 gnd 0.006932f
C4316 vdd.n3027 gnd 0.005352f
C4317 vdd.n3028 gnd 0.009907f
C4318 vdd.n3029 gnd 0.005046f
C4319 vdd.n3030 gnd 0.006932f
C4320 vdd.n3031 gnd 0.006932f
C4321 vdd.n3032 gnd 0.006932f
C4322 vdd.n3033 gnd 0.006932f
C4323 vdd.n3034 gnd 0.006932f
C4324 vdd.n3035 gnd 0.006932f
C4325 vdd.n3036 gnd 0.006932f
C4326 vdd.n3037 gnd 0.006932f
C4327 vdd.n3038 gnd 0.006932f
C4328 vdd.n3039 gnd 0.006932f
C4329 vdd.n3040 gnd 0.006932f
C4330 vdd.n3041 gnd 0.006932f
C4331 vdd.n3042 gnd 0.006932f
C4332 vdd.n3043 gnd 0.006932f
C4333 vdd.n3044 gnd 0.006932f
C4334 vdd.n3045 gnd 0.006932f
C4335 vdd.n3046 gnd 0.006932f
C4336 vdd.n3047 gnd 0.006932f
C4337 vdd.n3048 gnd 0.006932f
C4338 vdd.n3049 gnd 0.006932f
C4339 vdd.n3050 gnd 0.006932f
C4340 vdd.n3051 gnd 0.006932f
C4341 vdd.n3052 gnd 0.006932f
C4342 vdd.n3053 gnd 0.006932f
C4343 vdd.n3054 gnd 0.006932f
C4344 vdd.n3055 gnd 0.006932f
C4345 vdd.n3056 gnd 0.006932f
C4346 vdd.n3057 gnd 0.006932f
C4347 vdd.n3058 gnd 0.006932f
C4348 vdd.n3059 gnd 0.006932f
C4349 vdd.n3060 gnd 0.006932f
C4350 vdd.n3061 gnd 0.006932f
C4351 vdd.n3062 gnd 0.006932f
C4352 vdd.n3063 gnd 0.006932f
C4353 vdd.n3064 gnd 0.006932f
C4354 vdd.n3065 gnd 0.006932f
C4355 vdd.n3066 gnd 0.006932f
C4356 vdd.n3067 gnd 0.006932f
C4357 vdd.n3068 gnd 0.006932f
C4358 vdd.n3069 gnd 0.006932f
C4359 vdd.n3070 gnd 0.006932f
C4360 vdd.n3071 gnd 0.006932f
C4361 vdd.n3072 gnd 0.006932f
C4362 vdd.n3073 gnd 0.006932f
C4363 vdd.n3074 gnd 0.006932f
C4364 vdd.n3075 gnd 0.006932f
C4365 vdd.n3076 gnd 0.006932f
C4366 vdd.n3077 gnd 0.006932f
C4367 vdd.n3078 gnd 0.006932f
C4368 vdd.n3079 gnd 0.006932f
C4369 vdd.n3080 gnd 0.006932f
C4370 vdd.n3081 gnd 0.006932f
C4371 vdd.n3082 gnd 0.006932f
C4372 vdd.n3083 gnd 0.006932f
C4373 vdd.n3084 gnd 0.006932f
C4374 vdd.n3085 gnd 0.006932f
C4375 vdd.n3086 gnd 0.006932f
C4376 vdd.n3087 gnd 0.006932f
C4377 vdd.n3088 gnd 0.864699f
C4378 vdd.n3090 gnd 0.01574f
C4379 vdd.n3091 gnd 0.01574f
C4380 vdd.n3092 gnd 0.014843f
C4381 vdd.n3093 gnd 0.006932f
C4382 vdd.n3094 gnd 0.006932f
C4383 vdd.n3095 gnd 0.416723f
C4384 vdd.n3096 gnd 0.006932f
C4385 vdd.n3097 gnd 0.006932f
C4386 vdd.n3098 gnd 0.006932f
C4387 vdd.n3099 gnd 0.006932f
C4388 vdd.n3100 gnd 0.006932f
C4389 vdd.n3101 gnd 0.421932f
C4390 vdd.n3102 gnd 0.006932f
C4391 vdd.n3103 gnd 0.006932f
C4392 vdd.n3104 gnd 0.006932f
C4393 vdd.n3105 gnd 0.006932f
C4394 vdd.n3106 gnd 0.006932f
C4395 vdd.n3107 gnd 0.708428f
C4396 vdd.n3108 gnd 0.006932f
C4397 vdd.n3109 gnd 0.006932f
C4398 vdd.n3110 gnd 0.006932f
C4399 vdd.n3111 gnd 0.006932f
C4400 vdd.n3112 gnd 0.006932f
C4401 vdd.n3113 gnd 0.510485f
C4402 vdd.n3114 gnd 0.006932f
C4403 vdd.n3115 gnd 0.006932f
C4404 vdd.n3116 gnd 0.006932f
C4405 vdd.n3117 gnd 0.006932f
C4406 vdd.n3118 gnd 0.006932f
C4407 vdd.n3119 gnd 0.640711f
C4408 vdd.n3120 gnd 0.006932f
C4409 vdd.n3121 gnd 0.006932f
C4410 vdd.n3122 gnd 0.006932f
C4411 vdd.n3123 gnd 0.006932f
C4412 vdd.n3124 gnd 0.006932f
C4413 vdd.n3125 gnd 0.526112f
C4414 vdd.n3126 gnd 0.006932f
C4415 vdd.n3127 gnd 0.006932f
C4416 vdd.n3128 gnd 0.006932f
C4417 vdd.n3129 gnd 0.006932f
C4418 vdd.n3130 gnd 0.006932f
C4419 vdd.n3131 gnd 0.369841f
C4420 vdd.n3132 gnd 0.006932f
C4421 vdd.n3133 gnd 0.006932f
C4422 vdd.n3134 gnd 0.006932f
C4423 vdd.n3135 gnd 0.006932f
C4424 vdd.n3136 gnd 0.006932f
C4425 vdd.n3137 gnd 0.223988f
C4426 vdd.n3138 gnd 0.006932f
C4427 vdd.n3139 gnd 0.006932f
C4428 vdd.n3140 gnd 0.006932f
C4429 vdd.n3141 gnd 0.006932f
C4430 vdd.n3142 gnd 0.006932f
C4431 vdd.n3143 gnd 0.651129f
C4432 vdd.n3144 gnd 0.006932f
C4433 vdd.n3145 gnd 0.006932f
C4434 vdd.n3146 gnd 0.006932f
C4435 vdd.n3147 gnd 0.004893f
C4436 vdd.n3148 gnd 0.006932f
C4437 vdd.n3149 gnd 0.006932f
C4438 vdd.n3150 gnd 0.708428f
C4439 vdd.n3151 gnd 0.006932f
C4440 vdd.n3152 gnd 0.006932f
C4441 vdd.n3153 gnd 0.006932f
C4442 vdd.n3154 gnd 0.006932f
C4443 vdd.n3155 gnd 0.006932f
C4444 vdd.n3156 gnd 0.562576f
C4445 vdd.n3157 gnd 0.006932f
C4446 vdd.n3158 gnd 0.005505f
C4447 vdd.n3159 gnd 0.006932f
C4448 vdd.n3160 gnd 0.006932f
C4449 vdd.n3161 gnd 0.006932f
C4450 vdd.n3162 gnd 0.453186f
C4451 vdd.n3163 gnd 0.006932f
C4452 vdd.n3164 gnd 0.006932f
C4453 vdd.n3165 gnd 0.006932f
C4454 vdd.n3166 gnd 0.006932f
C4455 vdd.n3167 gnd 0.006932f
C4456 vdd.n3168 gnd 0.411514f
C4457 vdd.n3169 gnd 0.006932f
C4458 vdd.n3170 gnd 0.006932f
C4459 vdd.n3171 gnd 0.006932f
C4460 vdd.n3172 gnd 0.006932f
C4461 vdd.n3173 gnd 0.006932f
C4462 vdd.n3174 gnd 0.567785f
C4463 vdd.n3175 gnd 0.006932f
C4464 vdd.n3176 gnd 0.006932f
C4465 vdd.n3177 gnd 0.006932f
C4466 vdd.n3178 gnd 0.006932f
C4467 vdd.n3179 gnd 0.006932f
C4468 vdd.n3180 gnd 0.708428f
C4469 vdd.n3181 gnd 0.006932f
C4470 vdd.n3182 gnd 0.006932f
C4471 vdd.n3183 gnd 0.006932f
C4472 vdd.n3184 gnd 0.006932f
C4473 vdd.n3185 gnd 0.006932f
C4474 vdd.n3186 gnd 0.692801f
C4475 vdd.n3187 gnd 0.006932f
C4476 vdd.n3188 gnd 0.006932f
C4477 vdd.n3189 gnd 0.006932f
C4478 vdd.n3190 gnd 0.006932f
C4479 vdd.n3191 gnd 0.006932f
C4480 vdd.n3192 gnd 0.53653f
C4481 vdd.n3193 gnd 0.006932f
C4482 vdd.n3194 gnd 0.006932f
C4483 vdd.n3195 gnd 0.006932f
C4484 vdd.n3196 gnd 0.006932f
C4485 vdd.n3197 gnd 0.006932f
C4486 vdd.n3198 gnd 0.380259f
C4487 vdd.n3199 gnd 0.006932f
C4488 vdd.n3200 gnd 0.006932f
C4489 vdd.n3201 gnd 0.006932f
C4490 vdd.n3202 gnd 0.006932f
C4491 vdd.n3203 gnd 0.006932f
C4492 vdd.n3204 gnd 0.708428f
C4493 vdd.n3205 gnd 0.006932f
C4494 vdd.n3206 gnd 0.006932f
C4495 vdd.n3207 gnd 0.006932f
C4496 vdd.n3208 gnd 0.006932f
C4497 vdd.n3209 gnd 0.006932f
C4498 vdd.n3210 gnd 0.006932f
C4499 vdd.n3212 gnd 0.006932f
C4500 vdd.n3213 gnd 0.006932f
C4501 vdd.n3215 gnd 0.006932f
C4502 vdd.n3216 gnd 0.006932f
C4503 vdd.n3219 gnd 0.006932f
C4504 vdd.n3220 gnd 0.006932f
C4505 vdd.n3221 gnd 0.006932f
C4506 vdd.n3222 gnd 0.006932f
C4507 vdd.n3224 gnd 0.006932f
C4508 vdd.n3225 gnd 0.006932f
C4509 vdd.n3226 gnd 0.006932f
C4510 vdd.n3227 gnd 0.006932f
C4511 vdd.n3228 gnd 0.006932f
C4512 vdd.n3229 gnd 0.006932f
C4513 vdd.n3231 gnd 0.006932f
C4514 vdd.n3232 gnd 0.006932f
C4515 vdd.n3233 gnd 0.006932f
C4516 vdd.n3234 gnd 0.006932f
C4517 vdd.n3235 gnd 0.006932f
C4518 vdd.n3236 gnd 0.006932f
C4519 vdd.n3238 gnd 0.006932f
C4520 vdd.n3239 gnd 0.006932f
C4521 vdd.n3240 gnd 0.006932f
C4522 vdd.n3241 gnd 0.006932f
C4523 vdd.n3242 gnd 0.006932f
C4524 vdd.n3243 gnd 0.006932f
C4525 vdd.n3245 gnd 0.006932f
C4526 vdd.n3246 gnd 0.01574f
C4527 vdd.n3247 gnd 0.01574f
C4528 vdd.n3248 gnd 0.014843f
C4529 vdd.n3249 gnd 0.006932f
C4530 vdd.n3250 gnd 0.006932f
C4531 vdd.n3251 gnd 0.006932f
C4532 vdd.n3252 gnd 0.006932f
C4533 vdd.n3253 gnd 0.006932f
C4534 vdd.n3254 gnd 0.006932f
C4535 vdd.n3255 gnd 0.708428f
C4536 vdd.n3256 gnd 0.006932f
C4537 vdd.n3257 gnd 0.006932f
C4538 vdd.n3258 gnd 0.006932f
C4539 vdd.n3259 gnd 0.006932f
C4540 vdd.n3260 gnd 0.006932f
C4541 vdd.n3261 gnd 0.505276f
C4542 vdd.n3262 gnd 0.006932f
C4543 vdd.n3263 gnd 0.006932f
C4544 vdd.n3264 gnd 0.006932f
C4545 vdd.n3265 gnd 0.01574f
C4546 vdd.n3266 gnd 0.014843f
C4547 vdd.n3267 gnd 0.01574f
C4548 vdd.n3269 gnd 0.006932f
C4549 vdd.n3270 gnd 0.006932f
C4550 vdd.n3271 gnd 0.005352f
C4551 vdd.n3272 gnd 0.009907f
C4552 vdd.n3273 gnd 0.005046f
C4553 vdd.n3274 gnd 0.006932f
C4554 vdd.n3275 gnd 0.006932f
C4555 vdd.n3277 gnd 0.006932f
C4556 vdd.n3278 gnd 0.006932f
C4557 vdd.n3279 gnd 0.006932f
C4558 vdd.n3280 gnd 0.006932f
C4559 vdd.n3281 gnd 0.006932f
C4560 vdd.n3282 gnd 0.006932f
C4561 vdd.n3284 gnd 0.006932f
C4562 vdd.n3285 gnd 0.006932f
C4563 vdd.n3286 gnd 0.006932f
C4564 vdd.n3287 gnd 0.006932f
C4565 vdd.n3288 gnd 0.006932f
C4566 vdd.n3289 gnd 0.006932f
C4567 vdd.n3291 gnd 0.006932f
C4568 vdd.n3292 gnd 0.006932f
C4569 vdd.n3293 gnd 0.006932f
C4570 vdd.n3294 gnd 0.006932f
C4571 vdd.n3295 gnd 0.006932f
C4572 vdd.n3296 gnd 0.006932f
C4573 vdd.n3298 gnd 0.006932f
C4574 vdd.n3299 gnd 0.006932f
C4575 vdd.n3300 gnd 0.006932f
C4576 vdd.n3302 gnd 0.006932f
C4577 vdd.n3303 gnd 0.006932f
C4578 vdd.n3304 gnd 0.006932f
C4579 vdd.n3305 gnd 0.006932f
C4580 vdd.n3306 gnd 0.006932f
C4581 vdd.n3307 gnd 0.006932f
C4582 vdd.n3309 gnd 0.006932f
C4583 vdd.n3310 gnd 0.006932f
C4584 vdd.n3311 gnd 0.006932f
C4585 vdd.n3312 gnd 0.006932f
C4586 vdd.n3313 gnd 0.006932f
C4587 vdd.n3314 gnd 0.006932f
C4588 vdd.n3316 gnd 0.006932f
C4589 vdd.n3317 gnd 0.006932f
C4590 vdd.n3318 gnd 0.006932f
C4591 vdd.n3319 gnd 0.006932f
C4592 vdd.n3320 gnd 0.006932f
C4593 vdd.n3321 gnd 0.006932f
C4594 vdd.n3323 gnd 0.006932f
C4595 vdd.n3324 gnd 0.006932f
C4596 vdd.n3326 gnd 0.006932f
C4597 vdd.n3327 gnd 0.006932f
C4598 vdd.n3328 gnd 0.01574f
C4599 vdd.n3329 gnd 0.014843f
C4600 vdd.n3330 gnd 0.014843f
C4601 vdd.n3331 gnd 0.958462f
C4602 vdd.n3332 gnd 0.014843f
C4603 vdd.n3333 gnd 0.01574f
C4604 vdd.n3334 gnd 0.014843f
C4605 vdd.n3335 gnd 0.006932f
C4606 vdd.n3336 gnd 0.005352f
C4607 vdd.n3337 gnd 0.006932f
C4608 vdd.n3339 gnd 0.006932f
C4609 vdd.n3340 gnd 0.006932f
C4610 vdd.n3341 gnd 0.006932f
C4611 vdd.n3342 gnd 0.006932f
C4612 vdd.n3343 gnd 0.006932f
C4613 vdd.n3344 gnd 0.006932f
C4614 vdd.n3346 gnd 0.006932f
C4615 vdd.n3347 gnd 0.006932f
C4616 vdd.n3348 gnd 0.006932f
C4617 vdd.n3349 gnd 0.006932f
C4618 vdd.n3350 gnd 0.006932f
C4619 vdd.n3351 gnd 0.006932f
C4620 vdd.n3353 gnd 0.006932f
C4621 vdd.n3354 gnd 0.006932f
C4622 vdd.n3355 gnd 0.006932f
C4623 vdd.n3356 gnd 0.006932f
C4624 vdd.n3357 gnd 0.006932f
C4625 vdd.n3358 gnd 0.006932f
C4626 vdd.n3360 gnd 0.006932f
C4627 vdd.n3361 gnd 0.006932f
C4628 vdd.n3363 gnd 0.006932f
C4629 vdd.n3364 gnd 0.042805f
C4630 vdd.n3365 gnd 1.08612f
C4631 vdd.n3367 gnd 0.004308f
C4632 vdd.n3368 gnd 0.008205f
C4633 vdd.n3369 gnd 0.010194f
C4634 vdd.n3370 gnd 0.010194f
C4635 vdd.n3371 gnd 0.008205f
C4636 vdd.n3372 gnd 0.008205f
C4637 vdd.n3373 gnd 0.010194f
C4638 vdd.n3374 gnd 0.010194f
C4639 vdd.n3375 gnd 0.008205f
C4640 vdd.n3376 gnd 0.008205f
C4641 vdd.n3377 gnd 0.010194f
C4642 vdd.n3378 gnd 0.010194f
C4643 vdd.n3379 gnd 0.008205f
C4644 vdd.n3380 gnd 0.008205f
C4645 vdd.n3381 gnd 0.010194f
C4646 vdd.n3382 gnd 0.010194f
C4647 vdd.n3383 gnd 0.008205f
C4648 vdd.n3384 gnd 0.008205f
C4649 vdd.n3385 gnd 0.010194f
C4650 vdd.n3386 gnd 0.010194f
C4651 vdd.n3387 gnd 0.008205f
C4652 vdd.n3388 gnd 0.008205f
C4653 vdd.n3389 gnd 0.010194f
C4654 vdd.n3390 gnd 0.010194f
C4655 vdd.n3391 gnd 0.008205f
C4656 vdd.n3392 gnd 0.008205f
C4657 vdd.n3393 gnd 0.010194f
C4658 vdd.n3394 gnd 0.010194f
C4659 vdd.n3395 gnd 0.008205f
C4660 vdd.n3396 gnd 0.008205f
C4661 vdd.n3397 gnd 0.010194f
C4662 vdd.n3398 gnd 0.010194f
C4663 vdd.n3399 gnd 0.008205f
C4664 vdd.n3400 gnd 0.008205f
C4665 vdd.n3401 gnd 0.010194f
C4666 vdd.n3402 gnd 0.010194f
C4667 vdd.n3403 gnd 0.008205f
C4668 vdd.n3404 gnd 0.010194f
C4669 vdd.n3405 gnd 0.010194f
C4670 vdd.n3406 gnd 0.008205f
C4671 vdd.n3407 gnd 0.010194f
C4672 vdd.n3408 gnd 0.010194f
C4673 vdd.n3409 gnd 0.010194f
C4674 vdd.n3410 gnd 0.016739f
C4675 vdd.n3411 gnd 0.010194f
C4676 vdd.n3412 gnd 0.010194f
C4677 vdd.n3413 gnd 0.00558f
C4678 vdd.n3414 gnd 0.008205f
C4679 vdd.n3415 gnd 0.010194f
C4680 vdd.n3416 gnd 0.010194f
C4681 vdd.n3417 gnd 0.008205f
C4682 vdd.n3418 gnd 0.008205f
C4683 vdd.n3419 gnd 0.010194f
C4684 vdd.n3420 gnd 0.010194f
C4685 vdd.n3421 gnd 0.008205f
C4686 vdd.n3422 gnd 0.008205f
C4687 vdd.n3423 gnd 0.010194f
C4688 vdd.n3424 gnd 0.010194f
C4689 vdd.n3425 gnd 0.008205f
C4690 vdd.n3426 gnd 0.008205f
C4691 vdd.n3427 gnd 0.010194f
C4692 vdd.n3428 gnd 0.010194f
C4693 vdd.n3429 gnd 0.008205f
C4694 vdd.n3430 gnd 0.008205f
C4695 vdd.n3431 gnd 0.010194f
C4696 vdd.n3432 gnd 0.010194f
C4697 vdd.n3433 gnd 0.008205f
C4698 vdd.n3434 gnd 0.008205f
C4699 vdd.n3435 gnd 0.010194f
C4700 vdd.n3436 gnd 0.010194f
C4701 vdd.n3437 gnd 0.008205f
C4702 vdd.n3438 gnd 0.008205f
C4703 vdd.n3439 gnd 0.010194f
C4704 vdd.n3440 gnd 0.010194f
C4705 vdd.n3441 gnd 0.008205f
C4706 vdd.n3442 gnd 0.008205f
C4707 vdd.n3443 gnd 0.010194f
C4708 vdd.n3444 gnd 0.010194f
C4709 vdd.n3445 gnd 0.008205f
C4710 vdd.n3446 gnd 0.008205f
C4711 vdd.n3447 gnd 0.010194f
C4712 vdd.n3448 gnd 0.010194f
C4713 vdd.n3449 gnd 0.008205f
C4714 vdd.n3450 gnd 0.010194f
C4715 vdd.n3451 gnd 0.010194f
C4716 vdd.n3452 gnd 0.008205f
C4717 vdd.n3453 gnd 0.010194f
C4718 vdd.n3454 gnd 0.010194f
C4719 vdd.n3455 gnd 0.010194f
C4720 vdd.t133 gnd 0.125416f
C4721 vdd.t134 gnd 0.134036f
C4722 vdd.t132 gnd 0.163792f
C4723 vdd.n3456 gnd 0.209958f
C4724 vdd.n3457 gnd 0.176403f
C4725 vdd.n3458 gnd 0.016739f
C4726 vdd.n3459 gnd 0.010194f
C4727 vdd.n3460 gnd 0.010194f
C4728 vdd.n3461 gnd 0.006851f
C4729 vdd.n3462 gnd 0.008205f
C4730 vdd.n3463 gnd 0.010194f
C4731 vdd.n3464 gnd 0.010194f
C4732 vdd.n3465 gnd 0.008205f
C4733 vdd.n3466 gnd 0.008205f
C4734 vdd.n3467 gnd 0.010194f
C4735 vdd.n3468 gnd 0.010194f
C4736 vdd.n3469 gnd 0.008205f
C4737 vdd.n3470 gnd 0.008205f
C4738 vdd.n3471 gnd 0.010194f
C4739 vdd.n3472 gnd 0.010194f
C4740 vdd.n3473 gnd 0.008205f
C4741 vdd.n3474 gnd 0.008205f
C4742 vdd.n3475 gnd 0.010194f
C4743 vdd.n3476 gnd 0.010194f
C4744 vdd.n3477 gnd 0.008205f
C4745 vdd.n3478 gnd 0.008205f
C4746 vdd.n3479 gnd 0.010194f
C4747 vdd.n3480 gnd 0.010194f
C4748 vdd.n3481 gnd 0.008205f
C4749 vdd.n3482 gnd 0.008205f
C4750 vdd.n3483 gnd 0.010194f
C4751 vdd.n3484 gnd 0.010194f
C4752 vdd.n3485 gnd 0.008205f
C4753 vdd.n3486 gnd 0.008205f
C4754 vdd.n3488 gnd 1.08612f
C4755 vdd.n3490 gnd 0.008205f
C4756 vdd.n3491 gnd 0.008205f
C4757 vdd.n3492 gnd 0.00681f
C4758 vdd.n3493 gnd 0.025189f
C4759 vdd.n3495 gnd 12.7205f
C4760 vdd.n3496 gnd 0.025189f
C4761 vdd.n3497 gnd 0.003897f
C4762 vdd.n3498 gnd 0.025189f
C4763 vdd.n3499 gnd 0.024661f
C4764 vdd.n3500 gnd 0.010194f
C4765 vdd.n3501 gnd 0.008205f
C4766 vdd.n3502 gnd 0.010194f
C4767 vdd.n3503 gnd 0.630293f
C4768 vdd.n3504 gnd 0.010194f
C4769 vdd.n3505 gnd 0.008205f
C4770 vdd.n3506 gnd 0.010194f
C4771 vdd.n3507 gnd 0.010194f
C4772 vdd.n3508 gnd 0.010194f
C4773 vdd.n3509 gnd 0.008205f
C4774 vdd.n3510 gnd 0.010194f
C4775 vdd.n3511 gnd 1.04181f
C4776 vdd.n3512 gnd 0.010194f
C4777 vdd.n3513 gnd 0.008205f
C4778 vdd.n3514 gnd 0.010194f
C4779 vdd.n3515 gnd 0.010194f
C4780 vdd.n3516 gnd 0.010194f
C4781 vdd.n3517 gnd 0.008205f
C4782 vdd.n3518 gnd 0.010194f
C4783 vdd.n3519 gnd 0.671965f
C4784 vdd.n3520 gnd 0.713638f
C4785 vdd.n3521 gnd 0.010194f
C4786 vdd.n3522 gnd 0.008205f
C4787 vdd.n3523 gnd 0.010194f
C4788 vdd.n3524 gnd 0.010194f
C4789 vdd.n3525 gnd 0.010194f
C4790 vdd.n3526 gnd 0.008205f
C4791 vdd.n3527 gnd 0.010194f
C4792 vdd.n3528 gnd 0.864699f
C4793 vdd.n3529 gnd 0.010194f
C4794 vdd.n3530 gnd 0.008205f
C4795 vdd.n3531 gnd 0.010194f
C4796 vdd.n3532 gnd 0.010194f
C4797 vdd.n3533 gnd 0.010194f
C4798 vdd.n3534 gnd 0.008205f
C4799 vdd.n3535 gnd 0.010194f
C4800 vdd.t54 gnd 0.520903f
C4801 vdd.n3536 gnd 0.838654f
C4802 vdd.n3537 gnd 0.010194f
C4803 vdd.n3538 gnd 0.008205f
C4804 vdd.n3539 gnd 0.010194f
C4805 vdd.n3540 gnd 0.010194f
C4806 vdd.n3541 gnd 0.010194f
C4807 vdd.n3542 gnd 0.008205f
C4808 vdd.n3543 gnd 0.010194f
C4809 vdd.n3544 gnd 0.661547f
C4810 vdd.n3545 gnd 0.010194f
C4811 vdd.n3546 gnd 0.008205f
C4812 vdd.n3547 gnd 0.010194f
C4813 vdd.n3548 gnd 0.010194f
C4814 vdd.n3549 gnd 0.010194f
C4815 vdd.n3550 gnd 0.008205f
C4816 vdd.n3551 gnd 0.010194f
C4817 vdd.n3552 gnd 0.828236f
C4818 vdd.n3553 gnd 0.557367f
C4819 vdd.n3554 gnd 0.010194f
C4820 vdd.n3555 gnd 0.008205f
C4821 vdd.n3556 gnd 0.010194f
C4822 vdd.n3557 gnd 0.010194f
C4823 vdd.n3558 gnd 0.010194f
C4824 vdd.n3559 gnd 0.008205f
C4825 vdd.n3560 gnd 0.010194f
C4826 vdd.n3561 gnd 0.734474f
C4827 vdd.n3562 gnd 0.010194f
C4828 vdd.n3563 gnd 0.008205f
C4829 vdd.n3564 gnd 0.010194f
C4830 vdd.n3565 gnd 0.010194f
C4831 vdd.n3566 gnd 0.010194f
C4832 vdd.n3567 gnd 0.010194f
C4833 vdd.n3568 gnd 0.010194f
C4834 vdd.n3569 gnd 0.008205f
C4835 vdd.n3570 gnd 0.008205f
C4836 vdd.n3571 gnd 0.010194f
C4837 vdd.t159 gnd 0.520903f
C4838 vdd.n3572 gnd 0.864699f
C4839 vdd.n3573 gnd 0.010194f
C4840 vdd.n3574 gnd 0.008205f
C4841 vdd.n3575 gnd 0.010194f
C4842 vdd.n3576 gnd 0.010194f
C4843 vdd.n3577 gnd 0.010194f
C4844 vdd.n3578 gnd 0.008205f
C4845 vdd.n3579 gnd 0.010194f
C4846 vdd.n3580 gnd 0.817818f
C4847 vdd.n3581 gnd 0.010194f
C4848 vdd.n3582 gnd 0.010194f
C4849 vdd.n3583 gnd 0.008205f
C4850 vdd.n3584 gnd 0.008205f
C4851 vdd.n3585 gnd 0.010194f
C4852 vdd.n3586 gnd 0.010194f
C4853 vdd.n3587 gnd 0.010194f
C4854 vdd.n3588 gnd 0.008205f
C4855 vdd.n3589 gnd 0.010194f
C4856 vdd.n3590 gnd 0.008205f
C4857 vdd.n3591 gnd 0.008205f
C4858 vdd.n3592 gnd 0.010194f
C4859 vdd.n3593 gnd 0.010194f
C4860 vdd.n3594 gnd 0.010194f
C4861 vdd.n3595 gnd 0.008205f
C4862 vdd.n3596 gnd 0.010194f
C4863 vdd.n3597 gnd 0.008205f
C4864 vdd.n3598 gnd 0.008205f
C4865 vdd.n3599 gnd 0.010194f
C4866 vdd.n3600 gnd 0.010194f
C4867 vdd.n3601 gnd 0.010194f
C4868 vdd.n3602 gnd 0.008205f
C4869 vdd.n3603 gnd 0.864699f
C4870 vdd.n3604 gnd 0.010194f
C4871 vdd.n3605 gnd 0.008205f
C4872 vdd.n3606 gnd 0.008205f
C4873 vdd.n3607 gnd 0.010194f
C4874 vdd.n3608 gnd 0.010194f
C4875 vdd.n3609 gnd 0.010194f
C4876 vdd.n3610 gnd 0.008205f
C4877 vdd.n3611 gnd 0.010194f
C4878 vdd.n3612 gnd 0.008205f
C4879 vdd.n3613 gnd 0.008205f
C4880 vdd.n3614 gnd 0.010194f
C4881 vdd.n3615 gnd 0.010194f
C4882 vdd.n3616 gnd 0.010194f
C4883 vdd.n3617 gnd 0.008205f
C4884 vdd.n3618 gnd 0.010194f
C4885 vdd.n3619 gnd 0.008205f
C4886 vdd.n3620 gnd 0.00681f
C4887 vdd.n3621 gnd 0.024661f
C4888 vdd.n3622 gnd 0.025189f
C4889 vdd.n3623 gnd 0.003897f
C4890 vdd.n3624 gnd 0.025189f
C4891 vdd.n3626 gnd 2.46908f
C4892 vdd.n3627 gnd 1.53666f
C4893 vdd.n3628 gnd 0.024661f
C4894 vdd.n3629 gnd 0.00681f
C4895 vdd.n3630 gnd 0.008205f
C4896 vdd.n3631 gnd 0.008205f
C4897 vdd.n3632 gnd 0.010194f
C4898 vdd.n3633 gnd 1.04181f
C4899 vdd.n3634 gnd 1.04181f
C4900 vdd.n3635 gnd 0.953253f
C4901 vdd.n3636 gnd 0.010194f
C4902 vdd.n3637 gnd 0.008205f
C4903 vdd.n3638 gnd 0.008205f
C4904 vdd.n3639 gnd 0.008205f
C4905 vdd.n3640 gnd 0.010194f
C4906 vdd.n3641 gnd 0.776146f
C4907 vdd.t186 gnd 0.520903f
C4908 vdd.n3642 gnd 0.786564f
C4909 vdd.n3643 gnd 0.599039f
C4910 vdd.n3644 gnd 0.010194f
C4911 vdd.n3645 gnd 0.008205f
C4912 vdd.n3646 gnd 0.008205f
C4913 vdd.n3647 gnd 0.008205f
C4914 vdd.n3648 gnd 0.010194f
C4915 vdd.n3649 gnd 0.619875f
C4916 vdd.n3650 gnd 0.765728f
C4917 vdd.t6 gnd 0.520903f
C4918 vdd.n3651 gnd 0.796982f
C4919 vdd.n3652 gnd 0.010194f
C4920 vdd.n3653 gnd 0.008205f
C4921 vdd.n3654 gnd 0.008205f
C4922 vdd.n3655 gnd 0.008205f
C4923 vdd.n3656 gnd 0.010194f
C4924 vdd.n3657 gnd 0.864699f
C4925 vdd.t51 gnd 0.520903f
C4926 vdd.n3658 gnd 0.630293f
C4927 vdd.n3659 gnd 0.75531f
C4928 vdd.n3660 gnd 0.010194f
C4929 vdd.n3661 gnd 0.008205f
C4930 vdd.n3662 gnd 0.008205f
C4931 vdd.n3663 gnd 0.008205f
C4932 vdd.n3664 gnd 0.010194f
C4933 vdd.n3665 gnd 0.578203f
C4934 vdd.t39 gnd 0.520903f
C4935 vdd.n3666 gnd 0.864699f
C4936 vdd.t70 gnd 0.520903f
C4937 vdd.n3667 gnd 0.640711f
C4938 vdd.n3668 gnd 0.010194f
C4939 vdd.n3669 gnd 0.008205f
C4940 vdd.n3670 gnd 0.007835f
C4941 vdd.n3671 gnd 0.601297f
C4942 vdd.n3672 gnd 2.97728f
C4943 a_n2982_13878.n0 gnd 2.69774f
C4944 a_n2982_13878.n1 gnd 3.89736f
C4945 a_n2982_13878.n2 gnd 3.76836f
C4946 a_n2982_13878.n3 gnd 3.09829f
C4947 a_n2982_13878.n4 gnd 0.208192f
C4948 a_n2982_13878.n5 gnd 0.208192f
C4949 a_n2982_13878.n6 gnd 0.838872f
C4950 a_n2982_13878.n7 gnd 0.208192f
C4951 a_n2982_13878.n8 gnd 0.272971f
C4952 a_n2982_13878.n9 gnd 0.965983f
C4953 a_n2982_13878.n10 gnd 0.208192f
C4954 a_n2982_13878.n11 gnd 0.208192f
C4955 a_n2982_13878.n12 gnd 0.474155f
C4956 a_n2982_13878.n13 gnd 0.208192f
C4957 a_n2982_13878.n14 gnd 0.272971f
C4958 a_n2982_13878.n15 gnd 0.898614f
C4959 a_n2982_13878.n16 gnd 0.19754f
C4960 a_n2982_13878.n17 gnd 0.145492f
C4961 a_n2982_13878.n18 gnd 0.228667f
C4962 a_n2982_13878.n19 gnd 0.176619f
C4963 a_n2982_13878.n20 gnd 0.19754f
C4964 a_n2982_13878.n21 gnd 1.31591f
C4965 a_n2982_13878.n22 gnd 0.145492f
C4966 a_n2982_13878.n23 gnd 0.950662f
C4967 a_n2982_13878.n24 gnd 0.208192f
C4968 a_n2982_13878.n25 gnd 0.732765f
C4969 a_n2982_13878.n26 gnd 0.208192f
C4970 a_n2982_13878.n27 gnd 0.208192f
C4971 a_n2982_13878.n28 gnd 0.474155f
C4972 a_n2982_13878.n29 gnd 0.272971f
C4973 a_n2982_13878.n30 gnd 0.208192f
C4974 a_n2982_13878.n31 gnd 0.526203f
C4975 a_n2982_13878.n32 gnd 0.208192f
C4976 a_n2982_13878.n33 gnd 0.208192f
C4977 a_n2982_13878.n34 gnd 0.926304f
C4978 a_n2982_13878.n35 gnd 0.272971f
C4979 a_n2982_13878.n36 gnd 1.71402f
C4980 a_n2982_13878.n37 gnd 1.15494f
C4981 a_n2982_13878.n38 gnd 2.30668f
C4982 a_n2982_13878.n39 gnd 2.10894f
C4983 a_n2982_13878.n40 gnd 1.15494f
C4984 a_n2982_13878.n41 gnd 1.71402f
C4985 a_n2982_13878.n42 gnd 0.008354f
C4986 a_n2982_13878.n43 gnd 4.03e-19
C4987 a_n2982_13878.n45 gnd 0.008061f
C4988 a_n2982_13878.n46 gnd 0.011721f
C4989 a_n2982_13878.n47 gnd 0.007754f
C4990 a_n2982_13878.n49 gnd 0.276148f
C4991 a_n2982_13878.n50 gnd 0.008354f
C4992 a_n2982_13878.n51 gnd 4.03e-19
C4993 a_n2982_13878.n53 gnd 0.008061f
C4994 a_n2982_13878.n54 gnd 0.011721f
C4995 a_n2982_13878.n55 gnd 0.007754f
C4996 a_n2982_13878.n57 gnd 0.276148f
C4997 a_n2982_13878.n58 gnd 0.008061f
C4998 a_n2982_13878.n59 gnd 0.275022f
C4999 a_n2982_13878.n60 gnd 0.008061f
C5000 a_n2982_13878.n61 gnd 0.275022f
C5001 a_n2982_13878.n62 gnd 0.008061f
C5002 a_n2982_13878.n63 gnd 0.275022f
C5003 a_n2982_13878.n64 gnd 0.008061f
C5004 a_n2982_13878.n65 gnd 0.275022f
C5005 a_n2982_13878.n66 gnd 0.008354f
C5006 a_n2982_13878.n67 gnd 4.03e-19
C5007 a_n2982_13878.n69 gnd 0.008061f
C5008 a_n2982_13878.n70 gnd 0.011721f
C5009 a_n2982_13878.n71 gnd 0.007754f
C5010 a_n2982_13878.n73 gnd 0.276148f
C5011 a_n2982_13878.n74 gnd 0.008354f
C5012 a_n2982_13878.n75 gnd 4.03e-19
C5013 a_n2982_13878.n77 gnd 0.008061f
C5014 a_n2982_13878.n78 gnd 0.011721f
C5015 a_n2982_13878.n79 gnd 0.007754f
C5016 a_n2982_13878.n81 gnd 0.276148f
C5017 a_n2982_13878.t38 gnd 0.144404f
C5018 a_n2982_13878.t35 gnd 0.685683f
C5019 a_n2982_13878.t59 gnd 0.671699f
C5020 a_n2982_13878.t17 gnd 0.671699f
C5021 a_n2982_13878.t45 gnd 0.671699f
C5022 a_n2982_13878.n82 gnd 0.295189f
C5023 a_n2982_13878.t61 gnd 0.671699f
C5024 a_n2982_13878.t43 gnd 0.671699f
C5025 a_n2982_13878.t27 gnd 0.671699f
C5026 a_n2982_13878.n83 gnd 0.291571f
C5027 a_n2982_13878.t37 gnd 0.671699f
C5028 a_n2982_13878.t15 gnd 0.671699f
C5029 a_n2982_13878.t29 gnd 0.671699f
C5030 a_n2982_13878.n84 gnd 0.295307f
C5031 a_n2982_13878.t53 gnd 0.671699f
C5032 a_n2982_13878.t41 gnd 0.682505f
C5033 a_n2982_13878.t2 gnd 0.112315f
C5034 a_n2982_13878.t8 gnd 0.112315f
C5035 a_n2982_13878.n85 gnd 0.995376f
C5036 a_n2982_13878.t5 gnd 0.112315f
C5037 a_n2982_13878.t7 gnd 0.112315f
C5038 a_n2982_13878.n86 gnd 0.99245f
C5039 a_n2982_13878.t9 gnd 0.112315f
C5040 a_n2982_13878.t63 gnd 0.112315f
C5041 a_n2982_13878.n87 gnd 0.995376f
C5042 a_n2982_13878.t13 gnd 0.112315f
C5043 a_n2982_13878.t14 gnd 0.112315f
C5044 a_n2982_13878.n88 gnd 0.99245f
C5045 a_n2982_13878.t0 gnd 0.112315f
C5046 a_n2982_13878.t1 gnd 0.112315f
C5047 a_n2982_13878.n89 gnd 0.992451f
C5048 a_n2982_13878.t10 gnd 0.112315f
C5049 a_n2982_13878.t11 gnd 0.112315f
C5050 a_n2982_13878.n90 gnd 0.992451f
C5051 a_n2982_13878.t3 gnd 0.112315f
C5052 a_n2982_13878.t4 gnd 0.112315f
C5053 a_n2982_13878.n91 gnd 0.995377f
C5054 a_n2982_13878.t12 gnd 0.112315f
C5055 a_n2982_13878.t6 gnd 0.112315f
C5056 a_n2982_13878.n92 gnd 0.992451f
C5057 a_n2982_13878.t102 gnd 0.685683f
C5058 a_n2982_13878.t79 gnd 0.671699f
C5059 a_n2982_13878.t84 gnd 0.671699f
C5060 a_n2982_13878.t72 gnd 0.671699f
C5061 a_n2982_13878.n93 gnd 0.295189f
C5062 a_n2982_13878.t89 gnd 0.671699f
C5063 a_n2982_13878.t98 gnd 0.671699f
C5064 a_n2982_13878.t99 gnd 0.671699f
C5065 a_n2982_13878.n94 gnd 0.291571f
C5066 a_n2982_13878.t66 gnd 0.671699f
C5067 a_n2982_13878.t81 gnd 0.671699f
C5068 a_n2982_13878.t69 gnd 0.671699f
C5069 a_n2982_13878.n95 gnd 0.295307f
C5070 a_n2982_13878.t76 gnd 0.671699f
C5071 a_n2982_13878.t95 gnd 0.682505f
C5072 a_n2982_13878.t58 gnd 1.35213f
C5073 a_n2982_13878.t22 gnd 0.144404f
C5074 a_n2982_13878.t40 gnd 0.144404f
C5075 a_n2982_13878.n96 gnd 1.01718f
C5076 a_n2982_13878.t52 gnd 0.144404f
C5077 a_n2982_13878.t26 gnd 0.144404f
C5078 a_n2982_13878.n97 gnd 1.01718f
C5079 a_n2982_13878.t20 gnd 0.144404f
C5080 a_n2982_13878.t48 gnd 0.144404f
C5081 a_n2982_13878.n98 gnd 1.01718f
C5082 a_n2982_13878.t50 gnd 0.144404f
C5083 a_n2982_13878.t24 gnd 0.144404f
C5084 a_n2982_13878.n99 gnd 1.01718f
C5085 a_n2982_13878.t32 gnd 0.144404f
C5086 a_n2982_13878.t34 gnd 0.144404f
C5087 a_n2982_13878.n100 gnd 1.01718f
C5088 a_n2982_13878.t56 gnd 1.34943f
C5089 a_n2982_13878.t31 gnd 0.671699f
C5090 a_n2982_13878.n101 gnd 0.295307f
C5091 a_n2982_13878.t33 gnd 0.671699f
C5092 a_n2982_13878.t49 gnd 0.671699f
C5093 a_n2982_13878.n102 gnd 0.286437f
C5094 a_n2982_13878.t25 gnd 0.671699f
C5095 a_n2982_13878.n103 gnd 0.297845f
C5096 a_n2982_13878.t19 gnd 0.671699f
C5097 a_n2982_13878.t39 gnd 0.671699f
C5098 a_n2982_13878.n104 gnd 0.29125f
C5099 a_n2982_13878.t57 gnd 0.685683f
C5100 a_n2982_13878.t78 gnd 0.671699f
C5101 a_n2982_13878.n105 gnd 0.295307f
C5102 a_n2982_13878.t88 gnd 0.671699f
C5103 a_n2982_13878.t93 gnd 0.671699f
C5104 a_n2982_13878.n106 gnd 0.286437f
C5105 a_n2982_13878.t97 gnd 0.671699f
C5106 a_n2982_13878.n107 gnd 0.297845f
C5107 a_n2982_13878.t68 gnd 0.671699f
C5108 a_n2982_13878.t71 gnd 0.671699f
C5109 a_n2982_13878.n108 gnd 0.29125f
C5110 a_n2982_13878.t101 gnd 0.685683f
C5111 a_n2982_13878.t70 gnd 0.671699f
C5112 a_n2982_13878.n109 gnd 0.297409f
C5113 a_n2982_13878.t96 gnd 0.671699f
C5114 a_n2982_13878.n110 gnd 0.295189f
C5115 a_n2982_13878.n111 gnd 0.295322f
C5116 a_n2982_13878.t92 gnd 0.671699f
C5117 a_n2982_13878.n112 gnd 0.291571f
C5118 a_n2982_13878.t65 gnd 0.671699f
C5119 a_n2982_13878.n113 gnd 0.291822f
C5120 a_n2982_13878.n114 gnd 0.297409f
C5121 a_n2982_13878.t67 gnd 0.682505f
C5122 a_n2982_13878.t21 gnd 0.671699f
C5123 a_n2982_13878.n115 gnd 0.297409f
C5124 a_n2982_13878.t51 gnd 0.671699f
C5125 a_n2982_13878.n116 gnd 0.295189f
C5126 a_n2982_13878.n117 gnd 0.295322f
C5127 a_n2982_13878.t47 gnd 0.671699f
C5128 a_n2982_13878.n118 gnd 0.291571f
C5129 a_n2982_13878.t23 gnd 0.671699f
C5130 a_n2982_13878.n119 gnd 0.291822f
C5131 a_n2982_13878.n120 gnd 0.297409f
C5132 a_n2982_13878.t55 gnd 0.682505f
C5133 a_n2982_13878.n121 gnd 1.30049f
C5134 a_n2982_13878.t75 gnd 0.671699f
C5135 a_n2982_13878.n122 gnd 0.291571f
C5136 a_n2982_13878.t83 gnd 0.671699f
C5137 a_n2982_13878.n123 gnd 0.291571f
C5138 a_n2982_13878.t73 gnd 0.671699f
C5139 a_n2982_13878.n124 gnd 0.291571f
C5140 a_n2982_13878.t87 gnd 0.671699f
C5141 a_n2982_13878.n125 gnd 0.291571f
C5142 a_n2982_13878.t77 gnd 0.671699f
C5143 a_n2982_13878.n126 gnd 0.286276f
C5144 a_n2982_13878.t103 gnd 0.671699f
C5145 a_n2982_13878.n127 gnd 0.295322f
C5146 a_n2982_13878.t80 gnd 0.682954f
C5147 a_n2982_13878.t90 gnd 0.671699f
C5148 a_n2982_13878.n128 gnd 0.286276f
C5149 a_n2982_13878.t74 gnd 0.671699f
C5150 a_n2982_13878.n129 gnd 0.295322f
C5151 a_n2982_13878.t85 gnd 0.682954f
C5152 a_n2982_13878.t94 gnd 0.671699f
C5153 a_n2982_13878.n130 gnd 0.286276f
C5154 a_n2982_13878.t82 gnd 0.671699f
C5155 a_n2982_13878.n131 gnd 0.295322f
C5156 a_n2982_13878.t100 gnd 0.682954f
C5157 a_n2982_13878.t86 gnd 0.671699f
C5158 a_n2982_13878.n132 gnd 0.286276f
C5159 a_n2982_13878.t64 gnd 0.671699f
C5160 a_n2982_13878.n133 gnd 0.295322f
C5161 a_n2982_13878.t91 gnd 0.682954f
C5162 a_n2982_13878.n134 gnd 1.63586f
C5163 a_n2982_13878.n135 gnd 0.297409f
C5164 a_n2982_13878.n136 gnd 0.291822f
C5165 a_n2982_13878.n137 gnd 0.286437f
C5166 a_n2982_13878.n138 gnd 0.295322f
C5167 a_n2982_13878.n139 gnd 0.297845f
C5168 a_n2982_13878.n140 gnd 0.29125f
C5169 a_n2982_13878.n141 gnd 0.297409f
C5170 a_n2982_13878.n142 gnd 0.297409f
C5171 a_n2982_13878.n143 gnd 0.291822f
C5172 a_n2982_13878.n144 gnd 0.286437f
C5173 a_n2982_13878.n145 gnd 0.295322f
C5174 a_n2982_13878.n146 gnd 0.297845f
C5175 a_n2982_13878.n147 gnd 0.29125f
C5176 a_n2982_13878.n148 gnd 0.297409f
C5177 a_n2982_13878.n149 gnd 0.988833f
C5178 a_n2982_13878.t36 gnd 1.34944f
C5179 a_n2982_13878.t60 gnd 0.144404f
C5180 a_n2982_13878.t18 gnd 0.144404f
C5181 a_n2982_13878.n150 gnd 1.01718f
C5182 a_n2982_13878.t46 gnd 0.144404f
C5183 a_n2982_13878.t62 gnd 0.144404f
C5184 a_n2982_13878.n151 gnd 1.01718f
C5185 a_n2982_13878.t44 gnd 0.144404f
C5186 a_n2982_13878.t28 gnd 0.144404f
C5187 a_n2982_13878.n152 gnd 1.01718f
C5188 a_n2982_13878.t42 gnd 1.35213f
C5189 a_n2982_13878.t30 gnd 0.144404f
C5190 a_n2982_13878.t54 gnd 0.144404f
C5191 a_n2982_13878.n153 gnd 1.01718f
C5192 a_n2982_13878.n154 gnd 1.01719f
C5193 a_n2982_13878.t16 gnd 0.144404f
C5194 CSoutput.n0 gnd 0.048358f
C5195 CSoutput.t186 gnd 0.319878f
C5196 CSoutput.n1 gnd 0.144441f
C5197 CSoutput.n2 gnd 0.048358f
C5198 CSoutput.t183 gnd 0.319878f
C5199 CSoutput.n3 gnd 0.038328f
C5200 CSoutput.n4 gnd 0.048358f
C5201 CSoutput.t173 gnd 0.319878f
C5202 CSoutput.n5 gnd 0.03305f
C5203 CSoutput.n6 gnd 0.048358f
C5204 CSoutput.t181 gnd 0.319878f
C5205 CSoutput.t168 gnd 0.319878f
C5206 CSoutput.n7 gnd 0.142867f
C5207 CSoutput.n8 gnd 0.048358f
C5208 CSoutput.t172 gnd 0.319878f
C5209 CSoutput.n9 gnd 0.031512f
C5210 CSoutput.n10 gnd 0.048358f
C5211 CSoutput.t176 gnd 0.319878f
C5212 CSoutput.t182 gnd 0.319878f
C5213 CSoutput.n11 gnd 0.142867f
C5214 CSoutput.n12 gnd 0.048358f
C5215 CSoutput.t188 gnd 0.319878f
C5216 CSoutput.n13 gnd 0.03305f
C5217 CSoutput.n14 gnd 0.048358f
C5218 CSoutput.t174 gnd 0.319878f
C5219 CSoutput.t180 gnd 0.319878f
C5220 CSoutput.n15 gnd 0.142867f
C5221 CSoutput.n16 gnd 0.048358f
C5222 CSoutput.t187 gnd 0.319878f
C5223 CSoutput.n17 gnd 0.035299f
C5224 CSoutput.t175 gnd 0.382263f
C5225 CSoutput.t184 gnd 0.319878f
C5226 CSoutput.n18 gnd 0.182385f
C5227 CSoutput.n19 gnd 0.176977f
C5228 CSoutput.n20 gnd 0.205314f
C5229 CSoutput.n21 gnd 0.048358f
C5230 CSoutput.n22 gnd 0.04036f
C5231 CSoutput.n23 gnd 0.142867f
C5232 CSoutput.n24 gnd 0.038906f
C5233 CSoutput.n25 gnd 0.038328f
C5234 CSoutput.n26 gnd 0.048358f
C5235 CSoutput.n27 gnd 0.048358f
C5236 CSoutput.n28 gnd 0.04005f
C5237 CSoutput.n29 gnd 0.034003f
C5238 CSoutput.n30 gnd 0.146047f
C5239 CSoutput.n31 gnd 0.034472f
C5240 CSoutput.n32 gnd 0.048358f
C5241 CSoutput.n33 gnd 0.048358f
C5242 CSoutput.n34 gnd 0.048358f
C5243 CSoutput.n35 gnd 0.039623f
C5244 CSoutput.n36 gnd 0.142867f
C5245 CSoutput.n37 gnd 0.037894f
C5246 CSoutput.n38 gnd 0.03934f
C5247 CSoutput.n39 gnd 0.048358f
C5248 CSoutput.n40 gnd 0.048358f
C5249 CSoutput.n41 gnd 0.040352f
C5250 CSoutput.n42 gnd 0.036882f
C5251 CSoutput.n43 gnd 0.142867f
C5252 CSoutput.n44 gnd 0.037817f
C5253 CSoutput.n45 gnd 0.048358f
C5254 CSoutput.n46 gnd 0.048358f
C5255 CSoutput.n47 gnd 0.048358f
C5256 CSoutput.n48 gnd 0.037817f
C5257 CSoutput.n49 gnd 0.142867f
C5258 CSoutput.n50 gnd 0.036882f
C5259 CSoutput.n51 gnd 0.040352f
C5260 CSoutput.n52 gnd 0.048358f
C5261 CSoutput.n53 gnd 0.048358f
C5262 CSoutput.n54 gnd 0.03934f
C5263 CSoutput.n55 gnd 0.037894f
C5264 CSoutput.n56 gnd 0.142867f
C5265 CSoutput.n57 gnd 0.039623f
C5266 CSoutput.n58 gnd 0.048358f
C5267 CSoutput.n59 gnd 0.048358f
C5268 CSoutput.n60 gnd 0.048358f
C5269 CSoutput.n61 gnd 0.034472f
C5270 CSoutput.n62 gnd 0.146047f
C5271 CSoutput.n63 gnd 0.034003f
C5272 CSoutput.t169 gnd 0.319878f
C5273 CSoutput.n64 gnd 0.142867f
C5274 CSoutput.n65 gnd 0.04005f
C5275 CSoutput.n66 gnd 0.048358f
C5276 CSoutput.n67 gnd 0.048358f
C5277 CSoutput.n68 gnd 0.048358f
C5278 CSoutput.n69 gnd 0.038906f
C5279 CSoutput.n70 gnd 0.142867f
C5280 CSoutput.n71 gnd 0.04036f
C5281 CSoutput.n72 gnd 0.035299f
C5282 CSoutput.n73 gnd 0.048358f
C5283 CSoutput.n74 gnd 0.048358f
C5284 CSoutput.n75 gnd 0.036608f
C5285 CSoutput.n76 gnd 0.021742f
C5286 CSoutput.t179 gnd 0.359406f
C5287 CSoutput.n77 gnd 0.178538f
C5288 CSoutput.n78 gnd 0.763844f
C5289 CSoutput.t30 gnd 0.06032f
C5290 CSoutput.t17 gnd 0.06032f
C5291 CSoutput.n79 gnd 0.467016f
C5292 CSoutput.t83 gnd 0.06032f
C5293 CSoutput.t153 gnd 0.06032f
C5294 CSoutput.n80 gnd 0.466184f
C5295 CSoutput.n81 gnd 0.473176f
C5296 CSoutput.t15 gnd 0.06032f
C5297 CSoutput.t90 gnd 0.06032f
C5298 CSoutput.n82 gnd 0.466184f
C5299 CSoutput.n83 gnd 0.233161f
C5300 CSoutput.t45 gnd 0.06032f
C5301 CSoutput.t64 gnd 0.06032f
C5302 CSoutput.n84 gnd 0.466184f
C5303 CSoutput.n85 gnd 0.233161f
C5304 CSoutput.t46 gnd 0.06032f
C5305 CSoutput.t77 gnd 0.06032f
C5306 CSoutput.n86 gnd 0.466184f
C5307 CSoutput.n87 gnd 0.233161f
C5308 CSoutput.t61 gnd 0.06032f
C5309 CSoutput.t35 gnd 0.06032f
C5310 CSoutput.n88 gnd 0.466184f
C5311 CSoutput.n89 gnd 0.233161f
C5312 CSoutput.t165 gnd 0.06032f
C5313 CSoutput.t97 gnd 0.06032f
C5314 CSoutput.n90 gnd 0.466184f
C5315 CSoutput.n91 gnd 0.233161f
C5316 CSoutput.t2 gnd 0.06032f
C5317 CSoutput.t89 gnd 0.06032f
C5318 CSoutput.n92 gnd 0.466184f
C5319 CSoutput.n93 gnd 0.233161f
C5320 CSoutput.t44 gnd 0.06032f
C5321 CSoutput.t37 gnd 0.06032f
C5322 CSoutput.n94 gnd 0.466184f
C5323 CSoutput.n95 gnd 0.233161f
C5324 CSoutput.t93 gnd 0.06032f
C5325 CSoutput.t76 gnd 0.06032f
C5326 CSoutput.n96 gnd 0.466184f
C5327 CSoutput.n97 gnd 0.427564f
C5328 CSoutput.t57 gnd 0.06032f
C5329 CSoutput.t43 gnd 0.06032f
C5330 CSoutput.n98 gnd 0.467016f
C5331 CSoutput.t50 gnd 0.06032f
C5332 CSoutput.t65 gnd 0.06032f
C5333 CSoutput.n99 gnd 0.466184f
C5334 CSoutput.n100 gnd 0.473176f
C5335 CSoutput.t25 gnd 0.06032f
C5336 CSoutput.t78 gnd 0.06032f
C5337 CSoutput.n101 gnd 0.466184f
C5338 CSoutput.n102 gnd 0.233161f
C5339 CSoutput.t51 gnd 0.06032f
C5340 CSoutput.t41 gnd 0.06032f
C5341 CSoutput.n103 gnd 0.466184f
C5342 CSoutput.n104 gnd 0.233161f
C5343 CSoutput.t33 gnd 0.06032f
C5344 CSoutput.t81 gnd 0.06032f
C5345 CSoutput.n105 gnd 0.466184f
C5346 CSoutput.n106 gnd 0.233161f
C5347 CSoutput.t161 gnd 0.06032f
C5348 CSoutput.t67 gnd 0.06032f
C5349 CSoutput.n107 gnd 0.466184f
C5350 CSoutput.n108 gnd 0.233161f
C5351 CSoutput.t74 gnd 0.06032f
C5352 CSoutput.t18 gnd 0.06032f
C5353 CSoutput.n109 gnd 0.466184f
C5354 CSoutput.n110 gnd 0.233161f
C5355 CSoutput.t56 gnd 0.06032f
C5356 CSoutput.t42 gnd 0.06032f
C5357 CSoutput.n111 gnd 0.466184f
C5358 CSoutput.n112 gnd 0.233161f
C5359 CSoutput.t156 gnd 0.06032f
C5360 CSoutput.t96 gnd 0.06032f
C5361 CSoutput.n113 gnd 0.466184f
C5362 CSoutput.n114 gnd 0.233161f
C5363 CSoutput.t24 gnd 0.06032f
C5364 CSoutput.t16 gnd 0.06032f
C5365 CSoutput.n115 gnd 0.466184f
C5366 CSoutput.n116 gnd 0.347702f
C5367 CSoutput.n117 gnd 0.43845f
C5368 CSoutput.t10 gnd 0.06032f
C5369 CSoutput.t80 gnd 0.06032f
C5370 CSoutput.n118 gnd 0.467016f
C5371 CSoutput.t166 gnd 0.06032f
C5372 CSoutput.t158 gnd 0.06032f
C5373 CSoutput.n119 gnd 0.466184f
C5374 CSoutput.n120 gnd 0.473176f
C5375 CSoutput.t84 gnd 0.06032f
C5376 CSoutput.t22 gnd 0.06032f
C5377 CSoutput.n121 gnd 0.466184f
C5378 CSoutput.n122 gnd 0.233161f
C5379 CSoutput.t167 gnd 0.06032f
C5380 CSoutput.t82 gnd 0.06032f
C5381 CSoutput.n123 gnd 0.466184f
C5382 CSoutput.n124 gnd 0.233161f
C5383 CSoutput.t92 gnd 0.06032f
C5384 CSoutput.t164 gnd 0.06032f
C5385 CSoutput.n125 gnd 0.466184f
C5386 CSoutput.n126 gnd 0.233161f
C5387 CSoutput.t54 gnd 0.06032f
C5388 CSoutput.t69 gnd 0.06032f
C5389 CSoutput.n127 gnd 0.466184f
C5390 CSoutput.n128 gnd 0.233161f
C5391 CSoutput.t88 gnd 0.06032f
C5392 CSoutput.t72 gnd 0.06032f
C5393 CSoutput.n129 gnd 0.466184f
C5394 CSoutput.n130 gnd 0.233161f
C5395 CSoutput.t159 gnd 0.06032f
C5396 CSoutput.t163 gnd 0.06032f
C5397 CSoutput.n131 gnd 0.466184f
C5398 CSoutput.n132 gnd 0.233161f
C5399 CSoutput.t23 gnd 0.06032f
C5400 CSoutput.t86 gnd 0.06032f
C5401 CSoutput.n133 gnd 0.466184f
C5402 CSoutput.n134 gnd 0.233161f
C5403 CSoutput.t11 gnd 0.06032f
C5404 CSoutput.t85 gnd 0.06032f
C5405 CSoutput.n135 gnd 0.466184f
C5406 CSoutput.n136 gnd 0.347702f
C5407 CSoutput.n137 gnd 0.490075f
C5408 CSoutput.n138 gnd 9.38805f
C5409 CSoutput.n140 gnd 0.855445f
C5410 CSoutput.n141 gnd 0.641584f
C5411 CSoutput.n142 gnd 0.855445f
C5412 CSoutput.n143 gnd 0.855445f
C5413 CSoutput.n144 gnd 2.30312f
C5414 CSoutput.n145 gnd 0.855445f
C5415 CSoutput.n146 gnd 0.855445f
C5416 CSoutput.t185 gnd 1.06931f
C5417 CSoutput.n147 gnd 0.855445f
C5418 CSoutput.n148 gnd 0.855445f
C5419 CSoutput.n152 gnd 0.855445f
C5420 CSoutput.n156 gnd 0.855445f
C5421 CSoutput.n157 gnd 0.855445f
C5422 CSoutput.n159 gnd 0.855445f
C5423 CSoutput.n164 gnd 0.855445f
C5424 CSoutput.n166 gnd 0.855445f
C5425 CSoutput.n167 gnd 0.855445f
C5426 CSoutput.n169 gnd 0.855445f
C5427 CSoutput.n170 gnd 0.855445f
C5428 CSoutput.n172 gnd 0.855445f
C5429 CSoutput.t170 gnd 14.294401f
C5430 CSoutput.n174 gnd 0.855445f
C5431 CSoutput.n175 gnd 0.641584f
C5432 CSoutput.n176 gnd 0.855445f
C5433 CSoutput.n177 gnd 0.855445f
C5434 CSoutput.n178 gnd 2.30312f
C5435 CSoutput.n179 gnd 0.855445f
C5436 CSoutput.n180 gnd 0.855445f
C5437 CSoutput.t171 gnd 1.06931f
C5438 CSoutput.n181 gnd 0.855445f
C5439 CSoutput.n182 gnd 0.855445f
C5440 CSoutput.n186 gnd 0.855445f
C5441 CSoutput.n190 gnd 0.855445f
C5442 CSoutput.n191 gnd 0.855445f
C5443 CSoutput.n193 gnd 0.855445f
C5444 CSoutput.n198 gnd 0.855445f
C5445 CSoutput.n200 gnd 0.855445f
C5446 CSoutput.n201 gnd 0.855445f
C5447 CSoutput.n203 gnd 0.855445f
C5448 CSoutput.n204 gnd 0.855445f
C5449 CSoutput.n206 gnd 0.855445f
C5450 CSoutput.n207 gnd 0.641584f
C5451 CSoutput.n209 gnd 0.855445f
C5452 CSoutput.n210 gnd 0.641584f
C5453 CSoutput.n211 gnd 0.855445f
C5454 CSoutput.n212 gnd 0.855445f
C5455 CSoutput.n213 gnd 2.30312f
C5456 CSoutput.n214 gnd 0.855445f
C5457 CSoutput.n215 gnd 0.855445f
C5458 CSoutput.t178 gnd 1.06931f
C5459 CSoutput.n216 gnd 0.855445f
C5460 CSoutput.n217 gnd 2.30312f
C5461 CSoutput.n219 gnd 0.855445f
C5462 CSoutput.n220 gnd 0.855445f
C5463 CSoutput.n222 gnd 0.855445f
C5464 CSoutput.n223 gnd 0.855445f
C5465 CSoutput.t189 gnd 14.0614f
C5466 CSoutput.t177 gnd 14.294401f
C5467 CSoutput.n229 gnd 2.68366f
C5468 CSoutput.n230 gnd 10.9322f
C5469 CSoutput.n231 gnd 11.389701f
C5470 CSoutput.n236 gnd 2.90712f
C5471 CSoutput.n242 gnd 0.855445f
C5472 CSoutput.n244 gnd 0.855445f
C5473 CSoutput.n246 gnd 0.855445f
C5474 CSoutput.n248 gnd 0.855445f
C5475 CSoutput.n250 gnd 0.855445f
C5476 CSoutput.n256 gnd 0.855445f
C5477 CSoutput.n263 gnd 1.56941f
C5478 CSoutput.n264 gnd 1.56941f
C5479 CSoutput.n265 gnd 0.855445f
C5480 CSoutput.n266 gnd 0.855445f
C5481 CSoutput.n268 gnd 0.641584f
C5482 CSoutput.n269 gnd 0.549459f
C5483 CSoutput.n271 gnd 0.641584f
C5484 CSoutput.n272 gnd 0.549459f
C5485 CSoutput.n273 gnd 0.641584f
C5486 CSoutput.n275 gnd 0.855445f
C5487 CSoutput.n277 gnd 2.30312f
C5488 CSoutput.n278 gnd 2.68366f
C5489 CSoutput.n279 gnd 10.0549f
C5490 CSoutput.n281 gnd 0.641584f
C5491 CSoutput.n282 gnd 1.65083f
C5492 CSoutput.n283 gnd 0.641584f
C5493 CSoutput.n285 gnd 0.855445f
C5494 CSoutput.n287 gnd 2.30312f
C5495 CSoutput.n288 gnd 5.01604f
C5496 CSoutput.t8 gnd 0.06032f
C5497 CSoutput.t6 gnd 0.06032f
C5498 CSoutput.n289 gnd 0.467016f
C5499 CSoutput.t154 gnd 0.06032f
C5500 CSoutput.t68 gnd 0.06032f
C5501 CSoutput.n290 gnd 0.466184f
C5502 CSoutput.n291 gnd 0.473176f
C5503 CSoutput.t91 gnd 0.06032f
C5504 CSoutput.t4 gnd 0.06032f
C5505 CSoutput.n292 gnd 0.466184f
C5506 CSoutput.n293 gnd 0.233161f
C5507 CSoutput.t94 gnd 0.06032f
C5508 CSoutput.t162 gnd 0.06032f
C5509 CSoutput.n294 gnd 0.466184f
C5510 CSoutput.n295 gnd 0.233161f
C5511 CSoutput.t99 gnd 0.06032f
C5512 CSoutput.t47 gnd 0.06032f
C5513 CSoutput.n296 gnd 0.466184f
C5514 CSoutput.n297 gnd 0.233161f
C5515 CSoutput.t70 gnd 0.06032f
C5516 CSoutput.t60 gnd 0.06032f
C5517 CSoutput.n298 gnd 0.466184f
C5518 CSoutput.n299 gnd 0.233161f
C5519 CSoutput.t152 gnd 0.06032f
C5520 CSoutput.t62 gnd 0.06032f
C5521 CSoutput.n300 gnd 0.466184f
C5522 CSoutput.n301 gnd 0.233161f
C5523 CSoutput.t102 gnd 0.06032f
C5524 CSoutput.t3 gnd 0.06032f
C5525 CSoutput.n302 gnd 0.466184f
C5526 CSoutput.n303 gnd 0.233161f
C5527 CSoutput.t66 gnd 0.06032f
C5528 CSoutput.t0 gnd 0.06032f
C5529 CSoutput.n304 gnd 0.466184f
C5530 CSoutput.n305 gnd 0.233161f
C5531 CSoutput.t98 gnd 0.06032f
C5532 CSoutput.t73 gnd 0.06032f
C5533 CSoutput.n306 gnd 0.466184f
C5534 CSoutput.n307 gnd 0.427564f
C5535 CSoutput.t38 gnd 0.06032f
C5536 CSoutput.t75 gnd 0.06032f
C5537 CSoutput.n308 gnd 0.467016f
C5538 CSoutput.t26 gnd 0.06032f
C5539 CSoutput.t34 gnd 0.06032f
C5540 CSoutput.n309 gnd 0.466184f
C5541 CSoutput.n310 gnd 0.473176f
C5542 CSoutput.t155 gnd 0.06032f
C5543 CSoutput.t13 gnd 0.06032f
C5544 CSoutput.n311 gnd 0.466184f
C5545 CSoutput.n312 gnd 0.233161f
C5546 CSoutput.t9 gnd 0.06032f
C5547 CSoutput.t71 gnd 0.06032f
C5548 CSoutput.n313 gnd 0.466184f
C5549 CSoutput.n314 gnd 0.233161f
C5550 CSoutput.t87 gnd 0.06032f
C5551 CSoutput.t160 gnd 0.06032f
C5552 CSoutput.n315 gnd 0.466184f
C5553 CSoutput.n316 gnd 0.233161f
C5554 CSoutput.t32 gnd 0.06032f
C5555 CSoutput.t31 gnd 0.06032f
C5556 CSoutput.n317 gnd 0.466184f
C5557 CSoutput.n318 gnd 0.233161f
C5558 CSoutput.t7 gnd 0.06032f
C5559 CSoutput.t49 gnd 0.06032f
C5560 CSoutput.n319 gnd 0.466184f
C5561 CSoutput.n320 gnd 0.233161f
C5562 CSoutput.t39 gnd 0.06032f
C5563 CSoutput.t27 gnd 0.06032f
C5564 CSoutput.n321 gnd 0.466184f
C5565 CSoutput.n322 gnd 0.233161f
C5566 CSoutput.t52 gnd 0.06032f
C5567 CSoutput.t20 gnd 0.06032f
C5568 CSoutput.n323 gnd 0.466184f
C5569 CSoutput.n324 gnd 0.233161f
C5570 CSoutput.t59 gnd 0.06032f
C5571 CSoutput.t58 gnd 0.06032f
C5572 CSoutput.n325 gnd 0.466184f
C5573 CSoutput.n326 gnd 0.347702f
C5574 CSoutput.n327 gnd 0.43845f
C5575 CSoutput.t28 gnd 0.06032f
C5576 CSoutput.t103 gnd 0.06032f
C5577 CSoutput.n328 gnd 0.467016f
C5578 CSoutput.t53 gnd 0.06032f
C5579 CSoutput.t21 gnd 0.06032f
C5580 CSoutput.n329 gnd 0.466184f
C5581 CSoutput.n330 gnd 0.473176f
C5582 CSoutput.t100 gnd 0.06032f
C5583 CSoutput.t5 gnd 0.06032f
C5584 CSoutput.n331 gnd 0.466184f
C5585 CSoutput.n332 gnd 0.233161f
C5586 CSoutput.t48 gnd 0.06032f
C5587 CSoutput.t36 gnd 0.06032f
C5588 CSoutput.n333 gnd 0.466184f
C5589 CSoutput.n334 gnd 0.233161f
C5590 CSoutput.t40 gnd 0.06032f
C5591 CSoutput.t63 gnd 0.06032f
C5592 CSoutput.n335 gnd 0.466184f
C5593 CSoutput.n336 gnd 0.233161f
C5594 CSoutput.t95 gnd 0.06032f
C5595 CSoutput.t12 gnd 0.06032f
C5596 CSoutput.n337 gnd 0.466184f
C5597 CSoutput.n338 gnd 0.233161f
C5598 CSoutput.t55 gnd 0.06032f
C5599 CSoutput.t19 gnd 0.06032f
C5600 CSoutput.n339 gnd 0.466184f
C5601 CSoutput.n340 gnd 0.233161f
C5602 CSoutput.t29 gnd 0.06032f
C5603 CSoutput.t14 gnd 0.06032f
C5604 CSoutput.n341 gnd 0.466184f
C5605 CSoutput.n342 gnd 0.233161f
C5606 CSoutput.t1 gnd 0.06032f
C5607 CSoutput.t101 gnd 0.06032f
C5608 CSoutput.n343 gnd 0.466184f
C5609 CSoutput.n344 gnd 0.233161f
C5610 CSoutput.t157 gnd 0.06032f
C5611 CSoutput.t79 gnd 0.06032f
C5612 CSoutput.n345 gnd 0.466182f
C5613 CSoutput.n346 gnd 0.347703f
C5614 CSoutput.n347 gnd 0.490075f
C5615 CSoutput.n348 gnd 13.494201f
C5616 CSoutput.t142 gnd 0.05278f
C5617 CSoutput.t134 gnd 0.05278f
C5618 CSoutput.n349 gnd 0.467942f
C5619 CSoutput.t105 gnd 0.05278f
C5620 CSoutput.t107 gnd 0.05278f
C5621 CSoutput.n350 gnd 0.466381f
C5622 CSoutput.n351 gnd 0.43458f
C5623 CSoutput.t122 gnd 0.05278f
C5624 CSoutput.t128 gnd 0.05278f
C5625 CSoutput.n352 gnd 0.466381f
C5626 CSoutput.n353 gnd 0.214228f
C5627 CSoutput.t110 gnd 0.05278f
C5628 CSoutput.t143 gnd 0.05278f
C5629 CSoutput.n354 gnd 0.466381f
C5630 CSoutput.n355 gnd 0.214228f
C5631 CSoutput.t146 gnd 0.05278f
C5632 CSoutput.t120 gnd 0.05278f
C5633 CSoutput.n356 gnd 0.466381f
C5634 CSoutput.n357 gnd 0.214228f
C5635 CSoutput.t148 gnd 0.05278f
C5636 CSoutput.t113 gnd 0.05278f
C5637 CSoutput.n358 gnd 0.466381f
C5638 CSoutput.n359 gnd 0.395079f
C5639 CSoutput.t112 gnd 0.05278f
C5640 CSoutput.t126 gnd 0.05278f
C5641 CSoutput.n360 gnd 0.467942f
C5642 CSoutput.t150 gnd 0.05278f
C5643 CSoutput.t140 gnd 0.05278f
C5644 CSoutput.n361 gnd 0.466381f
C5645 CSoutput.n362 gnd 0.43458f
C5646 CSoutput.t147 gnd 0.05278f
C5647 CSoutput.t121 gnd 0.05278f
C5648 CSoutput.n363 gnd 0.466381f
C5649 CSoutput.n364 gnd 0.214228f
C5650 CSoutput.t137 gnd 0.05278f
C5651 CSoutput.t114 gnd 0.05278f
C5652 CSoutput.n365 gnd 0.466381f
C5653 CSoutput.n366 gnd 0.214228f
C5654 CSoutput.t117 gnd 0.05278f
C5655 CSoutput.t145 gnd 0.05278f
C5656 CSoutput.n367 gnd 0.466381f
C5657 CSoutput.n368 gnd 0.214228f
C5658 CSoutput.t116 gnd 0.05278f
C5659 CSoutput.t106 gnd 0.05278f
C5660 CSoutput.n369 gnd 0.466381f
C5661 CSoutput.n370 gnd 0.325243f
C5662 CSoutput.n371 gnd 0.604327f
C5663 CSoutput.n372 gnd 13.190599f
C5664 CSoutput.t136 gnd 0.05278f
C5665 CSoutput.t131 gnd 0.05278f
C5666 CSoutput.n373 gnd 0.467942f
C5667 CSoutput.t111 gnd 0.05278f
C5668 CSoutput.t109 gnd 0.05278f
C5669 CSoutput.n374 gnd 0.466381f
C5670 CSoutput.n375 gnd 0.43458f
C5671 CSoutput.t151 gnd 0.05278f
C5672 CSoutput.t127 gnd 0.05278f
C5673 CSoutput.n376 gnd 0.466381f
C5674 CSoutput.n377 gnd 0.214228f
C5675 CSoutput.t132 gnd 0.05278f
C5676 CSoutput.t141 gnd 0.05278f
C5677 CSoutput.n378 gnd 0.466381f
C5678 CSoutput.n379 gnd 0.214228f
C5679 CSoutput.t138 gnd 0.05278f
C5680 CSoutput.t118 gnd 0.05278f
C5681 CSoutput.n380 gnd 0.466381f
C5682 CSoutput.n381 gnd 0.214228f
C5683 CSoutput.t123 gnd 0.05278f
C5684 CSoutput.t115 gnd 0.05278f
C5685 CSoutput.n382 gnd 0.466381f
C5686 CSoutput.n383 gnd 0.395079f
C5687 CSoutput.t130 gnd 0.05278f
C5688 CSoutput.t124 gnd 0.05278f
C5689 CSoutput.n384 gnd 0.467942f
C5690 CSoutput.t104 gnd 0.05278f
C5691 CSoutput.t135 gnd 0.05278f
C5692 CSoutput.n385 gnd 0.466381f
C5693 CSoutput.n386 gnd 0.43458f
C5694 CSoutput.t139 gnd 0.05278f
C5695 CSoutput.t119 gnd 0.05278f
C5696 CSoutput.n387 gnd 0.466381f
C5697 CSoutput.n388 gnd 0.214228f
C5698 CSoutput.t125 gnd 0.05278f
C5699 CSoutput.t129 gnd 0.05278f
C5700 CSoutput.n389 gnd 0.466381f
C5701 CSoutput.n390 gnd 0.214228f
C5702 CSoutput.t133 gnd 0.05278f
C5703 CSoutput.t144 gnd 0.05278f
C5704 CSoutput.n391 gnd 0.466381f
C5705 CSoutput.n392 gnd 0.214228f
C5706 CSoutput.t149 gnd 0.05278f
C5707 CSoutput.t108 gnd 0.05278f
C5708 CSoutput.n393 gnd 0.466381f
C5709 CSoutput.n394 gnd 0.325243f
C5710 CSoutput.n395 gnd 0.604327f
C5711 CSoutput.n396 gnd 7.8742f
C5712 CSoutput.n397 gnd 15.4615f
C5713 commonsourceibias.n0 gnd 0.010306f
C5714 commonsourceibias.t71 gnd 0.156059f
C5715 commonsourceibias.t81 gnd 0.144299f
C5716 commonsourceibias.n1 gnd 0.057575f
C5717 commonsourceibias.n2 gnd 0.007723f
C5718 commonsourceibias.t55 gnd 0.144299f
C5719 commonsourceibias.n3 gnd 0.006248f
C5720 commonsourceibias.n4 gnd 0.007723f
C5721 commonsourceibias.t53 gnd 0.144299f
C5722 commonsourceibias.n5 gnd 0.007456f
C5723 commonsourceibias.n6 gnd 0.007723f
C5724 commonsourceibias.t76 gnd 0.144299f
C5725 commonsourceibias.n7 gnd 0.057575f
C5726 commonsourceibias.t87 gnd 0.144299f
C5727 commonsourceibias.n8 gnd 0.006238f
C5728 commonsourceibias.n9 gnd 0.010306f
C5729 commonsourceibias.t16 gnd 0.156059f
C5730 commonsourceibias.t32 gnd 0.144299f
C5731 commonsourceibias.n10 gnd 0.057575f
C5732 commonsourceibias.n11 gnd 0.007723f
C5733 commonsourceibias.t44 gnd 0.144299f
C5734 commonsourceibias.n12 gnd 0.006248f
C5735 commonsourceibias.n13 gnd 0.007723f
C5736 commonsourceibias.t14 gnd 0.144299f
C5737 commonsourceibias.n14 gnd 0.007456f
C5738 commonsourceibias.n15 gnd 0.007723f
C5739 commonsourceibias.t22 gnd 0.144299f
C5740 commonsourceibias.n16 gnd 0.057575f
C5741 commonsourceibias.t0 gnd 0.144299f
C5742 commonsourceibias.n17 gnd 0.006238f
C5743 commonsourceibias.n18 gnd 0.007723f
C5744 commonsourceibias.t8 gnd 0.144299f
C5745 commonsourceibias.t10 gnd 0.144299f
C5746 commonsourceibias.n19 gnd 0.057575f
C5747 commonsourceibias.n20 gnd 0.007723f
C5748 commonsourceibias.t18 gnd 0.144299f
C5749 commonsourceibias.n21 gnd 0.057575f
C5750 commonsourceibias.n22 gnd 0.007723f
C5751 commonsourceibias.t28 gnd 0.144299f
C5752 commonsourceibias.n23 gnd 0.057575f
C5753 commonsourceibias.n24 gnd 0.038882f
C5754 commonsourceibias.t4 gnd 0.144299f
C5755 commonsourceibias.t46 gnd 0.162824f
C5756 commonsourceibias.n25 gnd 0.066816f
C5757 commonsourceibias.n26 gnd 0.069172f
C5758 commonsourceibias.n27 gnd 0.009519f
C5759 commonsourceibias.n28 gnd 0.010531f
C5760 commonsourceibias.n29 gnd 0.007723f
C5761 commonsourceibias.n30 gnd 0.007723f
C5762 commonsourceibias.n31 gnd 0.010462f
C5763 commonsourceibias.n32 gnd 0.006248f
C5764 commonsourceibias.n33 gnd 0.010592f
C5765 commonsourceibias.n34 gnd 0.007723f
C5766 commonsourceibias.n35 gnd 0.007723f
C5767 commonsourceibias.n36 gnd 0.010657f
C5768 commonsourceibias.n37 gnd 0.009189f
C5769 commonsourceibias.n38 gnd 0.007456f
C5770 commonsourceibias.n39 gnd 0.007723f
C5771 commonsourceibias.n40 gnd 0.007723f
C5772 commonsourceibias.n41 gnd 0.009447f
C5773 commonsourceibias.n42 gnd 0.010603f
C5774 commonsourceibias.n43 gnd 0.057575f
C5775 commonsourceibias.n44 gnd 0.010532f
C5776 commonsourceibias.n45 gnd 0.007723f
C5777 commonsourceibias.n46 gnd 0.007723f
C5778 commonsourceibias.n47 gnd 0.007723f
C5779 commonsourceibias.n48 gnd 0.010532f
C5780 commonsourceibias.n49 gnd 0.057575f
C5781 commonsourceibias.n50 gnd 0.010603f
C5782 commonsourceibias.n51 gnd 0.009447f
C5783 commonsourceibias.n52 gnd 0.007723f
C5784 commonsourceibias.n53 gnd 0.007723f
C5785 commonsourceibias.n54 gnd 0.007723f
C5786 commonsourceibias.n55 gnd 0.009189f
C5787 commonsourceibias.n56 gnd 0.010657f
C5788 commonsourceibias.n57 gnd 0.057575f
C5789 commonsourceibias.n58 gnd 0.010592f
C5790 commonsourceibias.n59 gnd 0.007723f
C5791 commonsourceibias.n60 gnd 0.007723f
C5792 commonsourceibias.n61 gnd 0.007723f
C5793 commonsourceibias.n62 gnd 0.010462f
C5794 commonsourceibias.n63 gnd 0.057575f
C5795 commonsourceibias.n64 gnd 0.010531f
C5796 commonsourceibias.n65 gnd 0.009519f
C5797 commonsourceibias.n66 gnd 0.007723f
C5798 commonsourceibias.n67 gnd 0.007723f
C5799 commonsourceibias.n68 gnd 0.007835f
C5800 commonsourceibias.n69 gnd 0.0081f
C5801 commonsourceibias.n70 gnd 0.068889f
C5802 commonsourceibias.n71 gnd 0.076422f
C5803 commonsourceibias.t17 gnd 0.016666f
C5804 commonsourceibias.t33 gnd 0.016666f
C5805 commonsourceibias.n72 gnd 0.147271f
C5806 commonsourceibias.n73 gnd 0.127253f
C5807 commonsourceibias.t45 gnd 0.016666f
C5808 commonsourceibias.t15 gnd 0.016666f
C5809 commonsourceibias.n74 gnd 0.147271f
C5810 commonsourceibias.n75 gnd 0.067647f
C5811 commonsourceibias.t23 gnd 0.016666f
C5812 commonsourceibias.t1 gnd 0.016666f
C5813 commonsourceibias.n76 gnd 0.147271f
C5814 commonsourceibias.n77 gnd 0.056516f
C5815 commonsourceibias.t5 gnd 0.016666f
C5816 commonsourceibias.t47 gnd 0.016666f
C5817 commonsourceibias.n78 gnd 0.147764f
C5818 commonsourceibias.t19 gnd 0.016666f
C5819 commonsourceibias.t29 gnd 0.016666f
C5820 commonsourceibias.n79 gnd 0.147271f
C5821 commonsourceibias.n80 gnd 0.137229f
C5822 commonsourceibias.t9 gnd 0.016666f
C5823 commonsourceibias.t11 gnd 0.016666f
C5824 commonsourceibias.n81 gnd 0.147271f
C5825 commonsourceibias.n82 gnd 0.056516f
C5826 commonsourceibias.n83 gnd 0.068435f
C5827 commonsourceibias.n84 gnd 0.007723f
C5828 commonsourceibias.t50 gnd 0.144299f
C5829 commonsourceibias.t70 gnd 0.144299f
C5830 commonsourceibias.n85 gnd 0.057575f
C5831 commonsourceibias.n86 gnd 0.007723f
C5832 commonsourceibias.t67 gnd 0.144299f
C5833 commonsourceibias.n87 gnd 0.057575f
C5834 commonsourceibias.n88 gnd 0.007723f
C5835 commonsourceibias.t78 gnd 0.144299f
C5836 commonsourceibias.n89 gnd 0.057575f
C5837 commonsourceibias.n90 gnd 0.038882f
C5838 commonsourceibias.t65 gnd 0.144299f
C5839 commonsourceibias.t62 gnd 0.162824f
C5840 commonsourceibias.n91 gnd 0.066816f
C5841 commonsourceibias.n92 gnd 0.069172f
C5842 commonsourceibias.n93 gnd 0.009519f
C5843 commonsourceibias.n94 gnd 0.010531f
C5844 commonsourceibias.n95 gnd 0.007723f
C5845 commonsourceibias.n96 gnd 0.007723f
C5846 commonsourceibias.n97 gnd 0.010462f
C5847 commonsourceibias.n98 gnd 0.006248f
C5848 commonsourceibias.n99 gnd 0.010592f
C5849 commonsourceibias.n100 gnd 0.007723f
C5850 commonsourceibias.n101 gnd 0.007723f
C5851 commonsourceibias.n102 gnd 0.010657f
C5852 commonsourceibias.n103 gnd 0.009189f
C5853 commonsourceibias.n104 gnd 0.007456f
C5854 commonsourceibias.n105 gnd 0.007723f
C5855 commonsourceibias.n106 gnd 0.007723f
C5856 commonsourceibias.n107 gnd 0.009447f
C5857 commonsourceibias.n108 gnd 0.010603f
C5858 commonsourceibias.n109 gnd 0.057575f
C5859 commonsourceibias.n110 gnd 0.010532f
C5860 commonsourceibias.n111 gnd 0.007686f
C5861 commonsourceibias.n112 gnd 0.055832f
C5862 commonsourceibias.n113 gnd 0.007686f
C5863 commonsourceibias.n114 gnd 0.010532f
C5864 commonsourceibias.n115 gnd 0.057575f
C5865 commonsourceibias.n116 gnd 0.010603f
C5866 commonsourceibias.n117 gnd 0.009447f
C5867 commonsourceibias.n118 gnd 0.007723f
C5868 commonsourceibias.n119 gnd 0.007723f
C5869 commonsourceibias.n120 gnd 0.007723f
C5870 commonsourceibias.n121 gnd 0.009189f
C5871 commonsourceibias.n122 gnd 0.010657f
C5872 commonsourceibias.n123 gnd 0.057575f
C5873 commonsourceibias.n124 gnd 0.010592f
C5874 commonsourceibias.n125 gnd 0.007723f
C5875 commonsourceibias.n126 gnd 0.007723f
C5876 commonsourceibias.n127 gnd 0.007723f
C5877 commonsourceibias.n128 gnd 0.010462f
C5878 commonsourceibias.n129 gnd 0.057575f
C5879 commonsourceibias.n130 gnd 0.010531f
C5880 commonsourceibias.n131 gnd 0.009519f
C5881 commonsourceibias.n132 gnd 0.007723f
C5882 commonsourceibias.n133 gnd 0.007723f
C5883 commonsourceibias.n134 gnd 0.007835f
C5884 commonsourceibias.n135 gnd 0.0081f
C5885 commonsourceibias.n136 gnd 0.068889f
C5886 commonsourceibias.n137 gnd 0.044582f
C5887 commonsourceibias.n138 gnd 0.010306f
C5888 commonsourceibias.t72 gnd 0.144299f
C5889 commonsourceibias.n139 gnd 0.057575f
C5890 commonsourceibias.n140 gnd 0.007723f
C5891 commonsourceibias.t49 gnd 0.144299f
C5892 commonsourceibias.n141 gnd 0.006248f
C5893 commonsourceibias.n142 gnd 0.007723f
C5894 commonsourceibias.t95 gnd 0.144299f
C5895 commonsourceibias.n143 gnd 0.007456f
C5896 commonsourceibias.n144 gnd 0.007723f
C5897 commonsourceibias.t66 gnd 0.144299f
C5898 commonsourceibias.n145 gnd 0.057575f
C5899 commonsourceibias.t77 gnd 0.144299f
C5900 commonsourceibias.n146 gnd 0.006238f
C5901 commonsourceibias.n147 gnd 0.007723f
C5902 commonsourceibias.t91 gnd 0.144299f
C5903 commonsourceibias.t60 gnd 0.144299f
C5904 commonsourceibias.n148 gnd 0.057575f
C5905 commonsourceibias.n149 gnd 0.007723f
C5906 commonsourceibias.t58 gnd 0.144299f
C5907 commonsourceibias.n150 gnd 0.057575f
C5908 commonsourceibias.n151 gnd 0.007723f
C5909 commonsourceibias.t68 gnd 0.144299f
C5910 commonsourceibias.n152 gnd 0.057575f
C5911 commonsourceibias.n153 gnd 0.038882f
C5912 commonsourceibias.t57 gnd 0.144299f
C5913 commonsourceibias.t54 gnd 0.162824f
C5914 commonsourceibias.n154 gnd 0.066816f
C5915 commonsourceibias.n155 gnd 0.069172f
C5916 commonsourceibias.n156 gnd 0.009519f
C5917 commonsourceibias.n157 gnd 0.010531f
C5918 commonsourceibias.n158 gnd 0.007723f
C5919 commonsourceibias.n159 gnd 0.007723f
C5920 commonsourceibias.n160 gnd 0.010462f
C5921 commonsourceibias.n161 gnd 0.006248f
C5922 commonsourceibias.n162 gnd 0.010592f
C5923 commonsourceibias.n163 gnd 0.007723f
C5924 commonsourceibias.n164 gnd 0.007723f
C5925 commonsourceibias.n165 gnd 0.010657f
C5926 commonsourceibias.n166 gnd 0.009189f
C5927 commonsourceibias.n167 gnd 0.007456f
C5928 commonsourceibias.n168 gnd 0.007723f
C5929 commonsourceibias.n169 gnd 0.007723f
C5930 commonsourceibias.n170 gnd 0.009447f
C5931 commonsourceibias.n171 gnd 0.010603f
C5932 commonsourceibias.n172 gnd 0.057575f
C5933 commonsourceibias.n173 gnd 0.010532f
C5934 commonsourceibias.n174 gnd 0.007723f
C5935 commonsourceibias.n175 gnd 0.007723f
C5936 commonsourceibias.n176 gnd 0.007723f
C5937 commonsourceibias.n177 gnd 0.010532f
C5938 commonsourceibias.n178 gnd 0.057575f
C5939 commonsourceibias.n179 gnd 0.010603f
C5940 commonsourceibias.n180 gnd 0.009447f
C5941 commonsourceibias.n181 gnd 0.007723f
C5942 commonsourceibias.n182 gnd 0.007723f
C5943 commonsourceibias.n183 gnd 0.007723f
C5944 commonsourceibias.n184 gnd 0.009189f
C5945 commonsourceibias.n185 gnd 0.010657f
C5946 commonsourceibias.n186 gnd 0.057575f
C5947 commonsourceibias.n187 gnd 0.010592f
C5948 commonsourceibias.n188 gnd 0.007723f
C5949 commonsourceibias.n189 gnd 0.007723f
C5950 commonsourceibias.n190 gnd 0.007723f
C5951 commonsourceibias.n191 gnd 0.010462f
C5952 commonsourceibias.n192 gnd 0.057575f
C5953 commonsourceibias.n193 gnd 0.010531f
C5954 commonsourceibias.n194 gnd 0.009519f
C5955 commonsourceibias.n195 gnd 0.007723f
C5956 commonsourceibias.n196 gnd 0.007723f
C5957 commonsourceibias.n197 gnd 0.007835f
C5958 commonsourceibias.n198 gnd 0.0081f
C5959 commonsourceibias.t61 gnd 0.156059f
C5960 commonsourceibias.n199 gnd 0.068889f
C5961 commonsourceibias.n200 gnd 0.023444f
C5962 commonsourceibias.n201 gnd 0.388889f
C5963 commonsourceibias.n202 gnd 0.010306f
C5964 commonsourceibias.t84 gnd 0.156059f
C5965 commonsourceibias.t92 gnd 0.144299f
C5966 commonsourceibias.n203 gnd 0.057575f
C5967 commonsourceibias.n204 gnd 0.007723f
C5968 commonsourceibias.t51 gnd 0.144299f
C5969 commonsourceibias.n205 gnd 0.006248f
C5970 commonsourceibias.n206 gnd 0.007723f
C5971 commonsourceibias.t63 gnd 0.144299f
C5972 commonsourceibias.n207 gnd 0.007456f
C5973 commonsourceibias.n208 gnd 0.007723f
C5974 commonsourceibias.t48 gnd 0.144299f
C5975 commonsourceibias.n209 gnd 0.006238f
C5976 commonsourceibias.n210 gnd 0.007723f
C5977 commonsourceibias.t94 gnd 0.144299f
C5978 commonsourceibias.t83 gnd 0.144299f
C5979 commonsourceibias.n211 gnd 0.057575f
C5980 commonsourceibias.n212 gnd 0.007723f
C5981 commonsourceibias.t80 gnd 0.144299f
C5982 commonsourceibias.n213 gnd 0.057575f
C5983 commonsourceibias.n214 gnd 0.007723f
C5984 commonsourceibias.t90 gnd 0.144299f
C5985 commonsourceibias.n215 gnd 0.057575f
C5986 commonsourceibias.n216 gnd 0.038882f
C5987 commonsourceibias.t59 gnd 0.144299f
C5988 commonsourceibias.t75 gnd 0.162824f
C5989 commonsourceibias.n217 gnd 0.066816f
C5990 commonsourceibias.n218 gnd 0.069172f
C5991 commonsourceibias.n219 gnd 0.009519f
C5992 commonsourceibias.n220 gnd 0.010531f
C5993 commonsourceibias.n221 gnd 0.007723f
C5994 commonsourceibias.n222 gnd 0.007723f
C5995 commonsourceibias.n223 gnd 0.010462f
C5996 commonsourceibias.n224 gnd 0.006248f
C5997 commonsourceibias.n225 gnd 0.010592f
C5998 commonsourceibias.n226 gnd 0.007723f
C5999 commonsourceibias.n227 gnd 0.007723f
C6000 commonsourceibias.n228 gnd 0.010657f
C6001 commonsourceibias.n229 gnd 0.009189f
C6002 commonsourceibias.n230 gnd 0.007456f
C6003 commonsourceibias.n231 gnd 0.007723f
C6004 commonsourceibias.n232 gnd 0.007723f
C6005 commonsourceibias.n233 gnd 0.009447f
C6006 commonsourceibias.n234 gnd 0.010603f
C6007 commonsourceibias.n235 gnd 0.057575f
C6008 commonsourceibias.n236 gnd 0.010532f
C6009 commonsourceibias.n237 gnd 0.007686f
C6010 commonsourceibias.t27 gnd 0.016666f
C6011 commonsourceibias.t43 gnd 0.016666f
C6012 commonsourceibias.n238 gnd 0.147764f
C6013 commonsourceibias.t21 gnd 0.016666f
C6014 commonsourceibias.t39 gnd 0.016666f
C6015 commonsourceibias.n239 gnd 0.147271f
C6016 commonsourceibias.n240 gnd 0.137229f
C6017 commonsourceibias.t7 gnd 0.016666f
C6018 commonsourceibias.t31 gnd 0.016666f
C6019 commonsourceibias.n241 gnd 0.147271f
C6020 commonsourceibias.n242 gnd 0.056516f
C6021 commonsourceibias.n243 gnd 0.010306f
C6022 commonsourceibias.t24 gnd 0.144299f
C6023 commonsourceibias.n244 gnd 0.057575f
C6024 commonsourceibias.n245 gnd 0.007723f
C6025 commonsourceibias.t2 gnd 0.144299f
C6026 commonsourceibias.n246 gnd 0.006248f
C6027 commonsourceibias.n247 gnd 0.007723f
C6028 commonsourceibias.t34 gnd 0.144299f
C6029 commonsourceibias.n248 gnd 0.007456f
C6030 commonsourceibias.n249 gnd 0.007723f
C6031 commonsourceibias.t40 gnd 0.144299f
C6032 commonsourceibias.n250 gnd 0.006238f
C6033 commonsourceibias.n251 gnd 0.007723f
C6034 commonsourceibias.t30 gnd 0.144299f
C6035 commonsourceibias.t6 gnd 0.144299f
C6036 commonsourceibias.n252 gnd 0.057575f
C6037 commonsourceibias.n253 gnd 0.007723f
C6038 commonsourceibias.t38 gnd 0.144299f
C6039 commonsourceibias.n254 gnd 0.057575f
C6040 commonsourceibias.n255 gnd 0.007723f
C6041 commonsourceibias.t20 gnd 0.144299f
C6042 commonsourceibias.n256 gnd 0.057575f
C6043 commonsourceibias.n257 gnd 0.038882f
C6044 commonsourceibias.t42 gnd 0.144299f
C6045 commonsourceibias.t26 gnd 0.162824f
C6046 commonsourceibias.n258 gnd 0.066816f
C6047 commonsourceibias.n259 gnd 0.069172f
C6048 commonsourceibias.n260 gnd 0.009519f
C6049 commonsourceibias.n261 gnd 0.010531f
C6050 commonsourceibias.n262 gnd 0.007723f
C6051 commonsourceibias.n263 gnd 0.007723f
C6052 commonsourceibias.n264 gnd 0.010462f
C6053 commonsourceibias.n265 gnd 0.006248f
C6054 commonsourceibias.n266 gnd 0.010592f
C6055 commonsourceibias.n267 gnd 0.007723f
C6056 commonsourceibias.n268 gnd 0.007723f
C6057 commonsourceibias.n269 gnd 0.010657f
C6058 commonsourceibias.n270 gnd 0.009189f
C6059 commonsourceibias.n271 gnd 0.007456f
C6060 commonsourceibias.n272 gnd 0.007723f
C6061 commonsourceibias.n273 gnd 0.007723f
C6062 commonsourceibias.n274 gnd 0.009447f
C6063 commonsourceibias.n275 gnd 0.010603f
C6064 commonsourceibias.n276 gnd 0.057575f
C6065 commonsourceibias.n277 gnd 0.010532f
C6066 commonsourceibias.n278 gnd 0.007723f
C6067 commonsourceibias.n279 gnd 0.007723f
C6068 commonsourceibias.n280 gnd 0.007723f
C6069 commonsourceibias.n281 gnd 0.010532f
C6070 commonsourceibias.n282 gnd 0.057575f
C6071 commonsourceibias.n283 gnd 0.010603f
C6072 commonsourceibias.t12 gnd 0.144299f
C6073 commonsourceibias.n284 gnd 0.057575f
C6074 commonsourceibias.n285 gnd 0.009447f
C6075 commonsourceibias.n286 gnd 0.007723f
C6076 commonsourceibias.n287 gnd 0.007723f
C6077 commonsourceibias.n288 gnd 0.007723f
C6078 commonsourceibias.n289 gnd 0.009189f
C6079 commonsourceibias.n290 gnd 0.010657f
C6080 commonsourceibias.n291 gnd 0.057575f
C6081 commonsourceibias.n292 gnd 0.010592f
C6082 commonsourceibias.n293 gnd 0.007723f
C6083 commonsourceibias.n294 gnd 0.007723f
C6084 commonsourceibias.n295 gnd 0.007723f
C6085 commonsourceibias.n296 gnd 0.010462f
C6086 commonsourceibias.n297 gnd 0.057575f
C6087 commonsourceibias.n298 gnd 0.010531f
C6088 commonsourceibias.n299 gnd 0.009519f
C6089 commonsourceibias.n300 gnd 0.007723f
C6090 commonsourceibias.n301 gnd 0.007723f
C6091 commonsourceibias.n302 gnd 0.007835f
C6092 commonsourceibias.n303 gnd 0.0081f
C6093 commonsourceibias.t36 gnd 0.156059f
C6094 commonsourceibias.n304 gnd 0.068889f
C6095 commonsourceibias.n305 gnd 0.076422f
C6096 commonsourceibias.t25 gnd 0.016666f
C6097 commonsourceibias.t37 gnd 0.016666f
C6098 commonsourceibias.n306 gnd 0.147271f
C6099 commonsourceibias.n307 gnd 0.127253f
C6100 commonsourceibias.t35 gnd 0.016666f
C6101 commonsourceibias.t3 gnd 0.016666f
C6102 commonsourceibias.n308 gnd 0.147271f
C6103 commonsourceibias.n309 gnd 0.067647f
C6104 commonsourceibias.t41 gnd 0.016666f
C6105 commonsourceibias.t13 gnd 0.016666f
C6106 commonsourceibias.n310 gnd 0.147271f
C6107 commonsourceibias.n311 gnd 0.056516f
C6108 commonsourceibias.n312 gnd 0.068435f
C6109 commonsourceibias.n313 gnd 0.055832f
C6110 commonsourceibias.n314 gnd 0.007686f
C6111 commonsourceibias.n315 gnd 0.010532f
C6112 commonsourceibias.n316 gnd 0.057575f
C6113 commonsourceibias.n317 gnd 0.010603f
C6114 commonsourceibias.t88 gnd 0.144299f
C6115 commonsourceibias.n318 gnd 0.057575f
C6116 commonsourceibias.n319 gnd 0.009447f
C6117 commonsourceibias.n320 gnd 0.007723f
C6118 commonsourceibias.n321 gnd 0.007723f
C6119 commonsourceibias.n322 gnd 0.007723f
C6120 commonsourceibias.n323 gnd 0.009189f
C6121 commonsourceibias.n324 gnd 0.010657f
C6122 commonsourceibias.n325 gnd 0.057575f
C6123 commonsourceibias.n326 gnd 0.010592f
C6124 commonsourceibias.n327 gnd 0.007723f
C6125 commonsourceibias.n328 gnd 0.007723f
C6126 commonsourceibias.n329 gnd 0.007723f
C6127 commonsourceibias.n330 gnd 0.010462f
C6128 commonsourceibias.n331 gnd 0.057575f
C6129 commonsourceibias.n332 gnd 0.010531f
C6130 commonsourceibias.n333 gnd 0.009519f
C6131 commonsourceibias.n334 gnd 0.007723f
C6132 commonsourceibias.n335 gnd 0.007723f
C6133 commonsourceibias.n336 gnd 0.007835f
C6134 commonsourceibias.n337 gnd 0.0081f
C6135 commonsourceibias.n338 gnd 0.068889f
C6136 commonsourceibias.n339 gnd 0.044582f
C6137 commonsourceibias.n340 gnd 0.010306f
C6138 commonsourceibias.t85 gnd 0.144299f
C6139 commonsourceibias.n341 gnd 0.057575f
C6140 commonsourceibias.n342 gnd 0.007723f
C6141 commonsourceibias.t93 gnd 0.144299f
C6142 commonsourceibias.n343 gnd 0.006248f
C6143 commonsourceibias.n344 gnd 0.007723f
C6144 commonsourceibias.t56 gnd 0.144299f
C6145 commonsourceibias.n345 gnd 0.007456f
C6146 commonsourceibias.n346 gnd 0.007723f
C6147 commonsourceibias.t89 gnd 0.144299f
C6148 commonsourceibias.n347 gnd 0.006238f
C6149 commonsourceibias.n348 gnd 0.007723f
C6150 commonsourceibias.t86 gnd 0.144299f
C6151 commonsourceibias.t73 gnd 0.144299f
C6152 commonsourceibias.n349 gnd 0.057575f
C6153 commonsourceibias.n350 gnd 0.007723f
C6154 commonsourceibias.t69 gnd 0.144299f
C6155 commonsourceibias.n351 gnd 0.057575f
C6156 commonsourceibias.n352 gnd 0.007723f
C6157 commonsourceibias.t82 gnd 0.144299f
C6158 commonsourceibias.n353 gnd 0.057575f
C6159 commonsourceibias.n354 gnd 0.038882f
C6160 commonsourceibias.t52 gnd 0.144299f
C6161 commonsourceibias.t64 gnd 0.162824f
C6162 commonsourceibias.n355 gnd 0.066816f
C6163 commonsourceibias.n356 gnd 0.069172f
C6164 commonsourceibias.n357 gnd 0.009519f
C6165 commonsourceibias.n358 gnd 0.010531f
C6166 commonsourceibias.n359 gnd 0.007723f
C6167 commonsourceibias.n360 gnd 0.007723f
C6168 commonsourceibias.n361 gnd 0.010462f
C6169 commonsourceibias.n362 gnd 0.006248f
C6170 commonsourceibias.n363 gnd 0.010592f
C6171 commonsourceibias.n364 gnd 0.007723f
C6172 commonsourceibias.n365 gnd 0.007723f
C6173 commonsourceibias.n366 gnd 0.010657f
C6174 commonsourceibias.n367 gnd 0.009189f
C6175 commonsourceibias.n368 gnd 0.007456f
C6176 commonsourceibias.n369 gnd 0.007723f
C6177 commonsourceibias.n370 gnd 0.007723f
C6178 commonsourceibias.n371 gnd 0.009447f
C6179 commonsourceibias.n372 gnd 0.010603f
C6180 commonsourceibias.n373 gnd 0.057575f
C6181 commonsourceibias.n374 gnd 0.010532f
C6182 commonsourceibias.n375 gnd 0.007723f
C6183 commonsourceibias.n376 gnd 0.007723f
C6184 commonsourceibias.n377 gnd 0.007723f
C6185 commonsourceibias.n378 gnd 0.010532f
C6186 commonsourceibias.n379 gnd 0.057575f
C6187 commonsourceibias.n380 gnd 0.010603f
C6188 commonsourceibias.t79 gnd 0.144299f
C6189 commonsourceibias.n381 gnd 0.057575f
C6190 commonsourceibias.n382 gnd 0.009447f
C6191 commonsourceibias.n383 gnd 0.007723f
C6192 commonsourceibias.n384 gnd 0.007723f
C6193 commonsourceibias.n385 gnd 0.007723f
C6194 commonsourceibias.n386 gnd 0.009189f
C6195 commonsourceibias.n387 gnd 0.010657f
C6196 commonsourceibias.n388 gnd 0.057575f
C6197 commonsourceibias.n389 gnd 0.010592f
C6198 commonsourceibias.n390 gnd 0.007723f
C6199 commonsourceibias.n391 gnd 0.007723f
C6200 commonsourceibias.n392 gnd 0.007723f
C6201 commonsourceibias.n393 gnd 0.010462f
C6202 commonsourceibias.n394 gnd 0.057575f
C6203 commonsourceibias.n395 gnd 0.010531f
C6204 commonsourceibias.n396 gnd 0.009519f
C6205 commonsourceibias.n397 gnd 0.007723f
C6206 commonsourceibias.n398 gnd 0.007723f
C6207 commonsourceibias.n399 gnd 0.007835f
C6208 commonsourceibias.n400 gnd 0.0081f
C6209 commonsourceibias.t74 gnd 0.156059f
C6210 commonsourceibias.n401 gnd 0.068889f
C6211 commonsourceibias.n402 gnd 0.023444f
C6212 commonsourceibias.n403 gnd 0.213098f
C6213 commonsourceibias.n404 gnd 4.20869f
.ends

