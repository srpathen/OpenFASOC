* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t41 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X1 source.t43 plus.t1 drain_left.t22 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X2 a_n2874_n2088# a_n2874_n2088# a_n2874_n2088# a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.5
X3 drain_right.t23 minus.t0 source.t19 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X4 source.t38 plus.t2 drain_left.t21 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X5 drain_left.t20 plus.t3 source.t39 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X6 source.t42 plus.t4 drain_left.t19 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X7 source.t4 minus.t1 drain_right.t22 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X8 drain_right.t21 minus.t2 source.t11 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X9 source.t3 minus.t3 drain_right.t20 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X10 source.t7 minus.t4 drain_right.t19 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X11 source.t22 plus.t5 drain_left.t18 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X12 source.t28 plus.t6 drain_left.t17 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X13 source.t5 minus.t5 drain_right.t18 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X14 source.t20 minus.t6 drain_right.t17 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X15 drain_right.t16 minus.t7 source.t13 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X16 drain_right.t15 minus.t8 source.t12 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X17 drain_right.t14 minus.t9 source.t46 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X18 a_n2874_n2088# a_n2874_n2088# a_n2874_n2088# a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X19 drain_left.t16 plus.t7 source.t25 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X20 drain_right.t13 minus.t10 source.t47 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X21 source.t44 plus.t8 drain_left.t15 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X22 source.t34 plus.t9 drain_left.t14 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X23 source.t6 minus.t11 drain_right.t12 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X24 source.t0 minus.t12 drain_right.t11 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X25 drain_left.t13 plus.t10 source.t23 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X26 source.t29 plus.t11 drain_left.t12 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X27 source.t36 plus.t12 drain_left.t11 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X28 drain_left.t10 plus.t13 source.t24 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X29 drain_right.t10 minus.t13 source.t21 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X30 drain_right.t9 minus.t14 source.t15 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X31 a_n2874_n2088# a_n2874_n2088# a_n2874_n2088# a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X32 source.t18 minus.t15 drain_right.t8 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X33 drain_right.t7 minus.t16 source.t9 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X34 source.t37 plus.t14 drain_left.t9 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X35 drain_left.t8 plus.t15 source.t30 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X36 drain_left.t7 plus.t16 source.t45 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X37 drain_right.t6 minus.t17 source.t14 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X38 drain_right.t5 minus.t18 source.t17 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X39 source.t8 minus.t19 drain_right.t4 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X40 source.t10 minus.t20 drain_right.t3 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X41 drain_left.t6 plus.t17 source.t26 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X42 source.t31 plus.t18 drain_left.t5 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X43 source.t1 minus.t21 drain_right.t2 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X44 drain_left.t4 plus.t19 source.t32 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X45 source.t2 minus.t22 drain_right.t1 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X46 drain_left.t3 plus.t20 source.t33 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X47 source.t27 plus.t21 drain_left.t2 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X48 drain_left.t1 plus.t22 source.t35 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X49 drain_left.t0 plus.t23 source.t40 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X50 drain_right.t0 minus.t23 source.t16 a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X51 a_n2874_n2088# a_n2874_n2088# a_n2874_n2088# a_n2874_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
R0 plus.n11 plus.t6 394.125
R1 plus.n45 plus.t10 394.125
R2 plus.n32 plus.t3 367.767
R3 plus.n30 plus.t4 367.767
R4 plus.n29 plus.t13 367.767
R5 plus.n3 plus.t5 367.767
R6 plus.n23 plus.t20 367.767
R7 plus.n22 plus.t9 367.767
R8 plus.n6 plus.t23 367.767
R9 plus.n17 plus.t18 367.767
R10 plus.n15 plus.t7 367.767
R11 plus.n9 plus.t21 367.767
R12 plus.n10 plus.t16 367.767
R13 plus.n66 plus.t8 367.767
R14 plus.n64 plus.t17 367.767
R15 plus.n63 plus.t1 367.767
R16 plus.n37 plus.t0 367.767
R17 plus.n57 plus.t12 367.767
R18 plus.n56 plus.t19 367.767
R19 plus.n40 plus.t2 367.767
R20 plus.n51 plus.t15 367.767
R21 plus.n49 plus.t14 367.767
R22 plus.n43 plus.t22 367.767
R23 plus.n44 plus.t11 367.767
R24 plus.n12 plus.n9 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n15 plus.n8 161.3
R27 plus.n16 plus.n7 161.3
R28 plus.n18 plus.n17 161.3
R29 plus.n19 plus.n6 161.3
R30 plus.n21 plus.n20 161.3
R31 plus.n22 plus.n5 161.3
R32 plus.n23 plus.n4 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n26 plus.n3 161.3
R35 plus.n28 plus.n27 161.3
R36 plus.n29 plus.n2 161.3
R37 plus.n30 plus.n1 161.3
R38 plus.n31 plus.n0 161.3
R39 plus.n33 plus.n32 161.3
R40 plus.n46 plus.n43 161.3
R41 plus.n48 plus.n47 161.3
R42 plus.n49 plus.n42 161.3
R43 plus.n50 plus.n41 161.3
R44 plus.n52 plus.n51 161.3
R45 plus.n53 plus.n40 161.3
R46 plus.n55 plus.n54 161.3
R47 plus.n56 plus.n39 161.3
R48 plus.n57 plus.n38 161.3
R49 plus.n59 plus.n58 161.3
R50 plus.n60 plus.n37 161.3
R51 plus.n62 plus.n61 161.3
R52 plus.n63 plus.n36 161.3
R53 plus.n64 plus.n35 161.3
R54 plus.n65 plus.n34 161.3
R55 plus.n67 plus.n66 161.3
R56 plus.n30 plus.n29 48.2005
R57 plus.n23 plus.n22 48.2005
R58 plus.n17 plus.n6 48.2005
R59 plus.n10 plus.n9 48.2005
R60 plus.n64 plus.n63 48.2005
R61 plus.n57 plus.n56 48.2005
R62 plus.n51 plus.n40 48.2005
R63 plus.n44 plus.n43 48.2005
R64 plus.n24 plus.n3 47.4702
R65 plus.n16 plus.n15 47.4702
R66 plus.n58 plus.n37 47.4702
R67 plus.n50 plus.n49 47.4702
R68 plus.n32 plus.n31 46.0096
R69 plus.n66 plus.n65 46.0096
R70 plus.n12 plus.n11 45.0871
R71 plus.n46 plus.n45 45.0871
R72 plus plus.n67 31.643
R73 plus.n28 plus.n3 25.5611
R74 plus.n15 plus.n14 25.5611
R75 plus.n62 plus.n37 25.5611
R76 plus.n49 plus.n48 25.5611
R77 plus.n21 plus.n6 24.1005
R78 plus.n22 plus.n21 24.1005
R79 plus.n56 plus.n55 24.1005
R80 plus.n55 plus.n40 24.1005
R81 plus.n29 plus.n28 22.6399
R82 plus.n14 plus.n9 22.6399
R83 plus.n63 plus.n62 22.6399
R84 plus.n48 plus.n43 22.6399
R85 plus.n11 plus.n10 14.1472
R86 plus.n45 plus.n44 14.1472
R87 plus plus.n33 9.89823
R88 plus.n31 plus.n30 2.19141
R89 plus.n65 plus.n64 2.19141
R90 plus.n24 plus.n23 0.730803
R91 plus.n17 plus.n16 0.730803
R92 plus.n58 plus.n57 0.730803
R93 plus.n51 plus.n50 0.730803
R94 plus.n13 plus.n12 0.189894
R95 plus.n13 plus.n8 0.189894
R96 plus.n8 plus.n7 0.189894
R97 plus.n18 plus.n7 0.189894
R98 plus.n19 plus.n18 0.189894
R99 plus.n20 plus.n19 0.189894
R100 plus.n20 plus.n5 0.189894
R101 plus.n5 plus.n4 0.189894
R102 plus.n25 plus.n4 0.189894
R103 plus.n26 plus.n25 0.189894
R104 plus.n27 plus.n26 0.189894
R105 plus.n27 plus.n2 0.189894
R106 plus.n2 plus.n1 0.189894
R107 plus.n1 plus.n0 0.189894
R108 plus.n33 plus.n0 0.189894
R109 plus.n67 plus.n34 0.189894
R110 plus.n35 plus.n34 0.189894
R111 plus.n36 plus.n35 0.189894
R112 plus.n61 plus.n36 0.189894
R113 plus.n61 plus.n60 0.189894
R114 plus.n60 plus.n59 0.189894
R115 plus.n59 plus.n38 0.189894
R116 plus.n39 plus.n38 0.189894
R117 plus.n54 plus.n39 0.189894
R118 plus.n54 plus.n53 0.189894
R119 plus.n53 plus.n52 0.189894
R120 plus.n52 plus.n41 0.189894
R121 plus.n42 plus.n41 0.189894
R122 plus.n47 plus.n42 0.189894
R123 plus.n47 plus.n46 0.189894
R124 source.n290 source.n264 289.615
R125 source.n248 source.n222 289.615
R126 source.n216 source.n190 289.615
R127 source.n174 source.n148 289.615
R128 source.n26 source.n0 289.615
R129 source.n68 source.n42 289.615
R130 source.n100 source.n74 289.615
R131 source.n142 source.n116 289.615
R132 source.n275 source.n274 185
R133 source.n272 source.n271 185
R134 source.n281 source.n280 185
R135 source.n283 source.n282 185
R136 source.n268 source.n267 185
R137 source.n289 source.n288 185
R138 source.n291 source.n290 185
R139 source.n233 source.n232 185
R140 source.n230 source.n229 185
R141 source.n239 source.n238 185
R142 source.n241 source.n240 185
R143 source.n226 source.n225 185
R144 source.n247 source.n246 185
R145 source.n249 source.n248 185
R146 source.n201 source.n200 185
R147 source.n198 source.n197 185
R148 source.n207 source.n206 185
R149 source.n209 source.n208 185
R150 source.n194 source.n193 185
R151 source.n215 source.n214 185
R152 source.n217 source.n216 185
R153 source.n159 source.n158 185
R154 source.n156 source.n155 185
R155 source.n165 source.n164 185
R156 source.n167 source.n166 185
R157 source.n152 source.n151 185
R158 source.n173 source.n172 185
R159 source.n175 source.n174 185
R160 source.n27 source.n26 185
R161 source.n25 source.n24 185
R162 source.n4 source.n3 185
R163 source.n19 source.n18 185
R164 source.n17 source.n16 185
R165 source.n8 source.n7 185
R166 source.n11 source.n10 185
R167 source.n69 source.n68 185
R168 source.n67 source.n66 185
R169 source.n46 source.n45 185
R170 source.n61 source.n60 185
R171 source.n59 source.n58 185
R172 source.n50 source.n49 185
R173 source.n53 source.n52 185
R174 source.n101 source.n100 185
R175 source.n99 source.n98 185
R176 source.n78 source.n77 185
R177 source.n93 source.n92 185
R178 source.n91 source.n90 185
R179 source.n82 source.n81 185
R180 source.n85 source.n84 185
R181 source.n143 source.n142 185
R182 source.n141 source.n140 185
R183 source.n120 source.n119 185
R184 source.n135 source.n134 185
R185 source.n133 source.n132 185
R186 source.n124 source.n123 185
R187 source.n127 source.n126 185
R188 source.t9 source.n273 147.661
R189 source.t8 source.n231 147.661
R190 source.t23 source.n199 147.661
R191 source.t44 source.n157 147.661
R192 source.t39 source.n9 147.661
R193 source.t28 source.n51 147.661
R194 source.t21 source.n83 147.661
R195 source.t2 source.n125 147.661
R196 source.n274 source.n271 104.615
R197 source.n281 source.n271 104.615
R198 source.n282 source.n281 104.615
R199 source.n282 source.n267 104.615
R200 source.n289 source.n267 104.615
R201 source.n290 source.n289 104.615
R202 source.n232 source.n229 104.615
R203 source.n239 source.n229 104.615
R204 source.n240 source.n239 104.615
R205 source.n240 source.n225 104.615
R206 source.n247 source.n225 104.615
R207 source.n248 source.n247 104.615
R208 source.n200 source.n197 104.615
R209 source.n207 source.n197 104.615
R210 source.n208 source.n207 104.615
R211 source.n208 source.n193 104.615
R212 source.n215 source.n193 104.615
R213 source.n216 source.n215 104.615
R214 source.n158 source.n155 104.615
R215 source.n165 source.n155 104.615
R216 source.n166 source.n165 104.615
R217 source.n166 source.n151 104.615
R218 source.n173 source.n151 104.615
R219 source.n174 source.n173 104.615
R220 source.n26 source.n25 104.615
R221 source.n25 source.n3 104.615
R222 source.n18 source.n3 104.615
R223 source.n18 source.n17 104.615
R224 source.n17 source.n7 104.615
R225 source.n10 source.n7 104.615
R226 source.n68 source.n67 104.615
R227 source.n67 source.n45 104.615
R228 source.n60 source.n45 104.615
R229 source.n60 source.n59 104.615
R230 source.n59 source.n49 104.615
R231 source.n52 source.n49 104.615
R232 source.n100 source.n99 104.615
R233 source.n99 source.n77 104.615
R234 source.n92 source.n77 104.615
R235 source.n92 source.n91 104.615
R236 source.n91 source.n81 104.615
R237 source.n84 source.n81 104.615
R238 source.n142 source.n141 104.615
R239 source.n141 source.n119 104.615
R240 source.n134 source.n119 104.615
R241 source.n134 source.n133 104.615
R242 source.n133 source.n123 104.615
R243 source.n126 source.n123 104.615
R244 source.n274 source.t9 52.3082
R245 source.n232 source.t8 52.3082
R246 source.n200 source.t23 52.3082
R247 source.n158 source.t44 52.3082
R248 source.n10 source.t39 52.3082
R249 source.n52 source.t28 52.3082
R250 source.n84 source.t21 52.3082
R251 source.n126 source.t2 52.3082
R252 source.n33 source.n32 50.512
R253 source.n35 source.n34 50.512
R254 source.n37 source.n36 50.512
R255 source.n39 source.n38 50.512
R256 source.n41 source.n40 50.512
R257 source.n107 source.n106 50.512
R258 source.n109 source.n108 50.512
R259 source.n111 source.n110 50.512
R260 source.n113 source.n112 50.512
R261 source.n115 source.n114 50.512
R262 source.n263 source.n262 50.5119
R263 source.n261 source.n260 50.5119
R264 source.n259 source.n258 50.5119
R265 source.n257 source.n256 50.5119
R266 source.n255 source.n254 50.5119
R267 source.n189 source.n188 50.5119
R268 source.n187 source.n186 50.5119
R269 source.n185 source.n184 50.5119
R270 source.n183 source.n182 50.5119
R271 source.n181 source.n180 50.5119
R272 source.n295 source.n294 32.1853
R273 source.n253 source.n252 32.1853
R274 source.n221 source.n220 32.1853
R275 source.n179 source.n178 32.1853
R276 source.n31 source.n30 32.1853
R277 source.n73 source.n72 32.1853
R278 source.n105 source.n104 32.1853
R279 source.n147 source.n146 32.1853
R280 source.n179 source.n147 17.4578
R281 source.n275 source.n273 15.6674
R282 source.n233 source.n231 15.6674
R283 source.n201 source.n199 15.6674
R284 source.n159 source.n157 15.6674
R285 source.n11 source.n9 15.6674
R286 source.n53 source.n51 15.6674
R287 source.n85 source.n83 15.6674
R288 source.n127 source.n125 15.6674
R289 source.n276 source.n272 12.8005
R290 source.n234 source.n230 12.8005
R291 source.n202 source.n198 12.8005
R292 source.n160 source.n156 12.8005
R293 source.n12 source.n8 12.8005
R294 source.n54 source.n50 12.8005
R295 source.n86 source.n82 12.8005
R296 source.n128 source.n124 12.8005
R297 source.n280 source.n279 12.0247
R298 source.n238 source.n237 12.0247
R299 source.n206 source.n205 12.0247
R300 source.n164 source.n163 12.0247
R301 source.n16 source.n15 12.0247
R302 source.n58 source.n57 12.0247
R303 source.n90 source.n89 12.0247
R304 source.n132 source.n131 12.0247
R305 source.n296 source.n31 11.8371
R306 source.n283 source.n270 11.249
R307 source.n241 source.n228 11.249
R308 source.n209 source.n196 11.249
R309 source.n167 source.n154 11.249
R310 source.n19 source.n6 11.249
R311 source.n61 source.n48 11.249
R312 source.n93 source.n80 11.249
R313 source.n135 source.n122 11.249
R314 source.n284 source.n268 10.4732
R315 source.n242 source.n226 10.4732
R316 source.n210 source.n194 10.4732
R317 source.n168 source.n152 10.4732
R318 source.n20 source.n4 10.4732
R319 source.n62 source.n46 10.4732
R320 source.n94 source.n78 10.4732
R321 source.n136 source.n120 10.4732
R322 source.n288 source.n287 9.69747
R323 source.n246 source.n245 9.69747
R324 source.n214 source.n213 9.69747
R325 source.n172 source.n171 9.69747
R326 source.n24 source.n23 9.69747
R327 source.n66 source.n65 9.69747
R328 source.n98 source.n97 9.69747
R329 source.n140 source.n139 9.69747
R330 source.n294 source.n293 9.45567
R331 source.n252 source.n251 9.45567
R332 source.n220 source.n219 9.45567
R333 source.n178 source.n177 9.45567
R334 source.n30 source.n29 9.45567
R335 source.n72 source.n71 9.45567
R336 source.n104 source.n103 9.45567
R337 source.n146 source.n145 9.45567
R338 source.n293 source.n292 9.3005
R339 source.n266 source.n265 9.3005
R340 source.n287 source.n286 9.3005
R341 source.n285 source.n284 9.3005
R342 source.n270 source.n269 9.3005
R343 source.n279 source.n278 9.3005
R344 source.n277 source.n276 9.3005
R345 source.n251 source.n250 9.3005
R346 source.n224 source.n223 9.3005
R347 source.n245 source.n244 9.3005
R348 source.n243 source.n242 9.3005
R349 source.n228 source.n227 9.3005
R350 source.n237 source.n236 9.3005
R351 source.n235 source.n234 9.3005
R352 source.n219 source.n218 9.3005
R353 source.n192 source.n191 9.3005
R354 source.n213 source.n212 9.3005
R355 source.n211 source.n210 9.3005
R356 source.n196 source.n195 9.3005
R357 source.n205 source.n204 9.3005
R358 source.n203 source.n202 9.3005
R359 source.n177 source.n176 9.3005
R360 source.n150 source.n149 9.3005
R361 source.n171 source.n170 9.3005
R362 source.n169 source.n168 9.3005
R363 source.n154 source.n153 9.3005
R364 source.n163 source.n162 9.3005
R365 source.n161 source.n160 9.3005
R366 source.n29 source.n28 9.3005
R367 source.n2 source.n1 9.3005
R368 source.n23 source.n22 9.3005
R369 source.n21 source.n20 9.3005
R370 source.n6 source.n5 9.3005
R371 source.n15 source.n14 9.3005
R372 source.n13 source.n12 9.3005
R373 source.n71 source.n70 9.3005
R374 source.n44 source.n43 9.3005
R375 source.n65 source.n64 9.3005
R376 source.n63 source.n62 9.3005
R377 source.n48 source.n47 9.3005
R378 source.n57 source.n56 9.3005
R379 source.n55 source.n54 9.3005
R380 source.n103 source.n102 9.3005
R381 source.n76 source.n75 9.3005
R382 source.n97 source.n96 9.3005
R383 source.n95 source.n94 9.3005
R384 source.n80 source.n79 9.3005
R385 source.n89 source.n88 9.3005
R386 source.n87 source.n86 9.3005
R387 source.n145 source.n144 9.3005
R388 source.n118 source.n117 9.3005
R389 source.n139 source.n138 9.3005
R390 source.n137 source.n136 9.3005
R391 source.n122 source.n121 9.3005
R392 source.n131 source.n130 9.3005
R393 source.n129 source.n128 9.3005
R394 source.n291 source.n266 8.92171
R395 source.n249 source.n224 8.92171
R396 source.n217 source.n192 8.92171
R397 source.n175 source.n150 8.92171
R398 source.n27 source.n2 8.92171
R399 source.n69 source.n44 8.92171
R400 source.n101 source.n76 8.92171
R401 source.n143 source.n118 8.92171
R402 source.n292 source.n264 8.14595
R403 source.n250 source.n222 8.14595
R404 source.n218 source.n190 8.14595
R405 source.n176 source.n148 8.14595
R406 source.n28 source.n0 8.14595
R407 source.n70 source.n42 8.14595
R408 source.n102 source.n74 8.14595
R409 source.n144 source.n116 8.14595
R410 source.n294 source.n264 5.81868
R411 source.n252 source.n222 5.81868
R412 source.n220 source.n190 5.81868
R413 source.n178 source.n148 5.81868
R414 source.n30 source.n0 5.81868
R415 source.n72 source.n42 5.81868
R416 source.n104 source.n74 5.81868
R417 source.n146 source.n116 5.81868
R418 source.n296 source.n295 5.62119
R419 source.n292 source.n291 5.04292
R420 source.n250 source.n249 5.04292
R421 source.n218 source.n217 5.04292
R422 source.n176 source.n175 5.04292
R423 source.n28 source.n27 5.04292
R424 source.n70 source.n69 5.04292
R425 source.n102 source.n101 5.04292
R426 source.n144 source.n143 5.04292
R427 source.n277 source.n273 4.38594
R428 source.n235 source.n231 4.38594
R429 source.n203 source.n199 4.38594
R430 source.n161 source.n157 4.38594
R431 source.n13 source.n9 4.38594
R432 source.n55 source.n51 4.38594
R433 source.n87 source.n83 4.38594
R434 source.n129 source.n125 4.38594
R435 source.n288 source.n266 4.26717
R436 source.n246 source.n224 4.26717
R437 source.n214 source.n192 4.26717
R438 source.n172 source.n150 4.26717
R439 source.n24 source.n2 4.26717
R440 source.n66 source.n44 4.26717
R441 source.n98 source.n76 4.26717
R442 source.n140 source.n118 4.26717
R443 source.n287 source.n268 3.49141
R444 source.n245 source.n226 3.49141
R445 source.n213 source.n194 3.49141
R446 source.n171 source.n152 3.49141
R447 source.n23 source.n4 3.49141
R448 source.n65 source.n46 3.49141
R449 source.n97 source.n78 3.49141
R450 source.n139 source.n120 3.49141
R451 source.n262 source.t47 3.3005
R452 source.n262 source.t4 3.3005
R453 source.n260 source.t16 3.3005
R454 source.n260 source.t18 3.3005
R455 source.n258 source.t13 3.3005
R456 source.n258 source.t20 3.3005
R457 source.n256 source.t11 3.3005
R458 source.n256 source.t1 3.3005
R459 source.n254 source.t17 3.3005
R460 source.n254 source.t3 3.3005
R461 source.n188 source.t35 3.3005
R462 source.n188 source.t29 3.3005
R463 source.n186 source.t30 3.3005
R464 source.n186 source.t37 3.3005
R465 source.n184 source.t32 3.3005
R466 source.n184 source.t38 3.3005
R467 source.n182 source.t41 3.3005
R468 source.n182 source.t36 3.3005
R469 source.n180 source.t26 3.3005
R470 source.n180 source.t43 3.3005
R471 source.n32 source.t24 3.3005
R472 source.n32 source.t42 3.3005
R473 source.n34 source.t33 3.3005
R474 source.n34 source.t22 3.3005
R475 source.n36 source.t40 3.3005
R476 source.n36 source.t34 3.3005
R477 source.n38 source.t25 3.3005
R478 source.n38 source.t31 3.3005
R479 source.n40 source.t45 3.3005
R480 source.n40 source.t27 3.3005
R481 source.n106 source.t46 3.3005
R482 source.n106 source.t7 3.3005
R483 source.n108 source.t12 3.3005
R484 source.n108 source.t10 3.3005
R485 source.n110 source.t19 3.3005
R486 source.n110 source.t6 3.3005
R487 source.n112 source.t14 3.3005
R488 source.n112 source.t0 3.3005
R489 source.n114 source.t15 3.3005
R490 source.n114 source.t5 3.3005
R491 source.n284 source.n283 2.71565
R492 source.n242 source.n241 2.71565
R493 source.n210 source.n209 2.71565
R494 source.n168 source.n167 2.71565
R495 source.n20 source.n19 2.71565
R496 source.n62 source.n61 2.71565
R497 source.n94 source.n93 2.71565
R498 source.n136 source.n135 2.71565
R499 source.n280 source.n270 1.93989
R500 source.n238 source.n228 1.93989
R501 source.n206 source.n196 1.93989
R502 source.n164 source.n154 1.93989
R503 source.n16 source.n6 1.93989
R504 source.n58 source.n48 1.93989
R505 source.n90 source.n80 1.93989
R506 source.n132 source.n122 1.93989
R507 source.n279 source.n272 1.16414
R508 source.n237 source.n230 1.16414
R509 source.n205 source.n198 1.16414
R510 source.n163 source.n156 1.16414
R511 source.n15 source.n8 1.16414
R512 source.n57 source.n50 1.16414
R513 source.n89 source.n82 1.16414
R514 source.n131 source.n124 1.16414
R515 source.n147 source.n115 0.716017
R516 source.n115 source.n113 0.716017
R517 source.n113 source.n111 0.716017
R518 source.n111 source.n109 0.716017
R519 source.n109 source.n107 0.716017
R520 source.n107 source.n105 0.716017
R521 source.n73 source.n41 0.716017
R522 source.n41 source.n39 0.716017
R523 source.n39 source.n37 0.716017
R524 source.n37 source.n35 0.716017
R525 source.n35 source.n33 0.716017
R526 source.n33 source.n31 0.716017
R527 source.n181 source.n179 0.716017
R528 source.n183 source.n181 0.716017
R529 source.n185 source.n183 0.716017
R530 source.n187 source.n185 0.716017
R531 source.n189 source.n187 0.716017
R532 source.n221 source.n189 0.716017
R533 source.n255 source.n253 0.716017
R534 source.n257 source.n255 0.716017
R535 source.n259 source.n257 0.716017
R536 source.n261 source.n259 0.716017
R537 source.n263 source.n261 0.716017
R538 source.n295 source.n263 0.716017
R539 source.n105 source.n73 0.470328
R540 source.n253 source.n221 0.470328
R541 source.n276 source.n275 0.388379
R542 source.n234 source.n233 0.388379
R543 source.n202 source.n201 0.388379
R544 source.n160 source.n159 0.388379
R545 source.n12 source.n11 0.388379
R546 source.n54 source.n53 0.388379
R547 source.n86 source.n85 0.388379
R548 source.n128 source.n127 0.388379
R549 source source.n296 0.188
R550 source.n278 source.n277 0.155672
R551 source.n278 source.n269 0.155672
R552 source.n285 source.n269 0.155672
R553 source.n286 source.n285 0.155672
R554 source.n286 source.n265 0.155672
R555 source.n293 source.n265 0.155672
R556 source.n236 source.n235 0.155672
R557 source.n236 source.n227 0.155672
R558 source.n243 source.n227 0.155672
R559 source.n244 source.n243 0.155672
R560 source.n244 source.n223 0.155672
R561 source.n251 source.n223 0.155672
R562 source.n204 source.n203 0.155672
R563 source.n204 source.n195 0.155672
R564 source.n211 source.n195 0.155672
R565 source.n212 source.n211 0.155672
R566 source.n212 source.n191 0.155672
R567 source.n219 source.n191 0.155672
R568 source.n162 source.n161 0.155672
R569 source.n162 source.n153 0.155672
R570 source.n169 source.n153 0.155672
R571 source.n170 source.n169 0.155672
R572 source.n170 source.n149 0.155672
R573 source.n177 source.n149 0.155672
R574 source.n29 source.n1 0.155672
R575 source.n22 source.n1 0.155672
R576 source.n22 source.n21 0.155672
R577 source.n21 source.n5 0.155672
R578 source.n14 source.n5 0.155672
R579 source.n14 source.n13 0.155672
R580 source.n71 source.n43 0.155672
R581 source.n64 source.n43 0.155672
R582 source.n64 source.n63 0.155672
R583 source.n63 source.n47 0.155672
R584 source.n56 source.n47 0.155672
R585 source.n56 source.n55 0.155672
R586 source.n103 source.n75 0.155672
R587 source.n96 source.n75 0.155672
R588 source.n96 source.n95 0.155672
R589 source.n95 source.n79 0.155672
R590 source.n88 source.n79 0.155672
R591 source.n88 source.n87 0.155672
R592 source.n145 source.n117 0.155672
R593 source.n138 source.n117 0.155672
R594 source.n138 source.n137 0.155672
R595 source.n137 source.n121 0.155672
R596 source.n130 source.n121 0.155672
R597 source.n130 source.n129 0.155672
R598 drain_left.n13 drain_left.n11 67.9063
R599 drain_left.n7 drain_left.n5 67.9062
R600 drain_left.n2 drain_left.n0 67.9062
R601 drain_left.n19 drain_left.n18 67.1908
R602 drain_left.n17 drain_left.n16 67.1908
R603 drain_left.n15 drain_left.n14 67.1908
R604 drain_left.n13 drain_left.n12 67.1908
R605 drain_left.n21 drain_left.n20 67.1907
R606 drain_left.n7 drain_left.n6 67.1907
R607 drain_left.n9 drain_left.n8 67.1907
R608 drain_left.n4 drain_left.n3 67.1907
R609 drain_left.n2 drain_left.n1 67.1907
R610 drain_left drain_left.n10 29.619
R611 drain_left drain_left.n21 6.36873
R612 drain_left.n5 drain_left.t12 3.3005
R613 drain_left.n5 drain_left.t13 3.3005
R614 drain_left.n6 drain_left.t9 3.3005
R615 drain_left.n6 drain_left.t1 3.3005
R616 drain_left.n8 drain_left.t21 3.3005
R617 drain_left.n8 drain_left.t8 3.3005
R618 drain_left.n3 drain_left.t11 3.3005
R619 drain_left.n3 drain_left.t4 3.3005
R620 drain_left.n1 drain_left.t22 3.3005
R621 drain_left.n1 drain_left.t23 3.3005
R622 drain_left.n0 drain_left.t15 3.3005
R623 drain_left.n0 drain_left.t6 3.3005
R624 drain_left.n20 drain_left.t19 3.3005
R625 drain_left.n20 drain_left.t20 3.3005
R626 drain_left.n18 drain_left.t18 3.3005
R627 drain_left.n18 drain_left.t10 3.3005
R628 drain_left.n16 drain_left.t14 3.3005
R629 drain_left.n16 drain_left.t3 3.3005
R630 drain_left.n14 drain_left.t5 3.3005
R631 drain_left.n14 drain_left.t0 3.3005
R632 drain_left.n12 drain_left.t2 3.3005
R633 drain_left.n12 drain_left.t16 3.3005
R634 drain_left.n11 drain_left.t17 3.3005
R635 drain_left.n11 drain_left.t7 3.3005
R636 drain_left.n9 drain_left.n7 0.716017
R637 drain_left.n4 drain_left.n2 0.716017
R638 drain_left.n15 drain_left.n13 0.716017
R639 drain_left.n17 drain_left.n15 0.716017
R640 drain_left.n19 drain_left.n17 0.716017
R641 drain_left.n21 drain_left.n19 0.716017
R642 drain_left.n10 drain_left.n9 0.302913
R643 drain_left.n10 drain_left.n4 0.302913
R644 minus.n9 minus.t13 394.125
R645 minus.n43 minus.t19 394.125
R646 minus.n8 minus.t4 367.767
R647 minus.n7 minus.t9 367.767
R648 minus.n13 minus.t20 367.767
R649 minus.n5 minus.t8 367.767
R650 minus.n18 minus.t11 367.767
R651 minus.n20 minus.t0 367.767
R652 minus.n3 minus.t12 367.767
R653 minus.n25 minus.t17 367.767
R654 minus.n1 minus.t5 367.767
R655 minus.n30 minus.t14 367.767
R656 minus.n32 minus.t22 367.767
R657 minus.n42 minus.t18 367.767
R658 minus.n41 minus.t3 367.767
R659 minus.n47 minus.t2 367.767
R660 minus.n39 minus.t21 367.767
R661 minus.n52 minus.t7 367.767
R662 minus.n54 minus.t6 367.767
R663 minus.n37 minus.t23 367.767
R664 minus.n59 minus.t15 367.767
R665 minus.n35 minus.t10 367.767
R666 minus.n64 minus.t1 367.767
R667 minus.n66 minus.t16 367.767
R668 minus.n33 minus.n32 161.3
R669 minus.n31 minus.n0 161.3
R670 minus.n30 minus.n29 161.3
R671 minus.n28 minus.n1 161.3
R672 minus.n27 minus.n26 161.3
R673 minus.n25 minus.n2 161.3
R674 minus.n24 minus.n23 161.3
R675 minus.n22 minus.n3 161.3
R676 minus.n21 minus.n20 161.3
R677 minus.n19 minus.n4 161.3
R678 minus.n18 minus.n17 161.3
R679 minus.n16 minus.n5 161.3
R680 minus.n15 minus.n14 161.3
R681 minus.n13 minus.n6 161.3
R682 minus.n12 minus.n11 161.3
R683 minus.n10 minus.n7 161.3
R684 minus.n67 minus.n66 161.3
R685 minus.n65 minus.n34 161.3
R686 minus.n64 minus.n63 161.3
R687 minus.n62 minus.n35 161.3
R688 minus.n61 minus.n60 161.3
R689 minus.n59 minus.n36 161.3
R690 minus.n58 minus.n57 161.3
R691 minus.n56 minus.n37 161.3
R692 minus.n55 minus.n54 161.3
R693 minus.n53 minus.n38 161.3
R694 minus.n52 minus.n51 161.3
R695 minus.n50 minus.n39 161.3
R696 minus.n49 minus.n48 161.3
R697 minus.n47 minus.n40 161.3
R698 minus.n46 minus.n45 161.3
R699 minus.n44 minus.n41 161.3
R700 minus.n8 minus.n7 48.2005
R701 minus.n18 minus.n5 48.2005
R702 minus.n20 minus.n3 48.2005
R703 minus.n30 minus.n1 48.2005
R704 minus.n42 minus.n41 48.2005
R705 minus.n52 minus.n39 48.2005
R706 minus.n54 minus.n37 48.2005
R707 minus.n64 minus.n35 48.2005
R708 minus.n14 minus.n13 47.4702
R709 minus.n25 minus.n24 47.4702
R710 minus.n48 minus.n47 47.4702
R711 minus.n59 minus.n58 47.4702
R712 minus.n32 minus.n31 46.0096
R713 minus.n66 minus.n65 46.0096
R714 minus.n10 minus.n9 45.0871
R715 minus.n44 minus.n43 45.0871
R716 minus.n68 minus.n33 35.4891
R717 minus.n13 minus.n12 25.5611
R718 minus.n26 minus.n25 25.5611
R719 minus.n47 minus.n46 25.5611
R720 minus.n60 minus.n59 25.5611
R721 minus.n20 minus.n19 24.1005
R722 minus.n19 minus.n18 24.1005
R723 minus.n53 minus.n52 24.1005
R724 minus.n54 minus.n53 24.1005
R725 minus.n12 minus.n7 22.6399
R726 minus.n26 minus.n1 22.6399
R727 minus.n46 minus.n41 22.6399
R728 minus.n60 minus.n35 22.6399
R729 minus.n9 minus.n8 14.1472
R730 minus.n43 minus.n42 14.1472
R731 minus.n68 minus.n67 6.52702
R732 minus.n31 minus.n30 2.19141
R733 minus.n65 minus.n64 2.19141
R734 minus.n14 minus.n5 0.730803
R735 minus.n24 minus.n3 0.730803
R736 minus.n48 minus.n39 0.730803
R737 minus.n58 minus.n37 0.730803
R738 minus.n33 minus.n0 0.189894
R739 minus.n29 minus.n0 0.189894
R740 minus.n29 minus.n28 0.189894
R741 minus.n28 minus.n27 0.189894
R742 minus.n27 minus.n2 0.189894
R743 minus.n23 minus.n2 0.189894
R744 minus.n23 minus.n22 0.189894
R745 minus.n22 minus.n21 0.189894
R746 minus.n21 minus.n4 0.189894
R747 minus.n17 minus.n4 0.189894
R748 minus.n17 minus.n16 0.189894
R749 minus.n16 minus.n15 0.189894
R750 minus.n15 minus.n6 0.189894
R751 minus.n11 minus.n6 0.189894
R752 minus.n11 minus.n10 0.189894
R753 minus.n45 minus.n44 0.189894
R754 minus.n45 minus.n40 0.189894
R755 minus.n49 minus.n40 0.189894
R756 minus.n50 minus.n49 0.189894
R757 minus.n51 minus.n50 0.189894
R758 minus.n51 minus.n38 0.189894
R759 minus.n55 minus.n38 0.189894
R760 minus.n56 minus.n55 0.189894
R761 minus.n57 minus.n56 0.189894
R762 minus.n57 minus.n36 0.189894
R763 minus.n61 minus.n36 0.189894
R764 minus.n62 minus.n61 0.189894
R765 minus.n63 minus.n62 0.189894
R766 minus.n63 minus.n34 0.189894
R767 minus.n67 minus.n34 0.189894
R768 minus minus.n68 0.188
R769 drain_right.n7 drain_right.n5 67.9062
R770 drain_right.n2 drain_right.n0 67.9062
R771 drain_right.n13 drain_right.n11 67.9062
R772 drain_right.n13 drain_right.n12 67.1908
R773 drain_right.n15 drain_right.n14 67.1908
R774 drain_right.n17 drain_right.n16 67.1908
R775 drain_right.n19 drain_right.n18 67.1908
R776 drain_right.n21 drain_right.n20 67.1908
R777 drain_right.n7 drain_right.n6 67.1907
R778 drain_right.n9 drain_right.n8 67.1907
R779 drain_right.n4 drain_right.n3 67.1907
R780 drain_right.n2 drain_right.n1 67.1907
R781 drain_right drain_right.n10 29.0658
R782 drain_right drain_right.n21 6.36873
R783 drain_right.n5 drain_right.t22 3.3005
R784 drain_right.n5 drain_right.t7 3.3005
R785 drain_right.n6 drain_right.t8 3.3005
R786 drain_right.n6 drain_right.t13 3.3005
R787 drain_right.n8 drain_right.t17 3.3005
R788 drain_right.n8 drain_right.t0 3.3005
R789 drain_right.n3 drain_right.t2 3.3005
R790 drain_right.n3 drain_right.t16 3.3005
R791 drain_right.n1 drain_right.t20 3.3005
R792 drain_right.n1 drain_right.t21 3.3005
R793 drain_right.n0 drain_right.t4 3.3005
R794 drain_right.n0 drain_right.t5 3.3005
R795 drain_right.n11 drain_right.t19 3.3005
R796 drain_right.n11 drain_right.t10 3.3005
R797 drain_right.n12 drain_right.t3 3.3005
R798 drain_right.n12 drain_right.t14 3.3005
R799 drain_right.n14 drain_right.t12 3.3005
R800 drain_right.n14 drain_right.t15 3.3005
R801 drain_right.n16 drain_right.t11 3.3005
R802 drain_right.n16 drain_right.t23 3.3005
R803 drain_right.n18 drain_right.t18 3.3005
R804 drain_right.n18 drain_right.t6 3.3005
R805 drain_right.n20 drain_right.t1 3.3005
R806 drain_right.n20 drain_right.t9 3.3005
R807 drain_right.n9 drain_right.n7 0.716017
R808 drain_right.n4 drain_right.n2 0.716017
R809 drain_right.n21 drain_right.n19 0.716017
R810 drain_right.n19 drain_right.n17 0.716017
R811 drain_right.n17 drain_right.n15 0.716017
R812 drain_right.n15 drain_right.n13 0.716017
R813 drain_right.n10 drain_right.n9 0.302913
R814 drain_right.n10 drain_right.n4 0.302913
C0 drain_right drain_left 1.55979f
C1 minus drain_left 0.173624f
C2 drain_right minus 6.43784f
C3 source drain_left 19.1134f
C4 drain_right source 19.1149f
C5 minus source 6.83086f
C6 drain_left plus 6.72416f
C7 drain_right plus 0.443411f
C8 minus plus 5.63042f
C9 source plus 6.84488f
C10 drain_right a_n2874_n2088# 6.320179f
C11 drain_left a_n2874_n2088# 6.73654f
C12 source a_n2874_n2088# 5.765634f
C13 minus a_n2874_n2088# 10.999641f
C14 plus a_n2874_n2088# 12.63716f
C15 drain_right.t4 a_n2874_n2088# 0.138006f
C16 drain_right.t5 a_n2874_n2088# 0.138006f
C17 drain_right.n0 a_n2874_n2088# 1.155f
C18 drain_right.t20 a_n2874_n2088# 0.138006f
C19 drain_right.t21 a_n2874_n2088# 0.138006f
C20 drain_right.n1 a_n2874_n2088# 1.15097f
C21 drain_right.n2 a_n2874_n2088# 0.748604f
C22 drain_right.t2 a_n2874_n2088# 0.138006f
C23 drain_right.t16 a_n2874_n2088# 0.138006f
C24 drain_right.n3 a_n2874_n2088# 1.15097f
C25 drain_right.n4 a_n2874_n2088# 0.333941f
C26 drain_right.t22 a_n2874_n2088# 0.138006f
C27 drain_right.t7 a_n2874_n2088# 0.138006f
C28 drain_right.n5 a_n2874_n2088# 1.155f
C29 drain_right.t8 a_n2874_n2088# 0.138006f
C30 drain_right.t13 a_n2874_n2088# 0.138006f
C31 drain_right.n6 a_n2874_n2088# 1.15097f
C32 drain_right.n7 a_n2874_n2088# 0.748604f
C33 drain_right.t17 a_n2874_n2088# 0.138006f
C34 drain_right.t0 a_n2874_n2088# 0.138006f
C35 drain_right.n8 a_n2874_n2088# 1.15097f
C36 drain_right.n9 a_n2874_n2088# 0.333941f
C37 drain_right.n10 a_n2874_n2088# 1.30742f
C38 drain_right.t19 a_n2874_n2088# 0.138006f
C39 drain_right.t10 a_n2874_n2088# 0.138006f
C40 drain_right.n11 a_n2874_n2088# 1.155f
C41 drain_right.t3 a_n2874_n2088# 0.138006f
C42 drain_right.t14 a_n2874_n2088# 0.138006f
C43 drain_right.n12 a_n2874_n2088# 1.15097f
C44 drain_right.n13 a_n2874_n2088# 0.748599f
C45 drain_right.t12 a_n2874_n2088# 0.138006f
C46 drain_right.t15 a_n2874_n2088# 0.138006f
C47 drain_right.n14 a_n2874_n2088# 1.15097f
C48 drain_right.n15 a_n2874_n2088# 0.370448f
C49 drain_right.t11 a_n2874_n2088# 0.138006f
C50 drain_right.t23 a_n2874_n2088# 0.138006f
C51 drain_right.n16 a_n2874_n2088# 1.15097f
C52 drain_right.n17 a_n2874_n2088# 0.370448f
C53 drain_right.t18 a_n2874_n2088# 0.138006f
C54 drain_right.t6 a_n2874_n2088# 0.138006f
C55 drain_right.n18 a_n2874_n2088# 1.15097f
C56 drain_right.n19 a_n2874_n2088# 0.370448f
C57 drain_right.t1 a_n2874_n2088# 0.138006f
C58 drain_right.t9 a_n2874_n2088# 0.138006f
C59 drain_right.n20 a_n2874_n2088# 1.15097f
C60 drain_right.n21 a_n2874_n2088# 0.620515f
C61 minus.n0 a_n2874_n2088# 0.043616f
C62 minus.t5 a_n2874_n2088# 0.379533f
C63 minus.n1 a_n2874_n2088# 0.182951f
C64 minus.t14 a_n2874_n2088# 0.379533f
C65 minus.n2 a_n2874_n2088# 0.043616f
C66 minus.t12 a_n2874_n2088# 0.379533f
C67 minus.n3 a_n2874_n2088# 0.178917f
C68 minus.n4 a_n2874_n2088# 0.043616f
C69 minus.t8 a_n2874_n2088# 0.379533f
C70 minus.n5 a_n2874_n2088# 0.178917f
C71 minus.t11 a_n2874_n2088# 0.379533f
C72 minus.n6 a_n2874_n2088# 0.043616f
C73 minus.t9 a_n2874_n2088# 0.379533f
C74 minus.n7 a_n2874_n2088# 0.182951f
C75 minus.t13 a_n2874_n2088# 0.391486f
C76 minus.t4 a_n2874_n2088# 0.379533f
C77 minus.n8 a_n2874_n2088# 0.188112f
C78 minus.n9 a_n2874_n2088# 0.168259f
C79 minus.n10 a_n2874_n2088# 0.1771f
C80 minus.n11 a_n2874_n2088# 0.043616f
C81 minus.n12 a_n2874_n2088# 0.009897f
C82 minus.t20 a_n2874_n2088# 0.379533f
C83 minus.n13 a_n2874_n2088# 0.183354f
C84 minus.n14 a_n2874_n2088# 0.009897f
C85 minus.n15 a_n2874_n2088# 0.043616f
C86 minus.n16 a_n2874_n2088# 0.043616f
C87 minus.n17 a_n2874_n2088# 0.043616f
C88 minus.n18 a_n2874_n2088# 0.18322f
C89 minus.n19 a_n2874_n2088# 0.009897f
C90 minus.t0 a_n2874_n2088# 0.379533f
C91 minus.n20 a_n2874_n2088# 0.18322f
C92 minus.n21 a_n2874_n2088# 0.043616f
C93 minus.n22 a_n2874_n2088# 0.043616f
C94 minus.n23 a_n2874_n2088# 0.043616f
C95 minus.n24 a_n2874_n2088# 0.009897f
C96 minus.t17 a_n2874_n2088# 0.379533f
C97 minus.n25 a_n2874_n2088# 0.183354f
C98 minus.n26 a_n2874_n2088# 0.009897f
C99 minus.n27 a_n2874_n2088# 0.043616f
C100 minus.n28 a_n2874_n2088# 0.043616f
C101 minus.n29 a_n2874_n2088# 0.043616f
C102 minus.n30 a_n2874_n2088# 0.179186f
C103 minus.n31 a_n2874_n2088# 0.009897f
C104 minus.t22 a_n2874_n2088# 0.379533f
C105 minus.n32 a_n2874_n2088# 0.178379f
C106 minus.n33 a_n2874_n2088# 1.49551f
C107 minus.n34 a_n2874_n2088# 0.043616f
C108 minus.t10 a_n2874_n2088# 0.379533f
C109 minus.n35 a_n2874_n2088# 0.182951f
C110 minus.n36 a_n2874_n2088# 0.043616f
C111 minus.t23 a_n2874_n2088# 0.379533f
C112 minus.n37 a_n2874_n2088# 0.178917f
C113 minus.n38 a_n2874_n2088# 0.043616f
C114 minus.t21 a_n2874_n2088# 0.379533f
C115 minus.n39 a_n2874_n2088# 0.178917f
C116 minus.n40 a_n2874_n2088# 0.043616f
C117 minus.t3 a_n2874_n2088# 0.379533f
C118 minus.n41 a_n2874_n2088# 0.182951f
C119 minus.t19 a_n2874_n2088# 0.391486f
C120 minus.t18 a_n2874_n2088# 0.379533f
C121 minus.n42 a_n2874_n2088# 0.188112f
C122 minus.n43 a_n2874_n2088# 0.168259f
C123 minus.n44 a_n2874_n2088# 0.1771f
C124 minus.n45 a_n2874_n2088# 0.043616f
C125 minus.n46 a_n2874_n2088# 0.009897f
C126 minus.t2 a_n2874_n2088# 0.379533f
C127 minus.n47 a_n2874_n2088# 0.183354f
C128 minus.n48 a_n2874_n2088# 0.009897f
C129 minus.n49 a_n2874_n2088# 0.043616f
C130 minus.n50 a_n2874_n2088# 0.043616f
C131 minus.n51 a_n2874_n2088# 0.043616f
C132 minus.t7 a_n2874_n2088# 0.379533f
C133 minus.n52 a_n2874_n2088# 0.18322f
C134 minus.n53 a_n2874_n2088# 0.009897f
C135 minus.t6 a_n2874_n2088# 0.379533f
C136 minus.n54 a_n2874_n2088# 0.18322f
C137 minus.n55 a_n2874_n2088# 0.043616f
C138 minus.n56 a_n2874_n2088# 0.043616f
C139 minus.n57 a_n2874_n2088# 0.043616f
C140 minus.n58 a_n2874_n2088# 0.009897f
C141 minus.t15 a_n2874_n2088# 0.379533f
C142 minus.n59 a_n2874_n2088# 0.183354f
C143 minus.n60 a_n2874_n2088# 0.009897f
C144 minus.n61 a_n2874_n2088# 0.043616f
C145 minus.n62 a_n2874_n2088# 0.043616f
C146 minus.n63 a_n2874_n2088# 0.043616f
C147 minus.t1 a_n2874_n2088# 0.379533f
C148 minus.n64 a_n2874_n2088# 0.179186f
C149 minus.n65 a_n2874_n2088# 0.009897f
C150 minus.t16 a_n2874_n2088# 0.379533f
C151 minus.n66 a_n2874_n2088# 0.178379f
C152 minus.n67 a_n2874_n2088# 0.287924f
C153 minus.n68 a_n2874_n2088# 1.81936f
C154 drain_left.t15 a_n2874_n2088# 0.139009f
C155 drain_left.t6 a_n2874_n2088# 0.139009f
C156 drain_left.n0 a_n2874_n2088# 1.16339f
C157 drain_left.t22 a_n2874_n2088# 0.139009f
C158 drain_left.t23 a_n2874_n2088# 0.139009f
C159 drain_left.n1 a_n2874_n2088# 1.15933f
C160 drain_left.n2 a_n2874_n2088# 0.754044f
C161 drain_left.t11 a_n2874_n2088# 0.139009f
C162 drain_left.t4 a_n2874_n2088# 0.139009f
C163 drain_left.n3 a_n2874_n2088# 1.15933f
C164 drain_left.n4 a_n2874_n2088# 0.336368f
C165 drain_left.t12 a_n2874_n2088# 0.139009f
C166 drain_left.t13 a_n2874_n2088# 0.139009f
C167 drain_left.n5 a_n2874_n2088# 1.16339f
C168 drain_left.t9 a_n2874_n2088# 0.139009f
C169 drain_left.t1 a_n2874_n2088# 0.139009f
C170 drain_left.n6 a_n2874_n2088# 1.15933f
C171 drain_left.n7 a_n2874_n2088# 0.754044f
C172 drain_left.t21 a_n2874_n2088# 0.139009f
C173 drain_left.t8 a_n2874_n2088# 0.139009f
C174 drain_left.n8 a_n2874_n2088# 1.15933f
C175 drain_left.n9 a_n2874_n2088# 0.336368f
C176 drain_left.n10 a_n2874_n2088# 1.37551f
C177 drain_left.t17 a_n2874_n2088# 0.139009f
C178 drain_left.t7 a_n2874_n2088# 0.139009f
C179 drain_left.n11 a_n2874_n2088# 1.16339f
C180 drain_left.t2 a_n2874_n2088# 0.139009f
C181 drain_left.t16 a_n2874_n2088# 0.139009f
C182 drain_left.n12 a_n2874_n2088# 1.15934f
C183 drain_left.n13 a_n2874_n2088# 0.754033f
C184 drain_left.t5 a_n2874_n2088# 0.139009f
C185 drain_left.t0 a_n2874_n2088# 0.139009f
C186 drain_left.n14 a_n2874_n2088# 1.15934f
C187 drain_left.n15 a_n2874_n2088# 0.373141f
C188 drain_left.t14 a_n2874_n2088# 0.139009f
C189 drain_left.t3 a_n2874_n2088# 0.139009f
C190 drain_left.n16 a_n2874_n2088# 1.15934f
C191 drain_left.n17 a_n2874_n2088# 0.373141f
C192 drain_left.t18 a_n2874_n2088# 0.139009f
C193 drain_left.t10 a_n2874_n2088# 0.139009f
C194 drain_left.n18 a_n2874_n2088# 1.15934f
C195 drain_left.n19 a_n2874_n2088# 0.373141f
C196 drain_left.t19 a_n2874_n2088# 0.139009f
C197 drain_left.t20 a_n2874_n2088# 0.139009f
C198 drain_left.n20 a_n2874_n2088# 1.15933f
C199 drain_left.n21 a_n2874_n2088# 0.62503f
C200 source.n0 a_n2874_n2088# 0.039382f
C201 source.n1 a_n2874_n2088# 0.028018f
C202 source.n2 a_n2874_n2088# 0.015056f
C203 source.n3 a_n2874_n2088# 0.035586f
C204 source.n4 a_n2874_n2088# 0.015941f
C205 source.n5 a_n2874_n2088# 0.028018f
C206 source.n6 a_n2874_n2088# 0.015056f
C207 source.n7 a_n2874_n2088# 0.035586f
C208 source.n8 a_n2874_n2088# 0.015941f
C209 source.n9 a_n2874_n2088# 0.119897f
C210 source.t39 a_n2874_n2088# 0.058001f
C211 source.n10 a_n2874_n2088# 0.026689f
C212 source.n11 a_n2874_n2088# 0.02102f
C213 source.n12 a_n2874_n2088# 0.015056f
C214 source.n13 a_n2874_n2088# 0.666658f
C215 source.n14 a_n2874_n2088# 0.028018f
C216 source.n15 a_n2874_n2088# 0.015056f
C217 source.n16 a_n2874_n2088# 0.015941f
C218 source.n17 a_n2874_n2088# 0.035586f
C219 source.n18 a_n2874_n2088# 0.035586f
C220 source.n19 a_n2874_n2088# 0.015941f
C221 source.n20 a_n2874_n2088# 0.015056f
C222 source.n21 a_n2874_n2088# 0.028018f
C223 source.n22 a_n2874_n2088# 0.028018f
C224 source.n23 a_n2874_n2088# 0.015056f
C225 source.n24 a_n2874_n2088# 0.015941f
C226 source.n25 a_n2874_n2088# 0.035586f
C227 source.n26 a_n2874_n2088# 0.077038f
C228 source.n27 a_n2874_n2088# 0.015941f
C229 source.n28 a_n2874_n2088# 0.015056f
C230 source.n29 a_n2874_n2088# 0.064762f
C231 source.n30 a_n2874_n2088# 0.043106f
C232 source.n31 a_n2874_n2088# 0.705312f
C233 source.t24 a_n2874_n2088# 0.132843f
C234 source.t42 a_n2874_n2088# 0.132843f
C235 source.n32 a_n2874_n2088# 1.0346f
C236 source.n33 a_n2874_n2088# 0.391834f
C237 source.t33 a_n2874_n2088# 0.132843f
C238 source.t22 a_n2874_n2088# 0.132843f
C239 source.n34 a_n2874_n2088# 1.0346f
C240 source.n35 a_n2874_n2088# 0.391834f
C241 source.t40 a_n2874_n2088# 0.132843f
C242 source.t34 a_n2874_n2088# 0.132843f
C243 source.n36 a_n2874_n2088# 1.0346f
C244 source.n37 a_n2874_n2088# 0.391834f
C245 source.t25 a_n2874_n2088# 0.132843f
C246 source.t31 a_n2874_n2088# 0.132843f
C247 source.n38 a_n2874_n2088# 1.0346f
C248 source.n39 a_n2874_n2088# 0.391834f
C249 source.t45 a_n2874_n2088# 0.132843f
C250 source.t27 a_n2874_n2088# 0.132843f
C251 source.n40 a_n2874_n2088# 1.0346f
C252 source.n41 a_n2874_n2088# 0.391834f
C253 source.n42 a_n2874_n2088# 0.039382f
C254 source.n43 a_n2874_n2088# 0.028018f
C255 source.n44 a_n2874_n2088# 0.015056f
C256 source.n45 a_n2874_n2088# 0.035586f
C257 source.n46 a_n2874_n2088# 0.015941f
C258 source.n47 a_n2874_n2088# 0.028018f
C259 source.n48 a_n2874_n2088# 0.015056f
C260 source.n49 a_n2874_n2088# 0.035586f
C261 source.n50 a_n2874_n2088# 0.015941f
C262 source.n51 a_n2874_n2088# 0.119897f
C263 source.t28 a_n2874_n2088# 0.058001f
C264 source.n52 a_n2874_n2088# 0.026689f
C265 source.n53 a_n2874_n2088# 0.02102f
C266 source.n54 a_n2874_n2088# 0.015056f
C267 source.n55 a_n2874_n2088# 0.666658f
C268 source.n56 a_n2874_n2088# 0.028018f
C269 source.n57 a_n2874_n2088# 0.015056f
C270 source.n58 a_n2874_n2088# 0.015941f
C271 source.n59 a_n2874_n2088# 0.035586f
C272 source.n60 a_n2874_n2088# 0.035586f
C273 source.n61 a_n2874_n2088# 0.015941f
C274 source.n62 a_n2874_n2088# 0.015056f
C275 source.n63 a_n2874_n2088# 0.028018f
C276 source.n64 a_n2874_n2088# 0.028018f
C277 source.n65 a_n2874_n2088# 0.015056f
C278 source.n66 a_n2874_n2088# 0.015941f
C279 source.n67 a_n2874_n2088# 0.035586f
C280 source.n68 a_n2874_n2088# 0.077038f
C281 source.n69 a_n2874_n2088# 0.015941f
C282 source.n70 a_n2874_n2088# 0.015056f
C283 source.n71 a_n2874_n2088# 0.064762f
C284 source.n72 a_n2874_n2088# 0.043106f
C285 source.n73 a_n2874_n2088# 0.130942f
C286 source.n74 a_n2874_n2088# 0.039382f
C287 source.n75 a_n2874_n2088# 0.028018f
C288 source.n76 a_n2874_n2088# 0.015056f
C289 source.n77 a_n2874_n2088# 0.035586f
C290 source.n78 a_n2874_n2088# 0.015941f
C291 source.n79 a_n2874_n2088# 0.028018f
C292 source.n80 a_n2874_n2088# 0.015056f
C293 source.n81 a_n2874_n2088# 0.035586f
C294 source.n82 a_n2874_n2088# 0.015941f
C295 source.n83 a_n2874_n2088# 0.119897f
C296 source.t21 a_n2874_n2088# 0.058001f
C297 source.n84 a_n2874_n2088# 0.026689f
C298 source.n85 a_n2874_n2088# 0.02102f
C299 source.n86 a_n2874_n2088# 0.015056f
C300 source.n87 a_n2874_n2088# 0.666658f
C301 source.n88 a_n2874_n2088# 0.028018f
C302 source.n89 a_n2874_n2088# 0.015056f
C303 source.n90 a_n2874_n2088# 0.015941f
C304 source.n91 a_n2874_n2088# 0.035586f
C305 source.n92 a_n2874_n2088# 0.035586f
C306 source.n93 a_n2874_n2088# 0.015941f
C307 source.n94 a_n2874_n2088# 0.015056f
C308 source.n95 a_n2874_n2088# 0.028018f
C309 source.n96 a_n2874_n2088# 0.028018f
C310 source.n97 a_n2874_n2088# 0.015056f
C311 source.n98 a_n2874_n2088# 0.015941f
C312 source.n99 a_n2874_n2088# 0.035586f
C313 source.n100 a_n2874_n2088# 0.077038f
C314 source.n101 a_n2874_n2088# 0.015941f
C315 source.n102 a_n2874_n2088# 0.015056f
C316 source.n103 a_n2874_n2088# 0.064762f
C317 source.n104 a_n2874_n2088# 0.043106f
C318 source.n105 a_n2874_n2088# 0.130942f
C319 source.t46 a_n2874_n2088# 0.132843f
C320 source.t7 a_n2874_n2088# 0.132843f
C321 source.n106 a_n2874_n2088# 1.0346f
C322 source.n107 a_n2874_n2088# 0.391834f
C323 source.t12 a_n2874_n2088# 0.132843f
C324 source.t10 a_n2874_n2088# 0.132843f
C325 source.n108 a_n2874_n2088# 1.0346f
C326 source.n109 a_n2874_n2088# 0.391834f
C327 source.t19 a_n2874_n2088# 0.132843f
C328 source.t6 a_n2874_n2088# 0.132843f
C329 source.n110 a_n2874_n2088# 1.0346f
C330 source.n111 a_n2874_n2088# 0.391834f
C331 source.t14 a_n2874_n2088# 0.132843f
C332 source.t0 a_n2874_n2088# 0.132843f
C333 source.n112 a_n2874_n2088# 1.0346f
C334 source.n113 a_n2874_n2088# 0.391834f
C335 source.t15 a_n2874_n2088# 0.132843f
C336 source.t5 a_n2874_n2088# 0.132843f
C337 source.n114 a_n2874_n2088# 1.0346f
C338 source.n115 a_n2874_n2088# 0.391834f
C339 source.n116 a_n2874_n2088# 0.039382f
C340 source.n117 a_n2874_n2088# 0.028018f
C341 source.n118 a_n2874_n2088# 0.015056f
C342 source.n119 a_n2874_n2088# 0.035586f
C343 source.n120 a_n2874_n2088# 0.015941f
C344 source.n121 a_n2874_n2088# 0.028018f
C345 source.n122 a_n2874_n2088# 0.015056f
C346 source.n123 a_n2874_n2088# 0.035586f
C347 source.n124 a_n2874_n2088# 0.015941f
C348 source.n125 a_n2874_n2088# 0.119897f
C349 source.t2 a_n2874_n2088# 0.058001f
C350 source.n126 a_n2874_n2088# 0.026689f
C351 source.n127 a_n2874_n2088# 0.02102f
C352 source.n128 a_n2874_n2088# 0.015056f
C353 source.n129 a_n2874_n2088# 0.666658f
C354 source.n130 a_n2874_n2088# 0.028018f
C355 source.n131 a_n2874_n2088# 0.015056f
C356 source.n132 a_n2874_n2088# 0.015941f
C357 source.n133 a_n2874_n2088# 0.035586f
C358 source.n134 a_n2874_n2088# 0.035586f
C359 source.n135 a_n2874_n2088# 0.015941f
C360 source.n136 a_n2874_n2088# 0.015056f
C361 source.n137 a_n2874_n2088# 0.028018f
C362 source.n138 a_n2874_n2088# 0.028018f
C363 source.n139 a_n2874_n2088# 0.015056f
C364 source.n140 a_n2874_n2088# 0.015941f
C365 source.n141 a_n2874_n2088# 0.035586f
C366 source.n142 a_n2874_n2088# 0.077038f
C367 source.n143 a_n2874_n2088# 0.015941f
C368 source.n144 a_n2874_n2088# 0.015056f
C369 source.n145 a_n2874_n2088# 0.064762f
C370 source.n146 a_n2874_n2088# 0.043106f
C371 source.n147 a_n2874_n2088# 1.07048f
C372 source.n148 a_n2874_n2088# 0.039382f
C373 source.n149 a_n2874_n2088# 0.028018f
C374 source.n150 a_n2874_n2088# 0.015056f
C375 source.n151 a_n2874_n2088# 0.035586f
C376 source.n152 a_n2874_n2088# 0.015941f
C377 source.n153 a_n2874_n2088# 0.028018f
C378 source.n154 a_n2874_n2088# 0.015056f
C379 source.n155 a_n2874_n2088# 0.035586f
C380 source.n156 a_n2874_n2088# 0.015941f
C381 source.n157 a_n2874_n2088# 0.119897f
C382 source.t44 a_n2874_n2088# 0.058001f
C383 source.n158 a_n2874_n2088# 0.026689f
C384 source.n159 a_n2874_n2088# 0.02102f
C385 source.n160 a_n2874_n2088# 0.015056f
C386 source.n161 a_n2874_n2088# 0.666658f
C387 source.n162 a_n2874_n2088# 0.028018f
C388 source.n163 a_n2874_n2088# 0.015056f
C389 source.n164 a_n2874_n2088# 0.015941f
C390 source.n165 a_n2874_n2088# 0.035586f
C391 source.n166 a_n2874_n2088# 0.035586f
C392 source.n167 a_n2874_n2088# 0.015941f
C393 source.n168 a_n2874_n2088# 0.015056f
C394 source.n169 a_n2874_n2088# 0.028018f
C395 source.n170 a_n2874_n2088# 0.028018f
C396 source.n171 a_n2874_n2088# 0.015056f
C397 source.n172 a_n2874_n2088# 0.015941f
C398 source.n173 a_n2874_n2088# 0.035586f
C399 source.n174 a_n2874_n2088# 0.077038f
C400 source.n175 a_n2874_n2088# 0.015941f
C401 source.n176 a_n2874_n2088# 0.015056f
C402 source.n177 a_n2874_n2088# 0.064762f
C403 source.n178 a_n2874_n2088# 0.043106f
C404 source.n179 a_n2874_n2088# 1.07048f
C405 source.t26 a_n2874_n2088# 0.132843f
C406 source.t43 a_n2874_n2088# 0.132843f
C407 source.n180 a_n2874_n2088# 1.03459f
C408 source.n181 a_n2874_n2088# 0.391842f
C409 source.t41 a_n2874_n2088# 0.132843f
C410 source.t36 a_n2874_n2088# 0.132843f
C411 source.n182 a_n2874_n2088# 1.03459f
C412 source.n183 a_n2874_n2088# 0.391842f
C413 source.t32 a_n2874_n2088# 0.132843f
C414 source.t38 a_n2874_n2088# 0.132843f
C415 source.n184 a_n2874_n2088# 1.03459f
C416 source.n185 a_n2874_n2088# 0.391842f
C417 source.t30 a_n2874_n2088# 0.132843f
C418 source.t37 a_n2874_n2088# 0.132843f
C419 source.n186 a_n2874_n2088# 1.03459f
C420 source.n187 a_n2874_n2088# 0.391842f
C421 source.t35 a_n2874_n2088# 0.132843f
C422 source.t29 a_n2874_n2088# 0.132843f
C423 source.n188 a_n2874_n2088# 1.03459f
C424 source.n189 a_n2874_n2088# 0.391842f
C425 source.n190 a_n2874_n2088# 0.039382f
C426 source.n191 a_n2874_n2088# 0.028018f
C427 source.n192 a_n2874_n2088# 0.015056f
C428 source.n193 a_n2874_n2088# 0.035586f
C429 source.n194 a_n2874_n2088# 0.015941f
C430 source.n195 a_n2874_n2088# 0.028018f
C431 source.n196 a_n2874_n2088# 0.015056f
C432 source.n197 a_n2874_n2088# 0.035586f
C433 source.n198 a_n2874_n2088# 0.015941f
C434 source.n199 a_n2874_n2088# 0.119897f
C435 source.t23 a_n2874_n2088# 0.058001f
C436 source.n200 a_n2874_n2088# 0.026689f
C437 source.n201 a_n2874_n2088# 0.02102f
C438 source.n202 a_n2874_n2088# 0.015056f
C439 source.n203 a_n2874_n2088# 0.666658f
C440 source.n204 a_n2874_n2088# 0.028018f
C441 source.n205 a_n2874_n2088# 0.015056f
C442 source.n206 a_n2874_n2088# 0.015941f
C443 source.n207 a_n2874_n2088# 0.035586f
C444 source.n208 a_n2874_n2088# 0.035586f
C445 source.n209 a_n2874_n2088# 0.015941f
C446 source.n210 a_n2874_n2088# 0.015056f
C447 source.n211 a_n2874_n2088# 0.028018f
C448 source.n212 a_n2874_n2088# 0.028018f
C449 source.n213 a_n2874_n2088# 0.015056f
C450 source.n214 a_n2874_n2088# 0.015941f
C451 source.n215 a_n2874_n2088# 0.035586f
C452 source.n216 a_n2874_n2088# 0.077038f
C453 source.n217 a_n2874_n2088# 0.015941f
C454 source.n218 a_n2874_n2088# 0.015056f
C455 source.n219 a_n2874_n2088# 0.064762f
C456 source.n220 a_n2874_n2088# 0.043106f
C457 source.n221 a_n2874_n2088# 0.130942f
C458 source.n222 a_n2874_n2088# 0.039382f
C459 source.n223 a_n2874_n2088# 0.028018f
C460 source.n224 a_n2874_n2088# 0.015056f
C461 source.n225 a_n2874_n2088# 0.035586f
C462 source.n226 a_n2874_n2088# 0.015941f
C463 source.n227 a_n2874_n2088# 0.028018f
C464 source.n228 a_n2874_n2088# 0.015056f
C465 source.n229 a_n2874_n2088# 0.035586f
C466 source.n230 a_n2874_n2088# 0.015941f
C467 source.n231 a_n2874_n2088# 0.119897f
C468 source.t8 a_n2874_n2088# 0.058001f
C469 source.n232 a_n2874_n2088# 0.026689f
C470 source.n233 a_n2874_n2088# 0.02102f
C471 source.n234 a_n2874_n2088# 0.015056f
C472 source.n235 a_n2874_n2088# 0.666658f
C473 source.n236 a_n2874_n2088# 0.028018f
C474 source.n237 a_n2874_n2088# 0.015056f
C475 source.n238 a_n2874_n2088# 0.015941f
C476 source.n239 a_n2874_n2088# 0.035586f
C477 source.n240 a_n2874_n2088# 0.035586f
C478 source.n241 a_n2874_n2088# 0.015941f
C479 source.n242 a_n2874_n2088# 0.015056f
C480 source.n243 a_n2874_n2088# 0.028018f
C481 source.n244 a_n2874_n2088# 0.028018f
C482 source.n245 a_n2874_n2088# 0.015056f
C483 source.n246 a_n2874_n2088# 0.015941f
C484 source.n247 a_n2874_n2088# 0.035586f
C485 source.n248 a_n2874_n2088# 0.077038f
C486 source.n249 a_n2874_n2088# 0.015941f
C487 source.n250 a_n2874_n2088# 0.015056f
C488 source.n251 a_n2874_n2088# 0.064762f
C489 source.n252 a_n2874_n2088# 0.043106f
C490 source.n253 a_n2874_n2088# 0.130942f
C491 source.t17 a_n2874_n2088# 0.132843f
C492 source.t3 a_n2874_n2088# 0.132843f
C493 source.n254 a_n2874_n2088# 1.03459f
C494 source.n255 a_n2874_n2088# 0.391842f
C495 source.t11 a_n2874_n2088# 0.132843f
C496 source.t1 a_n2874_n2088# 0.132843f
C497 source.n256 a_n2874_n2088# 1.03459f
C498 source.n257 a_n2874_n2088# 0.391842f
C499 source.t13 a_n2874_n2088# 0.132843f
C500 source.t20 a_n2874_n2088# 0.132843f
C501 source.n258 a_n2874_n2088# 1.03459f
C502 source.n259 a_n2874_n2088# 0.391842f
C503 source.t16 a_n2874_n2088# 0.132843f
C504 source.t18 a_n2874_n2088# 0.132843f
C505 source.n260 a_n2874_n2088# 1.03459f
C506 source.n261 a_n2874_n2088# 0.391842f
C507 source.t47 a_n2874_n2088# 0.132843f
C508 source.t4 a_n2874_n2088# 0.132843f
C509 source.n262 a_n2874_n2088# 1.03459f
C510 source.n263 a_n2874_n2088# 0.391842f
C511 source.n264 a_n2874_n2088# 0.039382f
C512 source.n265 a_n2874_n2088# 0.028018f
C513 source.n266 a_n2874_n2088# 0.015056f
C514 source.n267 a_n2874_n2088# 0.035586f
C515 source.n268 a_n2874_n2088# 0.015941f
C516 source.n269 a_n2874_n2088# 0.028018f
C517 source.n270 a_n2874_n2088# 0.015056f
C518 source.n271 a_n2874_n2088# 0.035586f
C519 source.n272 a_n2874_n2088# 0.015941f
C520 source.n273 a_n2874_n2088# 0.119897f
C521 source.t9 a_n2874_n2088# 0.058001f
C522 source.n274 a_n2874_n2088# 0.026689f
C523 source.n275 a_n2874_n2088# 0.02102f
C524 source.n276 a_n2874_n2088# 0.015056f
C525 source.n277 a_n2874_n2088# 0.666658f
C526 source.n278 a_n2874_n2088# 0.028018f
C527 source.n279 a_n2874_n2088# 0.015056f
C528 source.n280 a_n2874_n2088# 0.015941f
C529 source.n281 a_n2874_n2088# 0.035586f
C530 source.n282 a_n2874_n2088# 0.035586f
C531 source.n283 a_n2874_n2088# 0.015941f
C532 source.n284 a_n2874_n2088# 0.015056f
C533 source.n285 a_n2874_n2088# 0.028018f
C534 source.n286 a_n2874_n2088# 0.028018f
C535 source.n287 a_n2874_n2088# 0.015056f
C536 source.n288 a_n2874_n2088# 0.015941f
C537 source.n289 a_n2874_n2088# 0.035586f
C538 source.n290 a_n2874_n2088# 0.077038f
C539 source.n291 a_n2874_n2088# 0.015941f
C540 source.n292 a_n2874_n2088# 0.015056f
C541 source.n293 a_n2874_n2088# 0.064762f
C542 source.n294 a_n2874_n2088# 0.043106f
C543 source.n295 a_n2874_n2088# 0.301473f
C544 source.n296 a_n2874_n2088# 1.15411f
C545 plus.n0 a_n2874_n2088# 0.044521f
C546 plus.t3 a_n2874_n2088# 0.387407f
C547 plus.t4 a_n2874_n2088# 0.387407f
C548 plus.n1 a_n2874_n2088# 0.044521f
C549 plus.t13 a_n2874_n2088# 0.387407f
C550 plus.n2 a_n2874_n2088# 0.044521f
C551 plus.t5 a_n2874_n2088# 0.387407f
C552 plus.n3 a_n2874_n2088# 0.187158f
C553 plus.n4 a_n2874_n2088# 0.044521f
C554 plus.t20 a_n2874_n2088# 0.387407f
C555 plus.t9 a_n2874_n2088# 0.387407f
C556 plus.n5 a_n2874_n2088# 0.044521f
C557 plus.t23 a_n2874_n2088# 0.387407f
C558 plus.n6 a_n2874_n2088# 0.187021f
C559 plus.n7 a_n2874_n2088# 0.044521f
C560 plus.t18 a_n2874_n2088# 0.387407f
C561 plus.t7 a_n2874_n2088# 0.387407f
C562 plus.n8 a_n2874_n2088# 0.044521f
C563 plus.t21 a_n2874_n2088# 0.387407f
C564 plus.n9 a_n2874_n2088# 0.186746f
C565 plus.t16 a_n2874_n2088# 0.387407f
C566 plus.n10 a_n2874_n2088# 0.192014f
C567 plus.t6 a_n2874_n2088# 0.399608f
C568 plus.n11 a_n2874_n2088# 0.17175f
C569 plus.n12 a_n2874_n2088# 0.180774f
C570 plus.n13 a_n2874_n2088# 0.044521f
C571 plus.n14 a_n2874_n2088# 0.010103f
C572 plus.n15 a_n2874_n2088# 0.187158f
C573 plus.n16 a_n2874_n2088# 0.010103f
C574 plus.n17 a_n2874_n2088# 0.182629f
C575 plus.n18 a_n2874_n2088# 0.044521f
C576 plus.n19 a_n2874_n2088# 0.044521f
C577 plus.n20 a_n2874_n2088# 0.044521f
C578 plus.n21 a_n2874_n2088# 0.010103f
C579 plus.n22 a_n2874_n2088# 0.187021f
C580 plus.n23 a_n2874_n2088# 0.182629f
C581 plus.n24 a_n2874_n2088# 0.010103f
C582 plus.n25 a_n2874_n2088# 0.044521f
C583 plus.n26 a_n2874_n2088# 0.044521f
C584 plus.n27 a_n2874_n2088# 0.044521f
C585 plus.n28 a_n2874_n2088# 0.010103f
C586 plus.n29 a_n2874_n2088# 0.186746f
C587 plus.n30 a_n2874_n2088# 0.182903f
C588 plus.n31 a_n2874_n2088# 0.010103f
C589 plus.n32 a_n2874_n2088# 0.18208f
C590 plus.n33 a_n2874_n2088# 0.384451f
C591 plus.n34 a_n2874_n2088# 0.044521f
C592 plus.t8 a_n2874_n2088# 0.387407f
C593 plus.n35 a_n2874_n2088# 0.044521f
C594 plus.t17 a_n2874_n2088# 0.387407f
C595 plus.n36 a_n2874_n2088# 0.044521f
C596 plus.t1 a_n2874_n2088# 0.387407f
C597 plus.t0 a_n2874_n2088# 0.387407f
C598 plus.n37 a_n2874_n2088# 0.187158f
C599 plus.n38 a_n2874_n2088# 0.044521f
C600 plus.t12 a_n2874_n2088# 0.387407f
C601 plus.n39 a_n2874_n2088# 0.044521f
C602 plus.t19 a_n2874_n2088# 0.387407f
C603 plus.t2 a_n2874_n2088# 0.387407f
C604 plus.n40 a_n2874_n2088# 0.187021f
C605 plus.n41 a_n2874_n2088# 0.044521f
C606 plus.t15 a_n2874_n2088# 0.387407f
C607 plus.n42 a_n2874_n2088# 0.044521f
C608 plus.t14 a_n2874_n2088# 0.387407f
C609 plus.t22 a_n2874_n2088# 0.387407f
C610 plus.n43 a_n2874_n2088# 0.186746f
C611 plus.t10 a_n2874_n2088# 0.399608f
C612 plus.t11 a_n2874_n2088# 0.387407f
C613 plus.n44 a_n2874_n2088# 0.192014f
C614 plus.n45 a_n2874_n2088# 0.17175f
C615 plus.n46 a_n2874_n2088# 0.180774f
C616 plus.n47 a_n2874_n2088# 0.044521f
C617 plus.n48 a_n2874_n2088# 0.010103f
C618 plus.n49 a_n2874_n2088# 0.187158f
C619 plus.n50 a_n2874_n2088# 0.010103f
C620 plus.n51 a_n2874_n2088# 0.182629f
C621 plus.n52 a_n2874_n2088# 0.044521f
C622 plus.n53 a_n2874_n2088# 0.044521f
C623 plus.n54 a_n2874_n2088# 0.044521f
C624 plus.n55 a_n2874_n2088# 0.010103f
C625 plus.n56 a_n2874_n2088# 0.187021f
C626 plus.n57 a_n2874_n2088# 0.182629f
C627 plus.n58 a_n2874_n2088# 0.010103f
C628 plus.n59 a_n2874_n2088# 0.044521f
C629 plus.n60 a_n2874_n2088# 0.044521f
C630 plus.n61 a_n2874_n2088# 0.044521f
C631 plus.n62 a_n2874_n2088# 0.010103f
C632 plus.n63 a_n2874_n2088# 0.186746f
C633 plus.n64 a_n2874_n2088# 0.182903f
C634 plus.n65 a_n2874_n2088# 0.010103f
C635 plus.n66 a_n2874_n2088# 0.18208f
C636 plus.n67 a_n2874_n2088# 1.38273f
.ends

