* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 CSoutput.t109 commonsourceibias.t48 gnd.t304 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 vdd.t175 a_n5644_8799.t36 CSoutput.t113 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n1986_8322.t11 a_n2848_n452.t48 vdd.t94 vdd.t93 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n1808_13878.t19 a_n2848_n452.t37 a_n2848_n452.t38 vdd.t110 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X4 CSoutput.t108 commonsourceibias.t49 gnd.t303 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 a_n5644_8799.t24 plus.t5 a_n3106_n452.t25 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X6 gnd.t302 commonsourceibias.t50 CSoutput.t107 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t106 commonsourceibias.t51 gnd.t301 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 a_n3106_n452.t24 plus.t6 a_n5644_8799.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X9 a_n2848_n452.t26 a_n2848_n452.t25 a_n1808_13878.t18 vdd.t111 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 a_n1808_13878.t17 a_n2848_n452.t39 a_n2848_n452.t40 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 vdd.t89 vdd.t87 vdd.t88 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X12 a_n1808_13878.t7 a_n2848_n452.t49 vdd.t96 vdd.t95 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 output.t3 outputibias.t8 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X14 CSoutput.t31 a_n5644_8799.t37 vdd.t174 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 vdd.t86 vdd.t84 vdd.t85 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X16 gnd.t300 commonsourceibias.t52 CSoutput.t105 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X17 CSoutput.t104 commonsourceibias.t53 gnd.t299 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 gnd.t298 commonsourceibias.t54 CSoutput.t103 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t102 commonsourceibias.t55 gnd.t297 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 gnd.t183 gnd.t180 gnd.t182 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X21 CSoutput.t101 commonsourceibias.t56 gnd.t296 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 a_n1986_8322.t23 a_n2848_n452.t50 a_n5644_8799.t18 vdd.t109 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X23 CSoutput.t100 commonsourceibias.t57 gnd.t295 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 a_n2848_n452.t45 minus.t5 a_n3106_n452.t49 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X25 a_n5644_8799.t29 plus.t7 a_n3106_n452.t23 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 plus.t4 gnd.t177 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 a_n2848_n452.t8 minus.t6 a_n3106_n452.t34 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 gnd.t294 commonsourceibias.t58 CSoutput.t99 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 CSoutput.t98 commonsourceibias.t59 gnd.t293 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 CSoutput.t97 commonsourceibias.t60 gnd.t292 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 gnd.t176 gnd.t174 gnd.t175 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X32 CSoutput.t120 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X33 CSoutput.t16 a_n5644_8799.t38 vdd.t173 vdd.t131 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X34 vdd.t172 a_n5644_8799.t39 CSoutput.t37 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n3106_n452.t22 plus.t8 a_n5644_8799.t26 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X36 CSoutput.t96 commonsourceibias.t61 gnd.t277 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 a_n5644_8799.t19 a_n2848_n452.t51 a_n1986_8322.t22 vdd.t110 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X38 CSoutput.t33 a_n5644_8799.t40 vdd.t171 vdd.t112 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X39 vdd.t170 a_n5644_8799.t41 CSoutput.t4 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X40 a_n3106_n452.t42 minus.t7 a_n2848_n452.t14 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X41 gnd.t278 commonsourceibias.t62 CSoutput.t95 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 a_n3106_n452.t55 diffpairibias.t16 gnd.t325 gnd.t324 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 CSoutput.t94 commonsourceibias.t63 gnd.t291 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X44 gnd.t290 commonsourceibias.t0 commonsourceibias.t1 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 gnd.t173 gnd.t170 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X46 output.t19 CSoutput.t121 vdd.t177 gnd.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X47 CSoutput.t93 commonsourceibias.t64 gnd.t289 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 CSoutput.t10 a_n5644_8799.t42 vdd.t169 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 vdd.t83 vdd.t81 vdd.t82 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X50 CSoutput.t92 commonsourceibias.t65 gnd.t288 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 gnd.t169 gnd.t167 gnd.t168 gnd.t102 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X52 outputibias.t7 outputibias.t6 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X53 gnd.t287 commonsourceibias.t66 CSoutput.t91 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 output.t18 CSoutput.t122 vdd.t190 gnd.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X55 CSoutput.t90 commonsourceibias.t67 gnd.t286 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 a_n3106_n452.t21 plus.t9 a_n5644_8799.t16 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X57 gnd.t166 gnd.t164 gnd.t165 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X58 CSoutput.t89 commonsourceibias.t68 gnd.t285 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 gnd.t284 commonsourceibias.t40 commonsourceibias.t41 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 gnd.t163 gnd.t161 gnd.t162 gnd.t78 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X61 a_n1808_13878.t16 a_n2848_n452.t27 a_n2848_n452.t28 vdd.t100 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X62 vdd.t168 a_n5644_8799.t43 CSoutput.t9 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 a_n3106_n452.t20 plus.t10 a_n5644_8799.t21 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X64 a_n3106_n452.t48 minus.t8 a_n2848_n452.t44 gnd.t305 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X65 diffpairibias.t15 diffpairibias.t14 gnd.t307 gnd.t306 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X66 a_n2848_n452.t18 a_n2848_n452.t17 a_n1808_13878.t15 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X67 CSoutput.t14 a_n5644_8799.t44 vdd.t167 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 CSoutput.t88 commonsourceibias.t69 gnd.t283 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X69 CSoutput.t87 commonsourceibias.t70 gnd.t282 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X70 vdd.t80 vdd.t78 vdd.t79 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X71 gnd.t281 commonsourceibias.t71 CSoutput.t86 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 gnd.t280 commonsourceibias.t72 CSoutput.t85 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 CSoutput.t84 commonsourceibias.t73 gnd.t279 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X74 diffpairibias.t13 diffpairibias.t12 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X75 gnd.t276 commonsourceibias.t38 commonsourceibias.t39 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 vdd.t77 vdd.t75 vdd.t76 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X77 CSoutput.t83 commonsourceibias.t74 gnd.t275 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 gnd.t256 commonsourceibias.t75 CSoutput.t82 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 CSoutput.t81 commonsourceibias.t76 gnd.t274 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 vdd.t166 a_n5644_8799.t45 CSoutput.t0 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 gnd.t273 commonsourceibias.t77 CSoutput.t80 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 output.t17 CSoutput.t123 vdd.t179 gnd.t57 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X83 vdd.t164 a_n5644_8799.t46 CSoutput.t119 vdd.t140 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 CSoutput.t5 a_n5644_8799.t47 vdd.t163 vdd.t112 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X85 a_n3106_n452.t29 minus.t9 a_n2848_n452.t4 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X86 a_n3106_n452.t19 plus.t11 a_n5644_8799.t31 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X87 vdd.t162 a_n5644_8799.t48 CSoutput.t7 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 a_n5644_8799.t28 plus.t12 a_n3106_n452.t18 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X89 gnd.t272 commonsourceibias.t78 CSoutput.t79 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 gnd.t160 gnd.t157 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X91 CSoutput.t13 a_n5644_8799.t49 vdd.t161 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 CSoutput.t1 a_n5644_8799.t50 vdd.t160 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 vdd.t180 CSoutput.t124 output.t16 gnd.t58 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X94 a_n3106_n452.t0 diffpairibias.t17 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X95 CSoutput.t28 a_n5644_8799.t51 vdd.t159 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 a_n3106_n452.t17 plus.t13 a_n5644_8799.t30 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X97 gnd.t271 commonsourceibias.t79 CSoutput.t78 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 gnd.t156 gnd.t154 gnd.t155 gnd.t82 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X99 vdd.t158 a_n5644_8799.t52 CSoutput.t18 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 gnd.t153 gnd.t151 gnd.t152 gnd.t82 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X101 a_n2848_n452.t34 a_n2848_n452.t33 a_n1808_13878.t14 vdd.t109 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X102 a_n2848_n452.t20 a_n2848_n452.t19 a_n1808_13878.t13 vdd.t13 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X103 vdd.t157 a_n5644_8799.t53 CSoutput.t26 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X104 a_n5644_8799.t10 a_n2848_n452.t52 a_n1986_8322.t21 vdd.t90 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X105 gnd.t270 commonsourceibias.t80 CSoutput.t77 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 vdd.t156 a_n5644_8799.t54 CSoutput.t116 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 a_n2848_n452.t1 minus.t10 a_n3106_n452.t26 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X108 gnd.t269 commonsourceibias.t81 CSoutput.t76 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 gnd.t268 commonsourceibias.t4 commonsourceibias.t5 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X110 vdd.t182 CSoutput.t125 output.t15 gnd.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X111 vdd.t74 vdd.t72 vdd.t73 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X112 output.t14 CSoutput.t126 vdd.t178 gnd.t50 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X113 CSoutput.t127 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X114 output.t2 outputibias.t9 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X115 vdd.t155 a_n5644_8799.t55 CSoutput.t20 vdd.t140 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 vdd.t71 vdd.t69 vdd.t70 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X117 vdd.t68 vdd.t65 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 CSoutput.t75 commonsourceibias.t82 gnd.t267 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 a_n3106_n452.t33 diffpairibias.t18 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X120 outputibias.t5 outputibias.t4 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X121 vdd.t64 vdd.t61 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X122 gnd.t150 gnd.t148 minus.t4 gnd.t149 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X123 gnd.t147 gnd.t145 gnd.t146 gnd.t78 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X124 CSoutput.t74 commonsourceibias.t83 gnd.t266 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 gnd.t144 gnd.t142 gnd.t143 gnd.t92 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X126 output.t13 CSoutput.t128 vdd.t183 gnd.t51 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X127 vdd.t92 a_n2848_n452.t53 a_n1986_8322.t10 vdd.t91 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 vdd.t60 vdd.t58 vdd.t59 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X129 CSoutput.t36 a_n5644_8799.t56 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X130 a_n1986_8322.t9 a_n2848_n452.t54 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X131 outputibias.t3 outputibias.t2 gnd.t311 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X132 vdd.t152 a_n5644_8799.t57 CSoutput.t111 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X133 gnd.t141 gnd.t139 gnd.t140 gnd.t82 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X134 vdd.t197 a_n2848_n452.t55 a_n1808_13878.t6 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X135 gnd.t138 gnd.t136 plus.t3 gnd.t137 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X136 a_n2848_n452.t7 minus.t11 a_n3106_n452.t32 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X137 a_n5644_8799.t8 plus.t14 a_n3106_n452.t16 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X138 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 a_n5644_8799.t4 plus.t15 a_n3106_n452.t15 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X140 a_n2848_n452.t10 minus.t12 a_n3106_n452.t36 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X141 diffpairibias.t11 diffpairibias.t10 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X142 vdd.t53 vdd.t50 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X143 vdd.t150 a_n5644_8799.t58 CSoutput.t112 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X144 CSoutput.t73 commonsourceibias.t84 gnd.t264 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 gnd.t265 commonsourceibias.t85 CSoutput.t72 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 commonsourceibias.t3 commonsourceibias.t2 gnd.t263 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 a_n5644_8799.t6 a_n2848_n452.t56 a_n1986_8322.t20 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X148 a_n1986_8322.t8 a_n2848_n452.t57 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X149 vdd.t49 vdd.t46 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X150 vdd.t185 CSoutput.t129 output.t12 gnd.t323 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X151 a_n2848_n452.t22 a_n2848_n452.t21 a_n1808_13878.t12 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X152 a_n3106_n452.t30 minus.t13 a_n2848_n452.t5 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X153 CSoutput.t130 a_n1986_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X154 a_n5644_8799.t34 a_n2848_n452.t58 a_n1986_8322.t19 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 CSoutput.t71 commonsourceibias.t86 gnd.t262 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 CSoutput.t131 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X157 a_n1808_13878.t11 a_n2848_n452.t23 a_n2848_n452.t24 vdd.t90 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X158 gnd.t261 commonsourceibias.t87 CSoutput.t70 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 gnd.t260 commonsourceibias.t88 CSoutput.t69 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 a_n3106_n452.t14 plus.t16 a_n5644_8799.t27 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X161 a_n2848_n452.t3 minus.t14 a_n3106_n452.t28 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X162 commonsourceibias.t31 commonsourceibias.t30 gnd.t259 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 gnd.t257 commonsourceibias.t89 CSoutput.t68 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X164 vdd.t199 a_n2848_n452.t59 a_n1986_8322.t7 vdd.t198 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X165 CSoutput.t67 commonsourceibias.t90 gnd.t255 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 outputibias.t1 outputibias.t0 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X167 vdd.t45 vdd.t43 vdd.t44 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X168 gnd.t135 gnd.t132 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X169 a_n3106_n452.t41 diffpairibias.t19 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X170 CSoutput.t6 a_n5644_8799.t59 vdd.t148 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 a_n5644_8799.t17 plus.t17 a_n3106_n452.t13 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X172 a_n3106_n452.t52 diffpairibias.t20 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X173 output.t1 outputibias.t10 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X174 commonsourceibias.t29 commonsourceibias.t28 gnd.t254 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 vdd.t147 a_n5644_8799.t60 CSoutput.t114 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X176 gnd.t131 gnd.t129 gnd.t130 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X177 gnd.t128 gnd.t125 gnd.t127 gnd.t126 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X178 a_n5644_8799.t1 plus.t18 a_n3106_n452.t12 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X179 CSoutput.t66 commonsourceibias.t91 gnd.t252 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 CSoutput.t65 commonsourceibias.t92 gnd.t251 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 vdd.t146 a_n5644_8799.t61 CSoutput.t32 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 output.t11 CSoutput.t132 vdd.t188 gnd.t314 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X183 gnd.t124 gnd.t122 gnd.t123 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X184 minus.t3 gnd.t119 gnd.t121 gnd.t120 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X185 commonsourceibias.t27 commonsourceibias.t26 gnd.t250 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 diffpairibias.t9 diffpairibias.t8 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X187 CSoutput.t64 commonsourceibias.t93 gnd.t249 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 CSoutput.t63 commonsourceibias.t94 gnd.t248 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 a_n2848_n452.t13 minus.t15 a_n3106_n452.t39 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X190 output.t10 CSoutput.t133 vdd.t176 gnd.t315 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X191 a_n3106_n452.t11 plus.t19 a_n5644_8799.t20 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X192 gnd.t247 commonsourceibias.t16 commonsourceibias.t17 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 CSoutput.t8 a_n5644_8799.t62 vdd.t145 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X194 commonsourceibias.t15 commonsourceibias.t14 gnd.t245 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 vdd.t42 vdd.t40 vdd.t41 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X196 a_n1808_13878.t5 a_n2848_n452.t60 vdd.t4 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X197 vdd.t6 a_n2848_n452.t61 a_n1808_13878.t4 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X198 gnd.t243 commonsourceibias.t95 CSoutput.t62 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 commonsourceibias.t13 commonsourceibias.t12 gnd.t242 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X200 vdd.t39 vdd.t36 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X201 a_n3106_n452.t44 minus.t16 a_n2848_n452.t16 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X202 gnd.t241 commonsourceibias.t10 commonsourceibias.t11 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 gnd.t118 gnd.t116 gnd.t117 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X204 diffpairibias.t7 diffpairibias.t6 gnd.t327 gnd.t326 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X205 commonsourceibias.t9 commonsourceibias.t8 gnd.t240 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X206 CSoutput.t23 a_n5644_8799.t63 vdd.t144 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 vdd.t142 a_n5644_8799.t64 CSoutput.t15 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X208 a_n3106_n452.t46 minus.t17 a_n2848_n452.t42 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X209 a_n3106_n452.t10 plus.t20 a_n5644_8799.t33 gnd.t305 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X210 a_n1986_8322.t18 a_n2848_n452.t62 a_n5644_8799.t23 vdd.t111 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X211 gnd.t239 commonsourceibias.t96 CSoutput.t61 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 a_n3106_n452.t31 minus.t18 a_n2848_n452.t6 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X213 vdd.t187 CSoutput.t134 output.t9 gnd.t316 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X214 output.t0 outputibias.t11 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X215 vdd.t181 CSoutput.t135 output.t8 gnd.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X216 vdd.t141 a_n5644_8799.t65 CSoutput.t29 vdd.t140 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 CSoutput.t117 a_n5644_8799.t66 vdd.t139 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 gnd.t238 commonsourceibias.t6 commonsourceibias.t7 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 vdd.t138 a_n5644_8799.t67 CSoutput.t11 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 vdd.t193 a_n2848_n452.t63 a_n1986_8322.t6 vdd.t192 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X221 a_n1808_13878.t3 a_n2848_n452.t64 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X222 gnd.t115 gnd.t112 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X223 minus.t2 gnd.t109 gnd.t111 gnd.t110 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X224 a_n3106_n452.t53 diffpairibias.t21 gnd.t320 gnd.t319 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X225 CSoutput.t3 a_n5644_8799.t68 vdd.t137 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 a_n5644_8799.t3 plus.t21 a_n3106_n452.t9 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X227 a_n2848_n452.t11 minus.t19 a_n3106_n452.t37 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X228 gnd.t236 commonsourceibias.t46 commonsourceibias.t47 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 CSoutput.t35 a_n5644_8799.t69 vdd.t136 vdd.t131 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X230 a_n3106_n452.t35 minus.t20 a_n2848_n452.t9 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X231 CSoutput.t136 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X232 vdd.t35 vdd.t33 vdd.t34 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X233 a_n1986_8322.t17 a_n2848_n452.t65 a_n5644_8799.t2 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X234 vdd.t102 a_n2848_n452.t66 a_n1986_8322.t5 vdd.t101 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X235 vdd.t135 a_n5644_8799.t70 CSoutput.t25 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X236 CSoutput.t30 a_n5644_8799.t71 vdd.t134 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 a_n3106_n452.t27 minus.t21 a_n2848_n452.t2 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X238 gnd.t235 commonsourceibias.t44 commonsourceibias.t45 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 a_n3106_n452.t51 minus.t22 a_n2848_n452.t47 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X240 CSoutput.t60 commonsourceibias.t97 gnd.t234 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 vdd.t189 CSoutput.t137 output.t7 gnd.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X242 diffpairibias.t5 diffpairibias.t4 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X243 output.t6 CSoutput.t138 vdd.t184 gnd.t60 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X244 vdd.t32 vdd.t29 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X245 vdd.t28 vdd.t25 vdd.t27 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X246 gnd.t108 gnd.t105 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X247 a_n1808_13878.t10 a_n2848_n452.t35 a_n2848_n452.t36 vdd.t104 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X248 CSoutput.t59 commonsourceibias.t98 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X249 a_n1986_8322.t16 a_n2848_n452.t67 a_n5644_8799.t13 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X250 gnd.t104 gnd.t101 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X251 a_n3106_n452.t50 minus.t23 a_n2848_n452.t46 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X252 gnd.t230 commonsourceibias.t99 CSoutput.t58 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 gnd.t100 gnd.t98 gnd.t99 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X254 CSoutput.t17 a_n5644_8799.t72 vdd.t132 vdd.t131 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X255 a_n1986_8322.t4 a_n2848_n452.t68 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X256 gnd.t97 gnd.t95 plus.t2 gnd.t96 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X257 gnd.t94 gnd.t91 gnd.t93 gnd.t92 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X258 gnd.t229 commonsourceibias.t100 CSoutput.t57 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 gnd.t228 commonsourceibias.t101 CSoutput.t56 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 vdd.t108 a_n2848_n452.t69 a_n1808_13878.t2 vdd.t107 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X261 gnd.t90 gnd.t88 gnd.t89 gnd.t78 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X262 commonsourceibias.t43 commonsourceibias.t42 gnd.t227 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 gnd.t215 commonsourceibias.t102 CSoutput.t55 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 vdd.t191 CSoutput.t139 output.t5 gnd.t61 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X265 vdd.t24 vdd.t21 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X266 a_n1986_8322.t15 a_n2848_n452.t70 a_n5644_8799.t14 vdd.t97 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X267 a_n3106_n452.t8 plus.t22 a_n5644_8799.t5 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X268 vdd.t20 vdd.t18 vdd.t19 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X269 a_n5644_8799.t15 a_n2848_n452.t71 a_n1986_8322.t14 vdd.t104 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X270 a_n1808_13878.t1 a_n2848_n452.t72 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X271 vdd.t130 a_n5644_8799.t73 CSoutput.t12 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 CSoutput.t19 a_n5644_8799.t74 vdd.t128 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 gnd.t87 gnd.t85 minus.t1 gnd.t86 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X274 gnd.t214 commonsourceibias.t103 CSoutput.t54 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n2848_n452.t15 minus.t24 a_n3106_n452.t43 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X276 a_n5644_8799.t9 plus.t23 a_n3106_n452.t7 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X277 commonsourceibias.t19 commonsourceibias.t18 gnd.t217 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 a_n2848_n452.t0 minus.t25 a_n3106_n452.t1 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X279 gnd.t225 commonsourceibias.t104 CSoutput.t53 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 gnd.t223 commonsourceibias.t24 commonsourceibias.t25 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 gnd.t222 commonsourceibias.t22 commonsourceibias.t23 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X282 commonsourceibias.t21 commonsourceibias.t20 gnd.t221 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 CSoutput.t115 a_n5644_8799.t75 vdd.t126 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 a_n1808_13878.t9 a_n2848_n452.t29 a_n2848_n452.t30 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X285 a_n3106_n452.t38 minus.t26 a_n2848_n452.t12 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X286 a_n3106_n452.t54 diffpairibias.t22 gnd.t322 gnd.t321 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X287 gnd.t219 commonsourceibias.t105 CSoutput.t52 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 CSoutput.t51 commonsourceibias.t106 gnd.t212 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X289 gnd.t211 commonsourceibias.t107 CSoutput.t50 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 gnd.t84 gnd.t81 gnd.t83 gnd.t82 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X291 gnd.t80 gnd.t77 gnd.t79 gnd.t78 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X292 a_n5644_8799.t25 plus.t24 a_n3106_n452.t6 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X293 CSoutput.t34 a_n5644_8799.t76 vdd.t125 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 CSoutput.t49 commonsourceibias.t108 gnd.t209 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 gnd.t208 commonsourceibias.t109 CSoutput.t48 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X296 commonsourceibias.t37 commonsourceibias.t36 gnd.t206 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 vdd.t124 a_n5644_8799.t77 CSoutput.t27 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 gnd.t76 gnd.t73 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X299 diffpairibias.t3 diffpairibias.t2 gnd.t309 gnd.t308 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X300 a_n5644_8799.t12 a_n2848_n452.t73 a_n1986_8322.t13 vdd.t100 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X301 a_n2848_n452.t32 a_n2848_n452.t31 a_n1808_13878.t8 vdd.t97 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X302 gnd.t72 gnd.t70 plus.t1 gnd.t71 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X303 gnd.t203 commonsourceibias.t110 CSoutput.t47 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 a_n2848_n452.t41 minus.t27 a_n3106_n452.t45 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X305 vdd.t123 a_n5644_8799.t78 CSoutput.t2 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 vdd.t17 vdd.t14 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X307 CSoutput.t140 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X308 diffpairibias.t1 diffpairibias.t0 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X309 gnd.t204 commonsourceibias.t111 CSoutput.t46 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X310 commonsourceibias.t35 commonsourceibias.t34 gnd.t202 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 CSoutput.t45 commonsourceibias.t112 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X312 plus.t0 gnd.t67 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X313 gnd.t199 commonsourceibias.t32 commonsourceibias.t33 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 gnd.t66 gnd.t64 minus.t0 gnd.t65 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X315 a_n5644_8799.t22 plus.t25 a_n3106_n452.t5 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X316 vdd.t12 a_n2848_n452.t74 a_n1808_13878.t0 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X317 CSoutput.t21 a_n5644_8799.t79 vdd.t121 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 a_n5644_8799.t35 plus.t26 a_n3106_n452.t4 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X319 a_n2848_n452.t43 minus.t28 a_n3106_n452.t47 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X320 gnd.t197 commonsourceibias.t113 CSoutput.t44 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X321 gnd.t195 commonsourceibias.t114 CSoutput.t43 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 vdd.t186 CSoutput.t141 output.t4 gnd.t184 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X323 gnd.t193 commonsourceibias.t115 CSoutput.t42 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 CSoutput.t24 a_n5644_8799.t80 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 gnd.t192 commonsourceibias.t116 CSoutput.t41 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 vdd.t117 a_n5644_8799.t81 CSoutput.t118 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 a_n1986_8322.t12 a_n2848_n452.t75 a_n5644_8799.t7 vdd.t13 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X328 CSoutput.t40 commonsourceibias.t117 gnd.t190 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 gnd.t188 commonsourceibias.t118 CSoutput.t39 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 CSoutput.t38 commonsourceibias.t119 gnd.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 a_n3106_n452.t3 plus.t27 a_n5644_8799.t11 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X332 vdd.t115 a_n5644_8799.t82 CSoutput.t22 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X333 CSoutput.t110 a_n5644_8799.t83 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X334 a_n3106_n452.t2 plus.t28 a_n5644_8799.t32 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X335 a_n3106_n452.t40 diffpairibias.t23 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 commonsourceibias.n25 commonsourceibias.t8 230.006
R1 commonsourceibias.n91 commonsourceibias.t73 230.006
R2 commonsourceibias.n218 commonsourceibias.t98 230.006
R3 commonsourceibias.n154 commonsourceibias.t69 230.006
R4 commonsourceibias.n322 commonsourceibias.t4 230.006
R5 commonsourceibias.n281 commonsourceibias.t111 230.006
R6 commonsourceibias.n483 commonsourceibias.t113 230.006
R7 commonsourceibias.n419 commonsourceibias.t54 230.006
R8 commonsourceibias.n70 commonsourceibias.t22 207.983
R9 commonsourceibias.n136 commonsourceibias.t89 207.983
R10 commonsourceibias.n263 commonsourceibias.t109 207.983
R11 commonsourceibias.n199 commonsourceibias.t52 207.983
R12 commonsourceibias.n368 commonsourceibias.t12 207.983
R13 commonsourceibias.n402 commonsourceibias.t70 207.983
R14 commonsourceibias.n529 commonsourceibias.t63 207.983
R15 commonsourceibias.n465 commonsourceibias.t112 207.983
R16 commonsourceibias.n10 commonsourceibias.t2 168.701
R17 commonsourceibias.n63 commonsourceibias.t32 168.701
R18 commonsourceibias.n57 commonsourceibias.t20 168.701
R19 commonsourceibias.n16 commonsourceibias.t40 168.701
R20 commonsourceibias.n49 commonsourceibias.t18 168.701
R21 commonsourceibias.n43 commonsourceibias.t6 168.701
R22 commonsourceibias.n19 commonsourceibias.t34 168.701
R23 commonsourceibias.n21 commonsourceibias.t24 168.701
R24 commonsourceibias.n23 commonsourceibias.t28 168.701
R25 commonsourceibias.n26 commonsourceibias.t44 168.701
R26 commonsourceibias.n1 commonsourceibias.t49 168.701
R27 commonsourceibias.n129 commonsourceibias.t95 168.701
R28 commonsourceibias.n123 commonsourceibias.t90 168.701
R29 commonsourceibias.n7 commonsourceibias.t100 168.701
R30 commonsourceibias.n115 commonsourceibias.t86 168.701
R31 commonsourceibias.n109 commonsourceibias.t77 168.701
R32 commonsourceibias.n85 commonsourceibias.t94 168.701
R33 commonsourceibias.n87 commonsourceibias.t88 168.701
R34 commonsourceibias.n89 commonsourceibias.t60 168.701
R35 commonsourceibias.n92 commonsourceibias.t80 168.701
R36 commonsourceibias.n219 commonsourceibias.t102 168.701
R37 commonsourceibias.n216 commonsourceibias.t48 168.701
R38 commonsourceibias.n214 commonsourceibias.t103 168.701
R39 commonsourceibias.n212 commonsourceibias.t108 168.701
R40 commonsourceibias.n236 commonsourceibias.t87 168.701
R41 commonsourceibias.n242 commonsourceibias.t67 168.701
R42 commonsourceibias.n209 commonsourceibias.t115 168.701
R43 commonsourceibias.n250 commonsourceibias.t93 168.701
R44 commonsourceibias.n256 commonsourceibias.t96 168.701
R45 commonsourceibias.n203 commonsourceibias.t57 168.701
R46 commonsourceibias.n139 commonsourceibias.t119 168.701
R47 commonsourceibias.n192 commonsourceibias.t110 168.701
R48 commonsourceibias.n186 commonsourceibias.t59 168.701
R49 commonsourceibias.n145 commonsourceibias.t118 168.701
R50 commonsourceibias.n178 commonsourceibias.t65 168.701
R51 commonsourceibias.n172 commonsourceibias.t58 168.701
R52 commonsourceibias.n148 commonsourceibias.t117 168.701
R53 commonsourceibias.n150 commonsourceibias.t71 168.701
R54 commonsourceibias.n152 commonsourceibias.t83 168.701
R55 commonsourceibias.n155 commonsourceibias.t116 168.701
R56 commonsourceibias.n323 commonsourceibias.t26 168.701
R57 commonsourceibias.n320 commonsourceibias.t38 168.701
R58 commonsourceibias.n318 commonsourceibias.t14 168.701
R59 commonsourceibias.n316 commonsourceibias.t46 168.701
R60 commonsourceibias.n340 commonsourceibias.t30 168.701
R61 commonsourceibias.n346 commonsourceibias.t16 168.701
R62 commonsourceibias.n348 commonsourceibias.t36 168.701
R63 commonsourceibias.n355 commonsourceibias.t10 168.701
R64 commonsourceibias.n361 commonsourceibias.t42 168.701
R65 commonsourceibias.n308 commonsourceibias.t0 168.701
R66 commonsourceibias.n267 commonsourceibias.t99 168.701
R67 commonsourceibias.n395 commonsourceibias.t84 168.701
R68 commonsourceibias.n389 commonsourceibias.t72 168.701
R69 commonsourceibias.n382 commonsourceibias.t92 168.701
R70 commonsourceibias.n380 commonsourceibias.t66 168.701
R71 commonsourceibias.n282 commonsourceibias.t64 168.701
R72 commonsourceibias.n279 commonsourceibias.t104 168.701
R73 commonsourceibias.n277 commonsourceibias.t68 168.701
R74 commonsourceibias.n275 commonsourceibias.t79 168.701
R75 commonsourceibias.n299 commonsourceibias.t56 168.701
R76 commonsourceibias.n484 commonsourceibias.t97 168.701
R77 commonsourceibias.n481 commonsourceibias.t78 168.701
R78 commonsourceibias.n479 commonsourceibias.t53 168.701
R79 commonsourceibias.n477 commonsourceibias.t62 168.701
R80 commonsourceibias.n501 commonsourceibias.t82 168.701
R81 commonsourceibias.n507 commonsourceibias.t85 168.701
R82 commonsourceibias.n509 commonsourceibias.t74 168.701
R83 commonsourceibias.n516 commonsourceibias.t101 168.701
R84 commonsourceibias.n522 commonsourceibias.t91 168.701
R85 commonsourceibias.n469 commonsourceibias.t81 168.701
R86 commonsourceibias.n420 commonsourceibias.t61 168.701
R87 commonsourceibias.n417 commonsourceibias.t75 168.701
R88 commonsourceibias.n415 commonsourceibias.t55 168.701
R89 commonsourceibias.n413 commonsourceibias.t105 168.701
R90 commonsourceibias.n437 commonsourceibias.t76 168.701
R91 commonsourceibias.n443 commonsourceibias.t50 168.701
R92 commonsourceibias.n445 commonsourceibias.t106 168.701
R93 commonsourceibias.n452 commonsourceibias.t114 168.701
R94 commonsourceibias.n458 commonsourceibias.t51 168.701
R95 commonsourceibias.n405 commonsourceibias.t107 168.701
R96 commonsourceibias.n27 commonsourceibias.n24 161.3
R97 commonsourceibias.n29 commonsourceibias.n28 161.3
R98 commonsourceibias.n31 commonsourceibias.n30 161.3
R99 commonsourceibias.n32 commonsourceibias.n22 161.3
R100 commonsourceibias.n34 commonsourceibias.n33 161.3
R101 commonsourceibias.n36 commonsourceibias.n35 161.3
R102 commonsourceibias.n37 commonsourceibias.n20 161.3
R103 commonsourceibias.n39 commonsourceibias.n38 161.3
R104 commonsourceibias.n41 commonsourceibias.n40 161.3
R105 commonsourceibias.n42 commonsourceibias.n18 161.3
R106 commonsourceibias.n45 commonsourceibias.n44 161.3
R107 commonsourceibias.n46 commonsourceibias.n17 161.3
R108 commonsourceibias.n48 commonsourceibias.n47 161.3
R109 commonsourceibias.n50 commonsourceibias.n15 161.3
R110 commonsourceibias.n52 commonsourceibias.n51 161.3
R111 commonsourceibias.n53 commonsourceibias.n14 161.3
R112 commonsourceibias.n55 commonsourceibias.n54 161.3
R113 commonsourceibias.n56 commonsourceibias.n13 161.3
R114 commonsourceibias.n59 commonsourceibias.n58 161.3
R115 commonsourceibias.n60 commonsourceibias.n12 161.3
R116 commonsourceibias.n62 commonsourceibias.n61 161.3
R117 commonsourceibias.n64 commonsourceibias.n11 161.3
R118 commonsourceibias.n66 commonsourceibias.n65 161.3
R119 commonsourceibias.n68 commonsourceibias.n67 161.3
R120 commonsourceibias.n69 commonsourceibias.n9 161.3
R121 commonsourceibias.n93 commonsourceibias.n90 161.3
R122 commonsourceibias.n95 commonsourceibias.n94 161.3
R123 commonsourceibias.n97 commonsourceibias.n96 161.3
R124 commonsourceibias.n98 commonsourceibias.n88 161.3
R125 commonsourceibias.n100 commonsourceibias.n99 161.3
R126 commonsourceibias.n102 commonsourceibias.n101 161.3
R127 commonsourceibias.n103 commonsourceibias.n86 161.3
R128 commonsourceibias.n105 commonsourceibias.n104 161.3
R129 commonsourceibias.n107 commonsourceibias.n106 161.3
R130 commonsourceibias.n108 commonsourceibias.n84 161.3
R131 commonsourceibias.n111 commonsourceibias.n110 161.3
R132 commonsourceibias.n112 commonsourceibias.n8 161.3
R133 commonsourceibias.n114 commonsourceibias.n113 161.3
R134 commonsourceibias.n116 commonsourceibias.n6 161.3
R135 commonsourceibias.n118 commonsourceibias.n117 161.3
R136 commonsourceibias.n119 commonsourceibias.n5 161.3
R137 commonsourceibias.n121 commonsourceibias.n120 161.3
R138 commonsourceibias.n122 commonsourceibias.n4 161.3
R139 commonsourceibias.n125 commonsourceibias.n124 161.3
R140 commonsourceibias.n126 commonsourceibias.n3 161.3
R141 commonsourceibias.n128 commonsourceibias.n127 161.3
R142 commonsourceibias.n130 commonsourceibias.n2 161.3
R143 commonsourceibias.n132 commonsourceibias.n131 161.3
R144 commonsourceibias.n134 commonsourceibias.n133 161.3
R145 commonsourceibias.n135 commonsourceibias.n0 161.3
R146 commonsourceibias.n262 commonsourceibias.n202 161.3
R147 commonsourceibias.n261 commonsourceibias.n260 161.3
R148 commonsourceibias.n259 commonsourceibias.n258 161.3
R149 commonsourceibias.n257 commonsourceibias.n204 161.3
R150 commonsourceibias.n255 commonsourceibias.n254 161.3
R151 commonsourceibias.n253 commonsourceibias.n205 161.3
R152 commonsourceibias.n252 commonsourceibias.n251 161.3
R153 commonsourceibias.n249 commonsourceibias.n206 161.3
R154 commonsourceibias.n248 commonsourceibias.n247 161.3
R155 commonsourceibias.n246 commonsourceibias.n207 161.3
R156 commonsourceibias.n245 commonsourceibias.n244 161.3
R157 commonsourceibias.n243 commonsourceibias.n208 161.3
R158 commonsourceibias.n241 commonsourceibias.n240 161.3
R159 commonsourceibias.n239 commonsourceibias.n210 161.3
R160 commonsourceibias.n238 commonsourceibias.n237 161.3
R161 commonsourceibias.n235 commonsourceibias.n211 161.3
R162 commonsourceibias.n234 commonsourceibias.n233 161.3
R163 commonsourceibias.n232 commonsourceibias.n231 161.3
R164 commonsourceibias.n230 commonsourceibias.n213 161.3
R165 commonsourceibias.n229 commonsourceibias.n228 161.3
R166 commonsourceibias.n227 commonsourceibias.n226 161.3
R167 commonsourceibias.n225 commonsourceibias.n215 161.3
R168 commonsourceibias.n224 commonsourceibias.n223 161.3
R169 commonsourceibias.n222 commonsourceibias.n221 161.3
R170 commonsourceibias.n220 commonsourceibias.n217 161.3
R171 commonsourceibias.n156 commonsourceibias.n153 161.3
R172 commonsourceibias.n158 commonsourceibias.n157 161.3
R173 commonsourceibias.n160 commonsourceibias.n159 161.3
R174 commonsourceibias.n161 commonsourceibias.n151 161.3
R175 commonsourceibias.n163 commonsourceibias.n162 161.3
R176 commonsourceibias.n165 commonsourceibias.n164 161.3
R177 commonsourceibias.n166 commonsourceibias.n149 161.3
R178 commonsourceibias.n168 commonsourceibias.n167 161.3
R179 commonsourceibias.n170 commonsourceibias.n169 161.3
R180 commonsourceibias.n171 commonsourceibias.n147 161.3
R181 commonsourceibias.n174 commonsourceibias.n173 161.3
R182 commonsourceibias.n175 commonsourceibias.n146 161.3
R183 commonsourceibias.n177 commonsourceibias.n176 161.3
R184 commonsourceibias.n179 commonsourceibias.n144 161.3
R185 commonsourceibias.n181 commonsourceibias.n180 161.3
R186 commonsourceibias.n182 commonsourceibias.n143 161.3
R187 commonsourceibias.n184 commonsourceibias.n183 161.3
R188 commonsourceibias.n185 commonsourceibias.n142 161.3
R189 commonsourceibias.n188 commonsourceibias.n187 161.3
R190 commonsourceibias.n189 commonsourceibias.n141 161.3
R191 commonsourceibias.n191 commonsourceibias.n190 161.3
R192 commonsourceibias.n193 commonsourceibias.n140 161.3
R193 commonsourceibias.n195 commonsourceibias.n194 161.3
R194 commonsourceibias.n197 commonsourceibias.n196 161.3
R195 commonsourceibias.n198 commonsourceibias.n138 161.3
R196 commonsourceibias.n367 commonsourceibias.n307 161.3
R197 commonsourceibias.n366 commonsourceibias.n365 161.3
R198 commonsourceibias.n364 commonsourceibias.n363 161.3
R199 commonsourceibias.n362 commonsourceibias.n309 161.3
R200 commonsourceibias.n360 commonsourceibias.n359 161.3
R201 commonsourceibias.n358 commonsourceibias.n310 161.3
R202 commonsourceibias.n357 commonsourceibias.n356 161.3
R203 commonsourceibias.n354 commonsourceibias.n311 161.3
R204 commonsourceibias.n353 commonsourceibias.n352 161.3
R205 commonsourceibias.n351 commonsourceibias.n312 161.3
R206 commonsourceibias.n350 commonsourceibias.n349 161.3
R207 commonsourceibias.n347 commonsourceibias.n313 161.3
R208 commonsourceibias.n345 commonsourceibias.n344 161.3
R209 commonsourceibias.n343 commonsourceibias.n314 161.3
R210 commonsourceibias.n342 commonsourceibias.n341 161.3
R211 commonsourceibias.n339 commonsourceibias.n315 161.3
R212 commonsourceibias.n338 commonsourceibias.n337 161.3
R213 commonsourceibias.n336 commonsourceibias.n335 161.3
R214 commonsourceibias.n334 commonsourceibias.n317 161.3
R215 commonsourceibias.n333 commonsourceibias.n332 161.3
R216 commonsourceibias.n331 commonsourceibias.n330 161.3
R217 commonsourceibias.n329 commonsourceibias.n319 161.3
R218 commonsourceibias.n328 commonsourceibias.n327 161.3
R219 commonsourceibias.n326 commonsourceibias.n325 161.3
R220 commonsourceibias.n324 commonsourceibias.n321 161.3
R221 commonsourceibias.n301 commonsourceibias.n300 161.3
R222 commonsourceibias.n298 commonsourceibias.n274 161.3
R223 commonsourceibias.n297 commonsourceibias.n296 161.3
R224 commonsourceibias.n295 commonsourceibias.n294 161.3
R225 commonsourceibias.n293 commonsourceibias.n276 161.3
R226 commonsourceibias.n292 commonsourceibias.n291 161.3
R227 commonsourceibias.n290 commonsourceibias.n289 161.3
R228 commonsourceibias.n288 commonsourceibias.n278 161.3
R229 commonsourceibias.n287 commonsourceibias.n286 161.3
R230 commonsourceibias.n285 commonsourceibias.n284 161.3
R231 commonsourceibias.n283 commonsourceibias.n280 161.3
R232 commonsourceibias.n377 commonsourceibias.n273 161.3
R233 commonsourceibias.n401 commonsourceibias.n266 161.3
R234 commonsourceibias.n400 commonsourceibias.n399 161.3
R235 commonsourceibias.n398 commonsourceibias.n397 161.3
R236 commonsourceibias.n396 commonsourceibias.n268 161.3
R237 commonsourceibias.n394 commonsourceibias.n393 161.3
R238 commonsourceibias.n392 commonsourceibias.n269 161.3
R239 commonsourceibias.n391 commonsourceibias.n390 161.3
R240 commonsourceibias.n388 commonsourceibias.n270 161.3
R241 commonsourceibias.n387 commonsourceibias.n386 161.3
R242 commonsourceibias.n385 commonsourceibias.n271 161.3
R243 commonsourceibias.n384 commonsourceibias.n383 161.3
R244 commonsourceibias.n381 commonsourceibias.n272 161.3
R245 commonsourceibias.n379 commonsourceibias.n378 161.3
R246 commonsourceibias.n528 commonsourceibias.n468 161.3
R247 commonsourceibias.n527 commonsourceibias.n526 161.3
R248 commonsourceibias.n525 commonsourceibias.n524 161.3
R249 commonsourceibias.n523 commonsourceibias.n470 161.3
R250 commonsourceibias.n521 commonsourceibias.n520 161.3
R251 commonsourceibias.n519 commonsourceibias.n471 161.3
R252 commonsourceibias.n518 commonsourceibias.n517 161.3
R253 commonsourceibias.n515 commonsourceibias.n472 161.3
R254 commonsourceibias.n514 commonsourceibias.n513 161.3
R255 commonsourceibias.n512 commonsourceibias.n473 161.3
R256 commonsourceibias.n511 commonsourceibias.n510 161.3
R257 commonsourceibias.n508 commonsourceibias.n474 161.3
R258 commonsourceibias.n506 commonsourceibias.n505 161.3
R259 commonsourceibias.n504 commonsourceibias.n475 161.3
R260 commonsourceibias.n503 commonsourceibias.n502 161.3
R261 commonsourceibias.n500 commonsourceibias.n476 161.3
R262 commonsourceibias.n499 commonsourceibias.n498 161.3
R263 commonsourceibias.n497 commonsourceibias.n496 161.3
R264 commonsourceibias.n495 commonsourceibias.n478 161.3
R265 commonsourceibias.n494 commonsourceibias.n493 161.3
R266 commonsourceibias.n492 commonsourceibias.n491 161.3
R267 commonsourceibias.n490 commonsourceibias.n480 161.3
R268 commonsourceibias.n489 commonsourceibias.n488 161.3
R269 commonsourceibias.n487 commonsourceibias.n486 161.3
R270 commonsourceibias.n485 commonsourceibias.n482 161.3
R271 commonsourceibias.n464 commonsourceibias.n404 161.3
R272 commonsourceibias.n463 commonsourceibias.n462 161.3
R273 commonsourceibias.n461 commonsourceibias.n460 161.3
R274 commonsourceibias.n459 commonsourceibias.n406 161.3
R275 commonsourceibias.n457 commonsourceibias.n456 161.3
R276 commonsourceibias.n455 commonsourceibias.n407 161.3
R277 commonsourceibias.n454 commonsourceibias.n453 161.3
R278 commonsourceibias.n451 commonsourceibias.n408 161.3
R279 commonsourceibias.n450 commonsourceibias.n449 161.3
R280 commonsourceibias.n448 commonsourceibias.n409 161.3
R281 commonsourceibias.n447 commonsourceibias.n446 161.3
R282 commonsourceibias.n444 commonsourceibias.n410 161.3
R283 commonsourceibias.n442 commonsourceibias.n441 161.3
R284 commonsourceibias.n440 commonsourceibias.n411 161.3
R285 commonsourceibias.n439 commonsourceibias.n438 161.3
R286 commonsourceibias.n436 commonsourceibias.n412 161.3
R287 commonsourceibias.n435 commonsourceibias.n434 161.3
R288 commonsourceibias.n433 commonsourceibias.n432 161.3
R289 commonsourceibias.n431 commonsourceibias.n414 161.3
R290 commonsourceibias.n430 commonsourceibias.n429 161.3
R291 commonsourceibias.n428 commonsourceibias.n427 161.3
R292 commonsourceibias.n426 commonsourceibias.n416 161.3
R293 commonsourceibias.n425 commonsourceibias.n424 161.3
R294 commonsourceibias.n423 commonsourceibias.n422 161.3
R295 commonsourceibias.n421 commonsourceibias.n418 161.3
R296 commonsourceibias.n80 commonsourceibias.n78 81.5057
R297 commonsourceibias.n304 commonsourceibias.n302 81.5057
R298 commonsourceibias.n80 commonsourceibias.n79 80.9324
R299 commonsourceibias.n82 commonsourceibias.n81 80.9324
R300 commonsourceibias.n77 commonsourceibias.n76 80.9324
R301 commonsourceibias.n75 commonsourceibias.n74 80.9324
R302 commonsourceibias.n73 commonsourceibias.n72 80.9324
R303 commonsourceibias.n371 commonsourceibias.n370 80.9324
R304 commonsourceibias.n373 commonsourceibias.n372 80.9324
R305 commonsourceibias.n375 commonsourceibias.n374 80.9324
R306 commonsourceibias.n306 commonsourceibias.n305 80.9324
R307 commonsourceibias.n304 commonsourceibias.n303 80.9324
R308 commonsourceibias.n71 commonsourceibias.n70 80.6037
R309 commonsourceibias.n137 commonsourceibias.n136 80.6037
R310 commonsourceibias.n264 commonsourceibias.n263 80.6037
R311 commonsourceibias.n200 commonsourceibias.n199 80.6037
R312 commonsourceibias.n369 commonsourceibias.n368 80.6037
R313 commonsourceibias.n403 commonsourceibias.n402 80.6037
R314 commonsourceibias.n530 commonsourceibias.n529 80.6037
R315 commonsourceibias.n466 commonsourceibias.n465 80.6037
R316 commonsourceibias.n65 commonsourceibias.n64 56.5617
R317 commonsourceibias.n51 commonsourceibias.n50 56.5617
R318 commonsourceibias.n42 commonsourceibias.n41 56.5617
R319 commonsourceibias.n28 commonsourceibias.n27 56.5617
R320 commonsourceibias.n131 commonsourceibias.n130 56.5617
R321 commonsourceibias.n117 commonsourceibias.n116 56.5617
R322 commonsourceibias.n108 commonsourceibias.n107 56.5617
R323 commonsourceibias.n94 commonsourceibias.n93 56.5617
R324 commonsourceibias.n221 commonsourceibias.n220 56.5617
R325 commonsourceibias.n235 commonsourceibias.n234 56.5617
R326 commonsourceibias.n244 commonsourceibias.n243 56.5617
R327 commonsourceibias.n258 commonsourceibias.n257 56.5617
R328 commonsourceibias.n194 commonsourceibias.n193 56.5617
R329 commonsourceibias.n180 commonsourceibias.n179 56.5617
R330 commonsourceibias.n171 commonsourceibias.n170 56.5617
R331 commonsourceibias.n157 commonsourceibias.n156 56.5617
R332 commonsourceibias.n325 commonsourceibias.n324 56.5617
R333 commonsourceibias.n339 commonsourceibias.n338 56.5617
R334 commonsourceibias.n349 commonsourceibias.n347 56.5617
R335 commonsourceibias.n363 commonsourceibias.n362 56.5617
R336 commonsourceibias.n397 commonsourceibias.n396 56.5617
R337 commonsourceibias.n383 commonsourceibias.n381 56.5617
R338 commonsourceibias.n284 commonsourceibias.n283 56.5617
R339 commonsourceibias.n298 commonsourceibias.n297 56.5617
R340 commonsourceibias.n486 commonsourceibias.n485 56.5617
R341 commonsourceibias.n500 commonsourceibias.n499 56.5617
R342 commonsourceibias.n510 commonsourceibias.n508 56.5617
R343 commonsourceibias.n524 commonsourceibias.n523 56.5617
R344 commonsourceibias.n422 commonsourceibias.n421 56.5617
R345 commonsourceibias.n436 commonsourceibias.n435 56.5617
R346 commonsourceibias.n446 commonsourceibias.n444 56.5617
R347 commonsourceibias.n460 commonsourceibias.n459 56.5617
R348 commonsourceibias.n56 commonsourceibias.n55 56.0773
R349 commonsourceibias.n37 commonsourceibias.n36 56.0773
R350 commonsourceibias.n122 commonsourceibias.n121 56.0773
R351 commonsourceibias.n103 commonsourceibias.n102 56.0773
R352 commonsourceibias.n230 commonsourceibias.n229 56.0773
R353 commonsourceibias.n249 commonsourceibias.n248 56.0773
R354 commonsourceibias.n185 commonsourceibias.n184 56.0773
R355 commonsourceibias.n166 commonsourceibias.n165 56.0773
R356 commonsourceibias.n334 commonsourceibias.n333 56.0773
R357 commonsourceibias.n354 commonsourceibias.n353 56.0773
R358 commonsourceibias.n388 commonsourceibias.n387 56.0773
R359 commonsourceibias.n293 commonsourceibias.n292 56.0773
R360 commonsourceibias.n495 commonsourceibias.n494 56.0773
R361 commonsourceibias.n515 commonsourceibias.n514 56.0773
R362 commonsourceibias.n431 commonsourceibias.n430 56.0773
R363 commonsourceibias.n451 commonsourceibias.n450 56.0773
R364 commonsourceibias.n70 commonsourceibias.n69 46.0096
R365 commonsourceibias.n136 commonsourceibias.n135 46.0096
R366 commonsourceibias.n263 commonsourceibias.n262 46.0096
R367 commonsourceibias.n199 commonsourceibias.n198 46.0096
R368 commonsourceibias.n368 commonsourceibias.n367 46.0096
R369 commonsourceibias.n402 commonsourceibias.n401 46.0096
R370 commonsourceibias.n529 commonsourceibias.n528 46.0096
R371 commonsourceibias.n465 commonsourceibias.n464 46.0096
R372 commonsourceibias.n58 commonsourceibias.n12 41.5458
R373 commonsourceibias.n33 commonsourceibias.n32 41.5458
R374 commonsourceibias.n124 commonsourceibias.n3 41.5458
R375 commonsourceibias.n99 commonsourceibias.n98 41.5458
R376 commonsourceibias.n226 commonsourceibias.n225 41.5458
R377 commonsourceibias.n251 commonsourceibias.n205 41.5458
R378 commonsourceibias.n187 commonsourceibias.n141 41.5458
R379 commonsourceibias.n162 commonsourceibias.n161 41.5458
R380 commonsourceibias.n330 commonsourceibias.n329 41.5458
R381 commonsourceibias.n356 commonsourceibias.n310 41.5458
R382 commonsourceibias.n390 commonsourceibias.n269 41.5458
R383 commonsourceibias.n289 commonsourceibias.n288 41.5458
R384 commonsourceibias.n491 commonsourceibias.n490 41.5458
R385 commonsourceibias.n517 commonsourceibias.n471 41.5458
R386 commonsourceibias.n427 commonsourceibias.n426 41.5458
R387 commonsourceibias.n453 commonsourceibias.n407 41.5458
R388 commonsourceibias.n48 commonsourceibias.n17 40.577
R389 commonsourceibias.n44 commonsourceibias.n17 40.577
R390 commonsourceibias.n114 commonsourceibias.n8 40.577
R391 commonsourceibias.n110 commonsourceibias.n8 40.577
R392 commonsourceibias.n237 commonsourceibias.n210 40.577
R393 commonsourceibias.n241 commonsourceibias.n210 40.577
R394 commonsourceibias.n177 commonsourceibias.n146 40.577
R395 commonsourceibias.n173 commonsourceibias.n146 40.577
R396 commonsourceibias.n341 commonsourceibias.n314 40.577
R397 commonsourceibias.n345 commonsourceibias.n314 40.577
R398 commonsourceibias.n379 commonsourceibias.n273 40.577
R399 commonsourceibias.n300 commonsourceibias.n273 40.577
R400 commonsourceibias.n502 commonsourceibias.n475 40.577
R401 commonsourceibias.n506 commonsourceibias.n475 40.577
R402 commonsourceibias.n438 commonsourceibias.n411 40.577
R403 commonsourceibias.n442 commonsourceibias.n411 40.577
R404 commonsourceibias.n62 commonsourceibias.n12 39.6083
R405 commonsourceibias.n32 commonsourceibias.n31 39.6083
R406 commonsourceibias.n128 commonsourceibias.n3 39.6083
R407 commonsourceibias.n98 commonsourceibias.n97 39.6083
R408 commonsourceibias.n225 commonsourceibias.n224 39.6083
R409 commonsourceibias.n255 commonsourceibias.n205 39.6083
R410 commonsourceibias.n191 commonsourceibias.n141 39.6083
R411 commonsourceibias.n161 commonsourceibias.n160 39.6083
R412 commonsourceibias.n329 commonsourceibias.n328 39.6083
R413 commonsourceibias.n360 commonsourceibias.n310 39.6083
R414 commonsourceibias.n394 commonsourceibias.n269 39.6083
R415 commonsourceibias.n288 commonsourceibias.n287 39.6083
R416 commonsourceibias.n490 commonsourceibias.n489 39.6083
R417 commonsourceibias.n521 commonsourceibias.n471 39.6083
R418 commonsourceibias.n426 commonsourceibias.n425 39.6083
R419 commonsourceibias.n457 commonsourceibias.n407 39.6083
R420 commonsourceibias.n26 commonsourceibias.n25 33.0515
R421 commonsourceibias.n92 commonsourceibias.n91 33.0515
R422 commonsourceibias.n155 commonsourceibias.n154 33.0515
R423 commonsourceibias.n219 commonsourceibias.n218 33.0515
R424 commonsourceibias.n323 commonsourceibias.n322 33.0515
R425 commonsourceibias.n282 commonsourceibias.n281 33.0515
R426 commonsourceibias.n484 commonsourceibias.n483 33.0515
R427 commonsourceibias.n420 commonsourceibias.n419 33.0515
R428 commonsourceibias.n25 commonsourceibias.n24 28.5514
R429 commonsourceibias.n91 commonsourceibias.n90 28.5514
R430 commonsourceibias.n218 commonsourceibias.n217 28.5514
R431 commonsourceibias.n154 commonsourceibias.n153 28.5514
R432 commonsourceibias.n322 commonsourceibias.n321 28.5514
R433 commonsourceibias.n281 commonsourceibias.n280 28.5514
R434 commonsourceibias.n483 commonsourceibias.n482 28.5514
R435 commonsourceibias.n419 commonsourceibias.n418 28.5514
R436 commonsourceibias.n69 commonsourceibias.n68 26.0455
R437 commonsourceibias.n135 commonsourceibias.n134 26.0455
R438 commonsourceibias.n262 commonsourceibias.n261 26.0455
R439 commonsourceibias.n198 commonsourceibias.n197 26.0455
R440 commonsourceibias.n367 commonsourceibias.n366 26.0455
R441 commonsourceibias.n401 commonsourceibias.n400 26.0455
R442 commonsourceibias.n528 commonsourceibias.n527 26.0455
R443 commonsourceibias.n464 commonsourceibias.n463 26.0455
R444 commonsourceibias.n55 commonsourceibias.n14 25.0767
R445 commonsourceibias.n38 commonsourceibias.n37 25.0767
R446 commonsourceibias.n121 commonsourceibias.n5 25.0767
R447 commonsourceibias.n104 commonsourceibias.n103 25.0767
R448 commonsourceibias.n231 commonsourceibias.n230 25.0767
R449 commonsourceibias.n248 commonsourceibias.n207 25.0767
R450 commonsourceibias.n184 commonsourceibias.n143 25.0767
R451 commonsourceibias.n167 commonsourceibias.n166 25.0767
R452 commonsourceibias.n335 commonsourceibias.n334 25.0767
R453 commonsourceibias.n353 commonsourceibias.n312 25.0767
R454 commonsourceibias.n387 commonsourceibias.n271 25.0767
R455 commonsourceibias.n294 commonsourceibias.n293 25.0767
R456 commonsourceibias.n496 commonsourceibias.n495 25.0767
R457 commonsourceibias.n514 commonsourceibias.n473 25.0767
R458 commonsourceibias.n432 commonsourceibias.n431 25.0767
R459 commonsourceibias.n450 commonsourceibias.n409 25.0767
R460 commonsourceibias.n51 commonsourceibias.n16 24.3464
R461 commonsourceibias.n41 commonsourceibias.n19 24.3464
R462 commonsourceibias.n117 commonsourceibias.n7 24.3464
R463 commonsourceibias.n107 commonsourceibias.n85 24.3464
R464 commonsourceibias.n234 commonsourceibias.n212 24.3464
R465 commonsourceibias.n244 commonsourceibias.n209 24.3464
R466 commonsourceibias.n180 commonsourceibias.n145 24.3464
R467 commonsourceibias.n170 commonsourceibias.n148 24.3464
R468 commonsourceibias.n338 commonsourceibias.n316 24.3464
R469 commonsourceibias.n349 commonsourceibias.n348 24.3464
R470 commonsourceibias.n383 commonsourceibias.n382 24.3464
R471 commonsourceibias.n297 commonsourceibias.n275 24.3464
R472 commonsourceibias.n499 commonsourceibias.n477 24.3464
R473 commonsourceibias.n510 commonsourceibias.n509 24.3464
R474 commonsourceibias.n435 commonsourceibias.n413 24.3464
R475 commonsourceibias.n446 commonsourceibias.n445 24.3464
R476 commonsourceibias.n65 commonsourceibias.n10 23.8546
R477 commonsourceibias.n27 commonsourceibias.n26 23.8546
R478 commonsourceibias.n131 commonsourceibias.n1 23.8546
R479 commonsourceibias.n93 commonsourceibias.n92 23.8546
R480 commonsourceibias.n220 commonsourceibias.n219 23.8546
R481 commonsourceibias.n258 commonsourceibias.n203 23.8546
R482 commonsourceibias.n194 commonsourceibias.n139 23.8546
R483 commonsourceibias.n156 commonsourceibias.n155 23.8546
R484 commonsourceibias.n324 commonsourceibias.n323 23.8546
R485 commonsourceibias.n363 commonsourceibias.n308 23.8546
R486 commonsourceibias.n397 commonsourceibias.n267 23.8546
R487 commonsourceibias.n283 commonsourceibias.n282 23.8546
R488 commonsourceibias.n485 commonsourceibias.n484 23.8546
R489 commonsourceibias.n524 commonsourceibias.n469 23.8546
R490 commonsourceibias.n421 commonsourceibias.n420 23.8546
R491 commonsourceibias.n460 commonsourceibias.n405 23.8546
R492 commonsourceibias.n64 commonsourceibias.n63 16.9689
R493 commonsourceibias.n28 commonsourceibias.n23 16.9689
R494 commonsourceibias.n130 commonsourceibias.n129 16.9689
R495 commonsourceibias.n94 commonsourceibias.n89 16.9689
R496 commonsourceibias.n221 commonsourceibias.n216 16.9689
R497 commonsourceibias.n257 commonsourceibias.n256 16.9689
R498 commonsourceibias.n193 commonsourceibias.n192 16.9689
R499 commonsourceibias.n157 commonsourceibias.n152 16.9689
R500 commonsourceibias.n325 commonsourceibias.n320 16.9689
R501 commonsourceibias.n362 commonsourceibias.n361 16.9689
R502 commonsourceibias.n396 commonsourceibias.n395 16.9689
R503 commonsourceibias.n284 commonsourceibias.n279 16.9689
R504 commonsourceibias.n486 commonsourceibias.n481 16.9689
R505 commonsourceibias.n523 commonsourceibias.n522 16.9689
R506 commonsourceibias.n422 commonsourceibias.n417 16.9689
R507 commonsourceibias.n459 commonsourceibias.n458 16.9689
R508 commonsourceibias.n50 commonsourceibias.n49 16.477
R509 commonsourceibias.n43 commonsourceibias.n42 16.477
R510 commonsourceibias.n116 commonsourceibias.n115 16.477
R511 commonsourceibias.n109 commonsourceibias.n108 16.477
R512 commonsourceibias.n236 commonsourceibias.n235 16.477
R513 commonsourceibias.n243 commonsourceibias.n242 16.477
R514 commonsourceibias.n179 commonsourceibias.n178 16.477
R515 commonsourceibias.n172 commonsourceibias.n171 16.477
R516 commonsourceibias.n340 commonsourceibias.n339 16.477
R517 commonsourceibias.n347 commonsourceibias.n346 16.477
R518 commonsourceibias.n381 commonsourceibias.n380 16.477
R519 commonsourceibias.n299 commonsourceibias.n298 16.477
R520 commonsourceibias.n501 commonsourceibias.n500 16.477
R521 commonsourceibias.n508 commonsourceibias.n507 16.477
R522 commonsourceibias.n437 commonsourceibias.n436 16.477
R523 commonsourceibias.n444 commonsourceibias.n443 16.477
R524 commonsourceibias.n57 commonsourceibias.n56 15.9852
R525 commonsourceibias.n36 commonsourceibias.n21 15.9852
R526 commonsourceibias.n123 commonsourceibias.n122 15.9852
R527 commonsourceibias.n102 commonsourceibias.n87 15.9852
R528 commonsourceibias.n229 commonsourceibias.n214 15.9852
R529 commonsourceibias.n250 commonsourceibias.n249 15.9852
R530 commonsourceibias.n186 commonsourceibias.n185 15.9852
R531 commonsourceibias.n165 commonsourceibias.n150 15.9852
R532 commonsourceibias.n333 commonsourceibias.n318 15.9852
R533 commonsourceibias.n355 commonsourceibias.n354 15.9852
R534 commonsourceibias.n389 commonsourceibias.n388 15.9852
R535 commonsourceibias.n292 commonsourceibias.n277 15.9852
R536 commonsourceibias.n494 commonsourceibias.n479 15.9852
R537 commonsourceibias.n516 commonsourceibias.n515 15.9852
R538 commonsourceibias.n430 commonsourceibias.n415 15.9852
R539 commonsourceibias.n452 commonsourceibias.n451 15.9852
R540 commonsourceibias.n73 commonsourceibias.n71 13.2057
R541 commonsourceibias.n371 commonsourceibias.n369 13.2057
R542 commonsourceibias.n532 commonsourceibias.n265 10.122
R543 commonsourceibias.n112 commonsourceibias.n83 9.50363
R544 commonsourceibias.n377 commonsourceibias.n376 9.50363
R545 commonsourceibias.n201 commonsourceibias.n137 8.7339
R546 commonsourceibias.n467 commonsourceibias.n403 8.7339
R547 commonsourceibias.n58 commonsourceibias.n57 8.60764
R548 commonsourceibias.n33 commonsourceibias.n21 8.60764
R549 commonsourceibias.n124 commonsourceibias.n123 8.60764
R550 commonsourceibias.n99 commonsourceibias.n87 8.60764
R551 commonsourceibias.n226 commonsourceibias.n214 8.60764
R552 commonsourceibias.n251 commonsourceibias.n250 8.60764
R553 commonsourceibias.n187 commonsourceibias.n186 8.60764
R554 commonsourceibias.n162 commonsourceibias.n150 8.60764
R555 commonsourceibias.n330 commonsourceibias.n318 8.60764
R556 commonsourceibias.n356 commonsourceibias.n355 8.60764
R557 commonsourceibias.n390 commonsourceibias.n389 8.60764
R558 commonsourceibias.n289 commonsourceibias.n277 8.60764
R559 commonsourceibias.n491 commonsourceibias.n479 8.60764
R560 commonsourceibias.n517 commonsourceibias.n516 8.60764
R561 commonsourceibias.n427 commonsourceibias.n415 8.60764
R562 commonsourceibias.n453 commonsourceibias.n452 8.60764
R563 commonsourceibias.n532 commonsourceibias.n531 8.46921
R564 commonsourceibias.n49 commonsourceibias.n48 8.11581
R565 commonsourceibias.n44 commonsourceibias.n43 8.11581
R566 commonsourceibias.n115 commonsourceibias.n114 8.11581
R567 commonsourceibias.n110 commonsourceibias.n109 8.11581
R568 commonsourceibias.n237 commonsourceibias.n236 8.11581
R569 commonsourceibias.n242 commonsourceibias.n241 8.11581
R570 commonsourceibias.n178 commonsourceibias.n177 8.11581
R571 commonsourceibias.n173 commonsourceibias.n172 8.11581
R572 commonsourceibias.n341 commonsourceibias.n340 8.11581
R573 commonsourceibias.n346 commonsourceibias.n345 8.11581
R574 commonsourceibias.n380 commonsourceibias.n379 8.11581
R575 commonsourceibias.n300 commonsourceibias.n299 8.11581
R576 commonsourceibias.n502 commonsourceibias.n501 8.11581
R577 commonsourceibias.n507 commonsourceibias.n506 8.11581
R578 commonsourceibias.n438 commonsourceibias.n437 8.11581
R579 commonsourceibias.n443 commonsourceibias.n442 8.11581
R580 commonsourceibias.n63 commonsourceibias.n62 7.62397
R581 commonsourceibias.n31 commonsourceibias.n23 7.62397
R582 commonsourceibias.n129 commonsourceibias.n128 7.62397
R583 commonsourceibias.n97 commonsourceibias.n89 7.62397
R584 commonsourceibias.n224 commonsourceibias.n216 7.62397
R585 commonsourceibias.n256 commonsourceibias.n255 7.62397
R586 commonsourceibias.n192 commonsourceibias.n191 7.62397
R587 commonsourceibias.n160 commonsourceibias.n152 7.62397
R588 commonsourceibias.n328 commonsourceibias.n320 7.62397
R589 commonsourceibias.n361 commonsourceibias.n360 7.62397
R590 commonsourceibias.n395 commonsourceibias.n394 7.62397
R591 commonsourceibias.n287 commonsourceibias.n279 7.62397
R592 commonsourceibias.n489 commonsourceibias.n481 7.62397
R593 commonsourceibias.n522 commonsourceibias.n521 7.62397
R594 commonsourceibias.n425 commonsourceibias.n417 7.62397
R595 commonsourceibias.n458 commonsourceibias.n457 7.62397
R596 commonsourceibias.n265 commonsourceibias.n264 5.00473
R597 commonsourceibias.n201 commonsourceibias.n200 5.00473
R598 commonsourceibias.n531 commonsourceibias.n530 5.00473
R599 commonsourceibias.n467 commonsourceibias.n466 5.00473
R600 commonsourceibias commonsourceibias.n532 3.87639
R601 commonsourceibias.n265 commonsourceibias.n201 3.72967
R602 commonsourceibias.n531 commonsourceibias.n467 3.72967
R603 commonsourceibias.n78 commonsourceibias.t45 2.82907
R604 commonsourceibias.n78 commonsourceibias.t9 2.82907
R605 commonsourceibias.n79 commonsourceibias.t25 2.82907
R606 commonsourceibias.n79 commonsourceibias.t29 2.82907
R607 commonsourceibias.n81 commonsourceibias.t7 2.82907
R608 commonsourceibias.n81 commonsourceibias.t35 2.82907
R609 commonsourceibias.n76 commonsourceibias.t41 2.82907
R610 commonsourceibias.n76 commonsourceibias.t19 2.82907
R611 commonsourceibias.n74 commonsourceibias.t33 2.82907
R612 commonsourceibias.n74 commonsourceibias.t21 2.82907
R613 commonsourceibias.n72 commonsourceibias.t23 2.82907
R614 commonsourceibias.n72 commonsourceibias.t3 2.82907
R615 commonsourceibias.n370 commonsourceibias.t1 2.82907
R616 commonsourceibias.n370 commonsourceibias.t13 2.82907
R617 commonsourceibias.n372 commonsourceibias.t11 2.82907
R618 commonsourceibias.n372 commonsourceibias.t43 2.82907
R619 commonsourceibias.n374 commonsourceibias.t17 2.82907
R620 commonsourceibias.n374 commonsourceibias.t37 2.82907
R621 commonsourceibias.n305 commonsourceibias.t47 2.82907
R622 commonsourceibias.n305 commonsourceibias.t31 2.82907
R623 commonsourceibias.n303 commonsourceibias.t39 2.82907
R624 commonsourceibias.n303 commonsourceibias.t15 2.82907
R625 commonsourceibias.n302 commonsourceibias.t5 2.82907
R626 commonsourceibias.n302 commonsourceibias.t27 2.82907
R627 commonsourceibias.n68 commonsourceibias.n10 0.738255
R628 commonsourceibias.n134 commonsourceibias.n1 0.738255
R629 commonsourceibias.n261 commonsourceibias.n203 0.738255
R630 commonsourceibias.n197 commonsourceibias.n139 0.738255
R631 commonsourceibias.n366 commonsourceibias.n308 0.738255
R632 commonsourceibias.n400 commonsourceibias.n267 0.738255
R633 commonsourceibias.n527 commonsourceibias.n469 0.738255
R634 commonsourceibias.n463 commonsourceibias.n405 0.738255
R635 commonsourceibias.n75 commonsourceibias.n73 0.573776
R636 commonsourceibias.n77 commonsourceibias.n75 0.573776
R637 commonsourceibias.n82 commonsourceibias.n80 0.573776
R638 commonsourceibias.n306 commonsourceibias.n304 0.573776
R639 commonsourceibias.n375 commonsourceibias.n373 0.573776
R640 commonsourceibias.n373 commonsourceibias.n371 0.573776
R641 commonsourceibias.n83 commonsourceibias.n77 0.287138
R642 commonsourceibias.n83 commonsourceibias.n82 0.287138
R643 commonsourceibias.n376 commonsourceibias.n306 0.287138
R644 commonsourceibias.n376 commonsourceibias.n375 0.287138
R645 commonsourceibias.n71 commonsourceibias.n9 0.285035
R646 commonsourceibias.n137 commonsourceibias.n0 0.285035
R647 commonsourceibias.n264 commonsourceibias.n202 0.285035
R648 commonsourceibias.n200 commonsourceibias.n138 0.285035
R649 commonsourceibias.n369 commonsourceibias.n307 0.285035
R650 commonsourceibias.n403 commonsourceibias.n266 0.285035
R651 commonsourceibias.n530 commonsourceibias.n468 0.285035
R652 commonsourceibias.n466 commonsourceibias.n404 0.285035
R653 commonsourceibias.n16 commonsourceibias.n14 0.246418
R654 commonsourceibias.n38 commonsourceibias.n19 0.246418
R655 commonsourceibias.n7 commonsourceibias.n5 0.246418
R656 commonsourceibias.n104 commonsourceibias.n85 0.246418
R657 commonsourceibias.n231 commonsourceibias.n212 0.246418
R658 commonsourceibias.n209 commonsourceibias.n207 0.246418
R659 commonsourceibias.n145 commonsourceibias.n143 0.246418
R660 commonsourceibias.n167 commonsourceibias.n148 0.246418
R661 commonsourceibias.n335 commonsourceibias.n316 0.246418
R662 commonsourceibias.n348 commonsourceibias.n312 0.246418
R663 commonsourceibias.n382 commonsourceibias.n271 0.246418
R664 commonsourceibias.n294 commonsourceibias.n275 0.246418
R665 commonsourceibias.n496 commonsourceibias.n477 0.246418
R666 commonsourceibias.n509 commonsourceibias.n473 0.246418
R667 commonsourceibias.n432 commonsourceibias.n413 0.246418
R668 commonsourceibias.n445 commonsourceibias.n409 0.246418
R669 commonsourceibias.n67 commonsourceibias.n9 0.189894
R670 commonsourceibias.n67 commonsourceibias.n66 0.189894
R671 commonsourceibias.n66 commonsourceibias.n11 0.189894
R672 commonsourceibias.n61 commonsourceibias.n11 0.189894
R673 commonsourceibias.n61 commonsourceibias.n60 0.189894
R674 commonsourceibias.n60 commonsourceibias.n59 0.189894
R675 commonsourceibias.n59 commonsourceibias.n13 0.189894
R676 commonsourceibias.n54 commonsourceibias.n13 0.189894
R677 commonsourceibias.n54 commonsourceibias.n53 0.189894
R678 commonsourceibias.n53 commonsourceibias.n52 0.189894
R679 commonsourceibias.n52 commonsourceibias.n15 0.189894
R680 commonsourceibias.n47 commonsourceibias.n15 0.189894
R681 commonsourceibias.n47 commonsourceibias.n46 0.189894
R682 commonsourceibias.n46 commonsourceibias.n45 0.189894
R683 commonsourceibias.n45 commonsourceibias.n18 0.189894
R684 commonsourceibias.n40 commonsourceibias.n18 0.189894
R685 commonsourceibias.n40 commonsourceibias.n39 0.189894
R686 commonsourceibias.n39 commonsourceibias.n20 0.189894
R687 commonsourceibias.n35 commonsourceibias.n20 0.189894
R688 commonsourceibias.n35 commonsourceibias.n34 0.189894
R689 commonsourceibias.n34 commonsourceibias.n22 0.189894
R690 commonsourceibias.n30 commonsourceibias.n22 0.189894
R691 commonsourceibias.n30 commonsourceibias.n29 0.189894
R692 commonsourceibias.n29 commonsourceibias.n24 0.189894
R693 commonsourceibias.n111 commonsourceibias.n84 0.189894
R694 commonsourceibias.n106 commonsourceibias.n84 0.189894
R695 commonsourceibias.n106 commonsourceibias.n105 0.189894
R696 commonsourceibias.n105 commonsourceibias.n86 0.189894
R697 commonsourceibias.n101 commonsourceibias.n86 0.189894
R698 commonsourceibias.n101 commonsourceibias.n100 0.189894
R699 commonsourceibias.n100 commonsourceibias.n88 0.189894
R700 commonsourceibias.n96 commonsourceibias.n88 0.189894
R701 commonsourceibias.n96 commonsourceibias.n95 0.189894
R702 commonsourceibias.n95 commonsourceibias.n90 0.189894
R703 commonsourceibias.n133 commonsourceibias.n0 0.189894
R704 commonsourceibias.n133 commonsourceibias.n132 0.189894
R705 commonsourceibias.n132 commonsourceibias.n2 0.189894
R706 commonsourceibias.n127 commonsourceibias.n2 0.189894
R707 commonsourceibias.n127 commonsourceibias.n126 0.189894
R708 commonsourceibias.n126 commonsourceibias.n125 0.189894
R709 commonsourceibias.n125 commonsourceibias.n4 0.189894
R710 commonsourceibias.n120 commonsourceibias.n4 0.189894
R711 commonsourceibias.n120 commonsourceibias.n119 0.189894
R712 commonsourceibias.n119 commonsourceibias.n118 0.189894
R713 commonsourceibias.n118 commonsourceibias.n6 0.189894
R714 commonsourceibias.n113 commonsourceibias.n6 0.189894
R715 commonsourceibias.n260 commonsourceibias.n202 0.189894
R716 commonsourceibias.n260 commonsourceibias.n259 0.189894
R717 commonsourceibias.n259 commonsourceibias.n204 0.189894
R718 commonsourceibias.n254 commonsourceibias.n204 0.189894
R719 commonsourceibias.n254 commonsourceibias.n253 0.189894
R720 commonsourceibias.n253 commonsourceibias.n252 0.189894
R721 commonsourceibias.n252 commonsourceibias.n206 0.189894
R722 commonsourceibias.n247 commonsourceibias.n206 0.189894
R723 commonsourceibias.n247 commonsourceibias.n246 0.189894
R724 commonsourceibias.n246 commonsourceibias.n245 0.189894
R725 commonsourceibias.n245 commonsourceibias.n208 0.189894
R726 commonsourceibias.n240 commonsourceibias.n208 0.189894
R727 commonsourceibias.n240 commonsourceibias.n239 0.189894
R728 commonsourceibias.n239 commonsourceibias.n238 0.189894
R729 commonsourceibias.n238 commonsourceibias.n211 0.189894
R730 commonsourceibias.n233 commonsourceibias.n211 0.189894
R731 commonsourceibias.n233 commonsourceibias.n232 0.189894
R732 commonsourceibias.n232 commonsourceibias.n213 0.189894
R733 commonsourceibias.n228 commonsourceibias.n213 0.189894
R734 commonsourceibias.n228 commonsourceibias.n227 0.189894
R735 commonsourceibias.n227 commonsourceibias.n215 0.189894
R736 commonsourceibias.n223 commonsourceibias.n215 0.189894
R737 commonsourceibias.n223 commonsourceibias.n222 0.189894
R738 commonsourceibias.n222 commonsourceibias.n217 0.189894
R739 commonsourceibias.n196 commonsourceibias.n138 0.189894
R740 commonsourceibias.n196 commonsourceibias.n195 0.189894
R741 commonsourceibias.n195 commonsourceibias.n140 0.189894
R742 commonsourceibias.n190 commonsourceibias.n140 0.189894
R743 commonsourceibias.n190 commonsourceibias.n189 0.189894
R744 commonsourceibias.n189 commonsourceibias.n188 0.189894
R745 commonsourceibias.n188 commonsourceibias.n142 0.189894
R746 commonsourceibias.n183 commonsourceibias.n142 0.189894
R747 commonsourceibias.n183 commonsourceibias.n182 0.189894
R748 commonsourceibias.n182 commonsourceibias.n181 0.189894
R749 commonsourceibias.n181 commonsourceibias.n144 0.189894
R750 commonsourceibias.n176 commonsourceibias.n144 0.189894
R751 commonsourceibias.n176 commonsourceibias.n175 0.189894
R752 commonsourceibias.n175 commonsourceibias.n174 0.189894
R753 commonsourceibias.n174 commonsourceibias.n147 0.189894
R754 commonsourceibias.n169 commonsourceibias.n147 0.189894
R755 commonsourceibias.n169 commonsourceibias.n168 0.189894
R756 commonsourceibias.n168 commonsourceibias.n149 0.189894
R757 commonsourceibias.n164 commonsourceibias.n149 0.189894
R758 commonsourceibias.n164 commonsourceibias.n163 0.189894
R759 commonsourceibias.n163 commonsourceibias.n151 0.189894
R760 commonsourceibias.n159 commonsourceibias.n151 0.189894
R761 commonsourceibias.n159 commonsourceibias.n158 0.189894
R762 commonsourceibias.n158 commonsourceibias.n153 0.189894
R763 commonsourceibias.n326 commonsourceibias.n321 0.189894
R764 commonsourceibias.n327 commonsourceibias.n326 0.189894
R765 commonsourceibias.n327 commonsourceibias.n319 0.189894
R766 commonsourceibias.n331 commonsourceibias.n319 0.189894
R767 commonsourceibias.n332 commonsourceibias.n331 0.189894
R768 commonsourceibias.n332 commonsourceibias.n317 0.189894
R769 commonsourceibias.n336 commonsourceibias.n317 0.189894
R770 commonsourceibias.n337 commonsourceibias.n336 0.189894
R771 commonsourceibias.n337 commonsourceibias.n315 0.189894
R772 commonsourceibias.n342 commonsourceibias.n315 0.189894
R773 commonsourceibias.n343 commonsourceibias.n342 0.189894
R774 commonsourceibias.n344 commonsourceibias.n343 0.189894
R775 commonsourceibias.n344 commonsourceibias.n313 0.189894
R776 commonsourceibias.n350 commonsourceibias.n313 0.189894
R777 commonsourceibias.n351 commonsourceibias.n350 0.189894
R778 commonsourceibias.n352 commonsourceibias.n351 0.189894
R779 commonsourceibias.n352 commonsourceibias.n311 0.189894
R780 commonsourceibias.n357 commonsourceibias.n311 0.189894
R781 commonsourceibias.n358 commonsourceibias.n357 0.189894
R782 commonsourceibias.n359 commonsourceibias.n358 0.189894
R783 commonsourceibias.n359 commonsourceibias.n309 0.189894
R784 commonsourceibias.n364 commonsourceibias.n309 0.189894
R785 commonsourceibias.n365 commonsourceibias.n364 0.189894
R786 commonsourceibias.n365 commonsourceibias.n307 0.189894
R787 commonsourceibias.n285 commonsourceibias.n280 0.189894
R788 commonsourceibias.n286 commonsourceibias.n285 0.189894
R789 commonsourceibias.n286 commonsourceibias.n278 0.189894
R790 commonsourceibias.n290 commonsourceibias.n278 0.189894
R791 commonsourceibias.n291 commonsourceibias.n290 0.189894
R792 commonsourceibias.n291 commonsourceibias.n276 0.189894
R793 commonsourceibias.n295 commonsourceibias.n276 0.189894
R794 commonsourceibias.n296 commonsourceibias.n295 0.189894
R795 commonsourceibias.n296 commonsourceibias.n274 0.189894
R796 commonsourceibias.n301 commonsourceibias.n274 0.189894
R797 commonsourceibias.n378 commonsourceibias.n272 0.189894
R798 commonsourceibias.n384 commonsourceibias.n272 0.189894
R799 commonsourceibias.n385 commonsourceibias.n384 0.189894
R800 commonsourceibias.n386 commonsourceibias.n385 0.189894
R801 commonsourceibias.n386 commonsourceibias.n270 0.189894
R802 commonsourceibias.n391 commonsourceibias.n270 0.189894
R803 commonsourceibias.n392 commonsourceibias.n391 0.189894
R804 commonsourceibias.n393 commonsourceibias.n392 0.189894
R805 commonsourceibias.n393 commonsourceibias.n268 0.189894
R806 commonsourceibias.n398 commonsourceibias.n268 0.189894
R807 commonsourceibias.n399 commonsourceibias.n398 0.189894
R808 commonsourceibias.n399 commonsourceibias.n266 0.189894
R809 commonsourceibias.n487 commonsourceibias.n482 0.189894
R810 commonsourceibias.n488 commonsourceibias.n487 0.189894
R811 commonsourceibias.n488 commonsourceibias.n480 0.189894
R812 commonsourceibias.n492 commonsourceibias.n480 0.189894
R813 commonsourceibias.n493 commonsourceibias.n492 0.189894
R814 commonsourceibias.n493 commonsourceibias.n478 0.189894
R815 commonsourceibias.n497 commonsourceibias.n478 0.189894
R816 commonsourceibias.n498 commonsourceibias.n497 0.189894
R817 commonsourceibias.n498 commonsourceibias.n476 0.189894
R818 commonsourceibias.n503 commonsourceibias.n476 0.189894
R819 commonsourceibias.n504 commonsourceibias.n503 0.189894
R820 commonsourceibias.n505 commonsourceibias.n504 0.189894
R821 commonsourceibias.n505 commonsourceibias.n474 0.189894
R822 commonsourceibias.n511 commonsourceibias.n474 0.189894
R823 commonsourceibias.n512 commonsourceibias.n511 0.189894
R824 commonsourceibias.n513 commonsourceibias.n512 0.189894
R825 commonsourceibias.n513 commonsourceibias.n472 0.189894
R826 commonsourceibias.n518 commonsourceibias.n472 0.189894
R827 commonsourceibias.n519 commonsourceibias.n518 0.189894
R828 commonsourceibias.n520 commonsourceibias.n519 0.189894
R829 commonsourceibias.n520 commonsourceibias.n470 0.189894
R830 commonsourceibias.n525 commonsourceibias.n470 0.189894
R831 commonsourceibias.n526 commonsourceibias.n525 0.189894
R832 commonsourceibias.n526 commonsourceibias.n468 0.189894
R833 commonsourceibias.n423 commonsourceibias.n418 0.189894
R834 commonsourceibias.n424 commonsourceibias.n423 0.189894
R835 commonsourceibias.n424 commonsourceibias.n416 0.189894
R836 commonsourceibias.n428 commonsourceibias.n416 0.189894
R837 commonsourceibias.n429 commonsourceibias.n428 0.189894
R838 commonsourceibias.n429 commonsourceibias.n414 0.189894
R839 commonsourceibias.n433 commonsourceibias.n414 0.189894
R840 commonsourceibias.n434 commonsourceibias.n433 0.189894
R841 commonsourceibias.n434 commonsourceibias.n412 0.189894
R842 commonsourceibias.n439 commonsourceibias.n412 0.189894
R843 commonsourceibias.n440 commonsourceibias.n439 0.189894
R844 commonsourceibias.n441 commonsourceibias.n440 0.189894
R845 commonsourceibias.n441 commonsourceibias.n410 0.189894
R846 commonsourceibias.n447 commonsourceibias.n410 0.189894
R847 commonsourceibias.n448 commonsourceibias.n447 0.189894
R848 commonsourceibias.n449 commonsourceibias.n448 0.189894
R849 commonsourceibias.n449 commonsourceibias.n408 0.189894
R850 commonsourceibias.n454 commonsourceibias.n408 0.189894
R851 commonsourceibias.n455 commonsourceibias.n454 0.189894
R852 commonsourceibias.n456 commonsourceibias.n455 0.189894
R853 commonsourceibias.n456 commonsourceibias.n406 0.189894
R854 commonsourceibias.n461 commonsourceibias.n406 0.189894
R855 commonsourceibias.n462 commonsourceibias.n461 0.189894
R856 commonsourceibias.n462 commonsourceibias.n404 0.189894
R857 commonsourceibias.n112 commonsourceibias.n111 0.170955
R858 commonsourceibias.n113 commonsourceibias.n112 0.170955
R859 commonsourceibias.n377 commonsourceibias.n301 0.170955
R860 commonsourceibias.n378 commonsourceibias.n377 0.170955
R861 gnd.n6638 gnd.n687 1087.89
R862 gnd.n4241 gnd.n3905 939.716
R863 gnd.n6968 gnd.n166 838.452
R864 gnd.n198 gnd.n164 838.452
R865 gnd.n1668 gnd.n1556 838.452
R866 gnd.n5633 gnd.n1670 838.452
R867 gnd.n1145 gnd.n1133 838.452
R868 gnd.n4716 gnd.n4715 838.452
R869 gnd.n4081 gnd.n3942 838.452
R870 gnd.n4120 gnd.n2433 838.452
R871 gnd.n6970 gnd.n161 783.196
R872 gnd.n490 gnd.n163 783.196
R873 gnd.n5636 gnd.n5635 783.196
R874 gnd.n5753 gnd.n1602 783.196
R875 gnd.n6085 gnd.n1138 783.196
R876 gnd.n4668 gnd.n2296 783.196
R877 gnd.n4244 gnd.n4243 783.196
R878 gnd.n4239 gnd.n2429 783.196
R879 gnd.n4756 gnd.n2263 771.183
R880 gnd.n5822 gnd.n1492 771.183
R881 gnd.n4737 gnd.n2266 771.183
R882 gnd.n5824 gnd.n1487 771.183
R883 gnd.n3813 gnd.n2444 766.379
R884 gnd.n3816 gnd.n3815 766.379
R885 gnd.n3054 gnd.n2957 766.379
R886 gnd.n3050 gnd.n2955 766.379
R887 gnd.n3904 gnd.n2466 756.769
R888 gnd.n3807 gnd.n3806 756.769
R889 gnd.n3147 gnd.n2864 756.769
R890 gnd.n3145 gnd.n2867 756.769
R891 gnd.n6310 gnd.n879 655.866
R892 gnd.n6637 gnd.n688 655.866
R893 gnd.n6850 gnd.n6849 655.866
R894 gnd.n6142 gnd.n1049 655.866
R895 gnd.n6311 gnd.n6310 585
R896 gnd.n6310 gnd.n6309 585
R897 gnd.n883 gnd.n882 585
R898 gnd.n6308 gnd.n883 585
R899 gnd.n6306 gnd.n6305 585
R900 gnd.n6307 gnd.n6306 585
R901 gnd.n6304 gnd.n885 585
R902 gnd.n885 gnd.n884 585
R903 gnd.n6303 gnd.n6302 585
R904 gnd.n6302 gnd.n6301 585
R905 gnd.n890 gnd.n889 585
R906 gnd.n6300 gnd.n890 585
R907 gnd.n6298 gnd.n6297 585
R908 gnd.n6299 gnd.n6298 585
R909 gnd.n6296 gnd.n892 585
R910 gnd.n892 gnd.n891 585
R911 gnd.n6295 gnd.n6294 585
R912 gnd.n6294 gnd.n6293 585
R913 gnd.n898 gnd.n897 585
R914 gnd.n6292 gnd.n898 585
R915 gnd.n6290 gnd.n6289 585
R916 gnd.n6291 gnd.n6290 585
R917 gnd.n6288 gnd.n900 585
R918 gnd.n900 gnd.n899 585
R919 gnd.n6287 gnd.n6286 585
R920 gnd.n6286 gnd.n6285 585
R921 gnd.n906 gnd.n905 585
R922 gnd.n6284 gnd.n906 585
R923 gnd.n6282 gnd.n6281 585
R924 gnd.n6283 gnd.n6282 585
R925 gnd.n6280 gnd.n908 585
R926 gnd.n908 gnd.n907 585
R927 gnd.n6279 gnd.n6278 585
R928 gnd.n6278 gnd.n6277 585
R929 gnd.n914 gnd.n913 585
R930 gnd.n6276 gnd.n914 585
R931 gnd.n6274 gnd.n6273 585
R932 gnd.n6275 gnd.n6274 585
R933 gnd.n6272 gnd.n916 585
R934 gnd.n916 gnd.n915 585
R935 gnd.n6271 gnd.n6270 585
R936 gnd.n6270 gnd.n6269 585
R937 gnd.n922 gnd.n921 585
R938 gnd.n6268 gnd.n922 585
R939 gnd.n6266 gnd.n6265 585
R940 gnd.n6267 gnd.n6266 585
R941 gnd.n6264 gnd.n924 585
R942 gnd.n924 gnd.n923 585
R943 gnd.n6263 gnd.n6262 585
R944 gnd.n6262 gnd.n6261 585
R945 gnd.n930 gnd.n929 585
R946 gnd.n6260 gnd.n930 585
R947 gnd.n6258 gnd.n6257 585
R948 gnd.n6259 gnd.n6258 585
R949 gnd.n6256 gnd.n932 585
R950 gnd.n932 gnd.n931 585
R951 gnd.n6255 gnd.n6254 585
R952 gnd.n6254 gnd.n6253 585
R953 gnd.n938 gnd.n937 585
R954 gnd.n6252 gnd.n938 585
R955 gnd.n6250 gnd.n6249 585
R956 gnd.n6251 gnd.n6250 585
R957 gnd.n6248 gnd.n940 585
R958 gnd.n940 gnd.n939 585
R959 gnd.n6247 gnd.n6246 585
R960 gnd.n6246 gnd.n6245 585
R961 gnd.n946 gnd.n945 585
R962 gnd.n6244 gnd.n946 585
R963 gnd.n6242 gnd.n6241 585
R964 gnd.n6243 gnd.n6242 585
R965 gnd.n6240 gnd.n948 585
R966 gnd.n948 gnd.n947 585
R967 gnd.n6239 gnd.n6238 585
R968 gnd.n6238 gnd.n6237 585
R969 gnd.n954 gnd.n953 585
R970 gnd.n6236 gnd.n954 585
R971 gnd.n6234 gnd.n6233 585
R972 gnd.n6235 gnd.n6234 585
R973 gnd.n6232 gnd.n956 585
R974 gnd.n956 gnd.n955 585
R975 gnd.n6231 gnd.n6230 585
R976 gnd.n6230 gnd.n6229 585
R977 gnd.n962 gnd.n961 585
R978 gnd.n6228 gnd.n962 585
R979 gnd.n6226 gnd.n6225 585
R980 gnd.n6227 gnd.n6226 585
R981 gnd.n6224 gnd.n964 585
R982 gnd.n964 gnd.n963 585
R983 gnd.n6223 gnd.n6222 585
R984 gnd.n6222 gnd.n6221 585
R985 gnd.n970 gnd.n969 585
R986 gnd.n6220 gnd.n970 585
R987 gnd.n6218 gnd.n6217 585
R988 gnd.n6219 gnd.n6218 585
R989 gnd.n6216 gnd.n972 585
R990 gnd.n972 gnd.n971 585
R991 gnd.n6215 gnd.n6214 585
R992 gnd.n6214 gnd.n6213 585
R993 gnd.n978 gnd.n977 585
R994 gnd.n6212 gnd.n978 585
R995 gnd.n6210 gnd.n6209 585
R996 gnd.n6211 gnd.n6210 585
R997 gnd.n6208 gnd.n980 585
R998 gnd.n980 gnd.n979 585
R999 gnd.n6207 gnd.n6206 585
R1000 gnd.n6206 gnd.n6205 585
R1001 gnd.n986 gnd.n985 585
R1002 gnd.n6204 gnd.n986 585
R1003 gnd.n6202 gnd.n6201 585
R1004 gnd.n6203 gnd.n6202 585
R1005 gnd.n6200 gnd.n988 585
R1006 gnd.n988 gnd.n987 585
R1007 gnd.n6199 gnd.n6198 585
R1008 gnd.n6198 gnd.n6197 585
R1009 gnd.n994 gnd.n993 585
R1010 gnd.n6196 gnd.n994 585
R1011 gnd.n6194 gnd.n6193 585
R1012 gnd.n6195 gnd.n6194 585
R1013 gnd.n6192 gnd.n996 585
R1014 gnd.n996 gnd.n995 585
R1015 gnd.n6191 gnd.n6190 585
R1016 gnd.n6190 gnd.n6189 585
R1017 gnd.n1002 gnd.n1001 585
R1018 gnd.n6188 gnd.n1002 585
R1019 gnd.n6186 gnd.n6185 585
R1020 gnd.n6187 gnd.n6186 585
R1021 gnd.n6184 gnd.n1004 585
R1022 gnd.n1004 gnd.n1003 585
R1023 gnd.n6183 gnd.n6182 585
R1024 gnd.n6182 gnd.n6181 585
R1025 gnd.n1010 gnd.n1009 585
R1026 gnd.n6180 gnd.n1010 585
R1027 gnd.n6178 gnd.n6177 585
R1028 gnd.n6179 gnd.n6178 585
R1029 gnd.n6176 gnd.n1012 585
R1030 gnd.n1012 gnd.n1011 585
R1031 gnd.n6175 gnd.n6174 585
R1032 gnd.n6174 gnd.n6173 585
R1033 gnd.n1018 gnd.n1017 585
R1034 gnd.n6172 gnd.n1018 585
R1035 gnd.n6170 gnd.n6169 585
R1036 gnd.n6171 gnd.n6170 585
R1037 gnd.n6168 gnd.n1020 585
R1038 gnd.n1020 gnd.n1019 585
R1039 gnd.n6167 gnd.n6166 585
R1040 gnd.n6166 gnd.n6165 585
R1041 gnd.n1026 gnd.n1025 585
R1042 gnd.n6164 gnd.n1026 585
R1043 gnd.n6162 gnd.n6161 585
R1044 gnd.n6163 gnd.n6162 585
R1045 gnd.n6160 gnd.n1028 585
R1046 gnd.n1028 gnd.n1027 585
R1047 gnd.n6159 gnd.n6158 585
R1048 gnd.n6158 gnd.n6157 585
R1049 gnd.n1034 gnd.n1033 585
R1050 gnd.n6156 gnd.n1034 585
R1051 gnd.n6154 gnd.n6153 585
R1052 gnd.n6155 gnd.n6154 585
R1053 gnd.n6152 gnd.n1036 585
R1054 gnd.n1036 gnd.n1035 585
R1055 gnd.n6151 gnd.n6150 585
R1056 gnd.n6150 gnd.n6149 585
R1057 gnd.n1042 gnd.n1041 585
R1058 gnd.n6148 gnd.n1042 585
R1059 gnd.n6146 gnd.n6145 585
R1060 gnd.n6147 gnd.n6146 585
R1061 gnd.n6144 gnd.n1044 585
R1062 gnd.n1044 gnd.n1043 585
R1063 gnd.n880 gnd.n879 585
R1064 gnd.n879 gnd.n878 585
R1065 gnd.n6316 gnd.n6315 585
R1066 gnd.n6317 gnd.n6316 585
R1067 gnd.n877 gnd.n876 585
R1068 gnd.n6318 gnd.n877 585
R1069 gnd.n6321 gnd.n6320 585
R1070 gnd.n6320 gnd.n6319 585
R1071 gnd.n874 gnd.n873 585
R1072 gnd.n873 gnd.n872 585
R1073 gnd.n6326 gnd.n6325 585
R1074 gnd.n6327 gnd.n6326 585
R1075 gnd.n871 gnd.n870 585
R1076 gnd.n6328 gnd.n871 585
R1077 gnd.n6331 gnd.n6330 585
R1078 gnd.n6330 gnd.n6329 585
R1079 gnd.n868 gnd.n867 585
R1080 gnd.n867 gnd.n866 585
R1081 gnd.n6336 gnd.n6335 585
R1082 gnd.n6337 gnd.n6336 585
R1083 gnd.n865 gnd.n864 585
R1084 gnd.n6338 gnd.n865 585
R1085 gnd.n6341 gnd.n6340 585
R1086 gnd.n6340 gnd.n6339 585
R1087 gnd.n862 gnd.n861 585
R1088 gnd.n861 gnd.n860 585
R1089 gnd.n6346 gnd.n6345 585
R1090 gnd.n6347 gnd.n6346 585
R1091 gnd.n859 gnd.n858 585
R1092 gnd.n6348 gnd.n859 585
R1093 gnd.n6351 gnd.n6350 585
R1094 gnd.n6350 gnd.n6349 585
R1095 gnd.n856 gnd.n855 585
R1096 gnd.n855 gnd.n854 585
R1097 gnd.n6356 gnd.n6355 585
R1098 gnd.n6357 gnd.n6356 585
R1099 gnd.n853 gnd.n852 585
R1100 gnd.n6358 gnd.n853 585
R1101 gnd.n6361 gnd.n6360 585
R1102 gnd.n6360 gnd.n6359 585
R1103 gnd.n850 gnd.n849 585
R1104 gnd.n849 gnd.n848 585
R1105 gnd.n6366 gnd.n6365 585
R1106 gnd.n6367 gnd.n6366 585
R1107 gnd.n847 gnd.n846 585
R1108 gnd.n6368 gnd.n847 585
R1109 gnd.n6371 gnd.n6370 585
R1110 gnd.n6370 gnd.n6369 585
R1111 gnd.n844 gnd.n843 585
R1112 gnd.n843 gnd.n842 585
R1113 gnd.n6376 gnd.n6375 585
R1114 gnd.n6377 gnd.n6376 585
R1115 gnd.n841 gnd.n840 585
R1116 gnd.n6378 gnd.n841 585
R1117 gnd.n6381 gnd.n6380 585
R1118 gnd.n6380 gnd.n6379 585
R1119 gnd.n838 gnd.n837 585
R1120 gnd.n837 gnd.n836 585
R1121 gnd.n6386 gnd.n6385 585
R1122 gnd.n6387 gnd.n6386 585
R1123 gnd.n835 gnd.n834 585
R1124 gnd.n6388 gnd.n835 585
R1125 gnd.n6391 gnd.n6390 585
R1126 gnd.n6390 gnd.n6389 585
R1127 gnd.n832 gnd.n831 585
R1128 gnd.n831 gnd.n830 585
R1129 gnd.n6396 gnd.n6395 585
R1130 gnd.n6397 gnd.n6396 585
R1131 gnd.n829 gnd.n828 585
R1132 gnd.n6398 gnd.n829 585
R1133 gnd.n6401 gnd.n6400 585
R1134 gnd.n6400 gnd.n6399 585
R1135 gnd.n826 gnd.n825 585
R1136 gnd.n825 gnd.n824 585
R1137 gnd.n6406 gnd.n6405 585
R1138 gnd.n6407 gnd.n6406 585
R1139 gnd.n823 gnd.n822 585
R1140 gnd.n6408 gnd.n823 585
R1141 gnd.n6411 gnd.n6410 585
R1142 gnd.n6410 gnd.n6409 585
R1143 gnd.n820 gnd.n819 585
R1144 gnd.n819 gnd.n818 585
R1145 gnd.n6416 gnd.n6415 585
R1146 gnd.n6417 gnd.n6416 585
R1147 gnd.n817 gnd.n816 585
R1148 gnd.n6418 gnd.n817 585
R1149 gnd.n6421 gnd.n6420 585
R1150 gnd.n6420 gnd.n6419 585
R1151 gnd.n814 gnd.n813 585
R1152 gnd.n813 gnd.n812 585
R1153 gnd.n6426 gnd.n6425 585
R1154 gnd.n6427 gnd.n6426 585
R1155 gnd.n811 gnd.n810 585
R1156 gnd.n6428 gnd.n811 585
R1157 gnd.n6431 gnd.n6430 585
R1158 gnd.n6430 gnd.n6429 585
R1159 gnd.n808 gnd.n807 585
R1160 gnd.n807 gnd.n806 585
R1161 gnd.n6436 gnd.n6435 585
R1162 gnd.n6437 gnd.n6436 585
R1163 gnd.n805 gnd.n804 585
R1164 gnd.n6438 gnd.n805 585
R1165 gnd.n6441 gnd.n6440 585
R1166 gnd.n6440 gnd.n6439 585
R1167 gnd.n802 gnd.n801 585
R1168 gnd.n801 gnd.n800 585
R1169 gnd.n6446 gnd.n6445 585
R1170 gnd.n6447 gnd.n6446 585
R1171 gnd.n799 gnd.n798 585
R1172 gnd.n6448 gnd.n799 585
R1173 gnd.n6451 gnd.n6450 585
R1174 gnd.n6450 gnd.n6449 585
R1175 gnd.n796 gnd.n795 585
R1176 gnd.n795 gnd.n794 585
R1177 gnd.n6456 gnd.n6455 585
R1178 gnd.n6457 gnd.n6456 585
R1179 gnd.n793 gnd.n792 585
R1180 gnd.n6458 gnd.n793 585
R1181 gnd.n6461 gnd.n6460 585
R1182 gnd.n6460 gnd.n6459 585
R1183 gnd.n790 gnd.n789 585
R1184 gnd.n789 gnd.n788 585
R1185 gnd.n6466 gnd.n6465 585
R1186 gnd.n6467 gnd.n6466 585
R1187 gnd.n787 gnd.n786 585
R1188 gnd.n6468 gnd.n787 585
R1189 gnd.n6471 gnd.n6470 585
R1190 gnd.n6470 gnd.n6469 585
R1191 gnd.n784 gnd.n783 585
R1192 gnd.n783 gnd.n782 585
R1193 gnd.n6476 gnd.n6475 585
R1194 gnd.n6477 gnd.n6476 585
R1195 gnd.n781 gnd.n780 585
R1196 gnd.n6478 gnd.n781 585
R1197 gnd.n6481 gnd.n6480 585
R1198 gnd.n6480 gnd.n6479 585
R1199 gnd.n778 gnd.n777 585
R1200 gnd.n777 gnd.n776 585
R1201 gnd.n6486 gnd.n6485 585
R1202 gnd.n6487 gnd.n6486 585
R1203 gnd.n775 gnd.n774 585
R1204 gnd.n6488 gnd.n775 585
R1205 gnd.n6491 gnd.n6490 585
R1206 gnd.n6490 gnd.n6489 585
R1207 gnd.n772 gnd.n771 585
R1208 gnd.n771 gnd.n770 585
R1209 gnd.n6496 gnd.n6495 585
R1210 gnd.n6497 gnd.n6496 585
R1211 gnd.n769 gnd.n768 585
R1212 gnd.n6498 gnd.n769 585
R1213 gnd.n6501 gnd.n6500 585
R1214 gnd.n6500 gnd.n6499 585
R1215 gnd.n766 gnd.n765 585
R1216 gnd.n765 gnd.n764 585
R1217 gnd.n6506 gnd.n6505 585
R1218 gnd.n6507 gnd.n6506 585
R1219 gnd.n763 gnd.n762 585
R1220 gnd.n6508 gnd.n763 585
R1221 gnd.n6511 gnd.n6510 585
R1222 gnd.n6510 gnd.n6509 585
R1223 gnd.n760 gnd.n759 585
R1224 gnd.n759 gnd.n758 585
R1225 gnd.n6516 gnd.n6515 585
R1226 gnd.n6517 gnd.n6516 585
R1227 gnd.n757 gnd.n756 585
R1228 gnd.n6518 gnd.n757 585
R1229 gnd.n6521 gnd.n6520 585
R1230 gnd.n6520 gnd.n6519 585
R1231 gnd.n754 gnd.n753 585
R1232 gnd.n753 gnd.n752 585
R1233 gnd.n6526 gnd.n6525 585
R1234 gnd.n6527 gnd.n6526 585
R1235 gnd.n751 gnd.n750 585
R1236 gnd.n6528 gnd.n751 585
R1237 gnd.n6531 gnd.n6530 585
R1238 gnd.n6530 gnd.n6529 585
R1239 gnd.n748 gnd.n747 585
R1240 gnd.n747 gnd.n746 585
R1241 gnd.n6536 gnd.n6535 585
R1242 gnd.n6537 gnd.n6536 585
R1243 gnd.n745 gnd.n744 585
R1244 gnd.n6538 gnd.n745 585
R1245 gnd.n6541 gnd.n6540 585
R1246 gnd.n6540 gnd.n6539 585
R1247 gnd.n742 gnd.n741 585
R1248 gnd.n741 gnd.n740 585
R1249 gnd.n6546 gnd.n6545 585
R1250 gnd.n6547 gnd.n6546 585
R1251 gnd.n739 gnd.n738 585
R1252 gnd.n6548 gnd.n739 585
R1253 gnd.n6551 gnd.n6550 585
R1254 gnd.n6550 gnd.n6549 585
R1255 gnd.n736 gnd.n735 585
R1256 gnd.n735 gnd.n734 585
R1257 gnd.n6556 gnd.n6555 585
R1258 gnd.n6557 gnd.n6556 585
R1259 gnd.n733 gnd.n732 585
R1260 gnd.n6558 gnd.n733 585
R1261 gnd.n6561 gnd.n6560 585
R1262 gnd.n6560 gnd.n6559 585
R1263 gnd.n730 gnd.n729 585
R1264 gnd.n729 gnd.n728 585
R1265 gnd.n6566 gnd.n6565 585
R1266 gnd.n6567 gnd.n6566 585
R1267 gnd.n727 gnd.n726 585
R1268 gnd.n6568 gnd.n727 585
R1269 gnd.n6571 gnd.n6570 585
R1270 gnd.n6570 gnd.n6569 585
R1271 gnd.n724 gnd.n723 585
R1272 gnd.n723 gnd.n722 585
R1273 gnd.n6576 gnd.n6575 585
R1274 gnd.n6577 gnd.n6576 585
R1275 gnd.n721 gnd.n720 585
R1276 gnd.n6578 gnd.n721 585
R1277 gnd.n6581 gnd.n6580 585
R1278 gnd.n6580 gnd.n6579 585
R1279 gnd.n718 gnd.n717 585
R1280 gnd.n717 gnd.n716 585
R1281 gnd.n6586 gnd.n6585 585
R1282 gnd.n6587 gnd.n6586 585
R1283 gnd.n715 gnd.n714 585
R1284 gnd.n6588 gnd.n715 585
R1285 gnd.n6591 gnd.n6590 585
R1286 gnd.n6590 gnd.n6589 585
R1287 gnd.n712 gnd.n711 585
R1288 gnd.n711 gnd.n710 585
R1289 gnd.n6596 gnd.n6595 585
R1290 gnd.n6597 gnd.n6596 585
R1291 gnd.n709 gnd.n708 585
R1292 gnd.n6598 gnd.n709 585
R1293 gnd.n6601 gnd.n6600 585
R1294 gnd.n6600 gnd.n6599 585
R1295 gnd.n706 gnd.n705 585
R1296 gnd.n705 gnd.n704 585
R1297 gnd.n6606 gnd.n6605 585
R1298 gnd.n6607 gnd.n6606 585
R1299 gnd.n703 gnd.n702 585
R1300 gnd.n6608 gnd.n703 585
R1301 gnd.n6611 gnd.n6610 585
R1302 gnd.n6610 gnd.n6609 585
R1303 gnd.n700 gnd.n699 585
R1304 gnd.n699 gnd.n698 585
R1305 gnd.n6616 gnd.n6615 585
R1306 gnd.n6617 gnd.n6616 585
R1307 gnd.n697 gnd.n696 585
R1308 gnd.n6618 gnd.n697 585
R1309 gnd.n6621 gnd.n6620 585
R1310 gnd.n6620 gnd.n6619 585
R1311 gnd.n694 gnd.n693 585
R1312 gnd.n693 gnd.n692 585
R1313 gnd.n6627 gnd.n6626 585
R1314 gnd.n6628 gnd.n6627 585
R1315 gnd.n691 gnd.n690 585
R1316 gnd.n6629 gnd.n691 585
R1317 gnd.n6632 gnd.n6631 585
R1318 gnd.n6631 gnd.n6630 585
R1319 gnd.n6633 gnd.n688 585
R1320 gnd.n688 gnd.n687 585
R1321 gnd.n563 gnd.n562 585
R1322 gnd.n6840 gnd.n562 585
R1323 gnd.n6843 gnd.n6842 585
R1324 gnd.n6842 gnd.n6841 585
R1325 gnd.n566 gnd.n565 585
R1326 gnd.n6839 gnd.n566 585
R1327 gnd.n6837 gnd.n6836 585
R1328 gnd.n6838 gnd.n6837 585
R1329 gnd.n569 gnd.n568 585
R1330 gnd.n568 gnd.n567 585
R1331 gnd.n6832 gnd.n6831 585
R1332 gnd.n6831 gnd.n6830 585
R1333 gnd.n572 gnd.n571 585
R1334 gnd.n6829 gnd.n572 585
R1335 gnd.n6827 gnd.n6826 585
R1336 gnd.n6828 gnd.n6827 585
R1337 gnd.n575 gnd.n574 585
R1338 gnd.n574 gnd.n573 585
R1339 gnd.n6822 gnd.n6821 585
R1340 gnd.n6821 gnd.n6820 585
R1341 gnd.n578 gnd.n577 585
R1342 gnd.n6819 gnd.n578 585
R1343 gnd.n6817 gnd.n6816 585
R1344 gnd.n6818 gnd.n6817 585
R1345 gnd.n581 gnd.n580 585
R1346 gnd.n580 gnd.n579 585
R1347 gnd.n6812 gnd.n6811 585
R1348 gnd.n6811 gnd.n6810 585
R1349 gnd.n584 gnd.n583 585
R1350 gnd.n6809 gnd.n584 585
R1351 gnd.n6807 gnd.n6806 585
R1352 gnd.n6808 gnd.n6807 585
R1353 gnd.n587 gnd.n586 585
R1354 gnd.n586 gnd.n585 585
R1355 gnd.n6802 gnd.n6801 585
R1356 gnd.n6801 gnd.n6800 585
R1357 gnd.n590 gnd.n589 585
R1358 gnd.n6799 gnd.n590 585
R1359 gnd.n6797 gnd.n6796 585
R1360 gnd.n6798 gnd.n6797 585
R1361 gnd.n593 gnd.n592 585
R1362 gnd.n592 gnd.n591 585
R1363 gnd.n6792 gnd.n6791 585
R1364 gnd.n6791 gnd.n6790 585
R1365 gnd.n596 gnd.n595 585
R1366 gnd.n6789 gnd.n596 585
R1367 gnd.n6787 gnd.n6786 585
R1368 gnd.n6788 gnd.n6787 585
R1369 gnd.n599 gnd.n598 585
R1370 gnd.n598 gnd.n597 585
R1371 gnd.n6782 gnd.n6781 585
R1372 gnd.n6781 gnd.n6780 585
R1373 gnd.n602 gnd.n601 585
R1374 gnd.n6779 gnd.n602 585
R1375 gnd.n6777 gnd.n6776 585
R1376 gnd.n6778 gnd.n6777 585
R1377 gnd.n605 gnd.n604 585
R1378 gnd.n604 gnd.n603 585
R1379 gnd.n6772 gnd.n6771 585
R1380 gnd.n6771 gnd.n6770 585
R1381 gnd.n608 gnd.n607 585
R1382 gnd.n6769 gnd.n608 585
R1383 gnd.n6767 gnd.n6766 585
R1384 gnd.n6768 gnd.n6767 585
R1385 gnd.n611 gnd.n610 585
R1386 gnd.n610 gnd.n609 585
R1387 gnd.n6762 gnd.n6761 585
R1388 gnd.n6761 gnd.n6760 585
R1389 gnd.n614 gnd.n613 585
R1390 gnd.n6759 gnd.n614 585
R1391 gnd.n6757 gnd.n6756 585
R1392 gnd.n6758 gnd.n6757 585
R1393 gnd.n617 gnd.n616 585
R1394 gnd.n616 gnd.n615 585
R1395 gnd.n6752 gnd.n6751 585
R1396 gnd.n6751 gnd.n6750 585
R1397 gnd.n620 gnd.n619 585
R1398 gnd.n6749 gnd.n620 585
R1399 gnd.n6747 gnd.n6746 585
R1400 gnd.n6748 gnd.n6747 585
R1401 gnd.n623 gnd.n622 585
R1402 gnd.n622 gnd.n621 585
R1403 gnd.n6742 gnd.n6741 585
R1404 gnd.n6741 gnd.n6740 585
R1405 gnd.n626 gnd.n625 585
R1406 gnd.n6739 gnd.n626 585
R1407 gnd.n6737 gnd.n6736 585
R1408 gnd.n6738 gnd.n6737 585
R1409 gnd.n629 gnd.n628 585
R1410 gnd.n628 gnd.n627 585
R1411 gnd.n6732 gnd.n6731 585
R1412 gnd.n6731 gnd.n6730 585
R1413 gnd.n632 gnd.n631 585
R1414 gnd.n6729 gnd.n632 585
R1415 gnd.n6727 gnd.n6726 585
R1416 gnd.n6728 gnd.n6727 585
R1417 gnd.n635 gnd.n634 585
R1418 gnd.n634 gnd.n633 585
R1419 gnd.n6722 gnd.n6721 585
R1420 gnd.n6721 gnd.n6720 585
R1421 gnd.n638 gnd.n637 585
R1422 gnd.n6719 gnd.n638 585
R1423 gnd.n6717 gnd.n6716 585
R1424 gnd.n6718 gnd.n6717 585
R1425 gnd.n641 gnd.n640 585
R1426 gnd.n640 gnd.n639 585
R1427 gnd.n6712 gnd.n6711 585
R1428 gnd.n6711 gnd.n6710 585
R1429 gnd.n644 gnd.n643 585
R1430 gnd.n6709 gnd.n644 585
R1431 gnd.n6707 gnd.n6706 585
R1432 gnd.n6708 gnd.n6707 585
R1433 gnd.n647 gnd.n646 585
R1434 gnd.n646 gnd.n645 585
R1435 gnd.n6702 gnd.n6701 585
R1436 gnd.n6701 gnd.n6700 585
R1437 gnd.n650 gnd.n649 585
R1438 gnd.n6699 gnd.n650 585
R1439 gnd.n6697 gnd.n6696 585
R1440 gnd.n6698 gnd.n6697 585
R1441 gnd.n653 gnd.n652 585
R1442 gnd.n652 gnd.n651 585
R1443 gnd.n6692 gnd.n6691 585
R1444 gnd.n6691 gnd.n6690 585
R1445 gnd.n656 gnd.n655 585
R1446 gnd.n6689 gnd.n656 585
R1447 gnd.n6687 gnd.n6686 585
R1448 gnd.n6688 gnd.n6687 585
R1449 gnd.n659 gnd.n658 585
R1450 gnd.n658 gnd.n657 585
R1451 gnd.n6682 gnd.n6681 585
R1452 gnd.n6681 gnd.n6680 585
R1453 gnd.n662 gnd.n661 585
R1454 gnd.n6679 gnd.n662 585
R1455 gnd.n6677 gnd.n6676 585
R1456 gnd.n6678 gnd.n6677 585
R1457 gnd.n665 gnd.n664 585
R1458 gnd.n664 gnd.n663 585
R1459 gnd.n6672 gnd.n6671 585
R1460 gnd.n6671 gnd.n6670 585
R1461 gnd.n668 gnd.n667 585
R1462 gnd.n6669 gnd.n668 585
R1463 gnd.n6667 gnd.n6666 585
R1464 gnd.n6668 gnd.n6667 585
R1465 gnd.n671 gnd.n670 585
R1466 gnd.n670 gnd.n669 585
R1467 gnd.n6662 gnd.n6661 585
R1468 gnd.n6661 gnd.n6660 585
R1469 gnd.n674 gnd.n673 585
R1470 gnd.n6659 gnd.n674 585
R1471 gnd.n6657 gnd.n6656 585
R1472 gnd.n6658 gnd.n6657 585
R1473 gnd.n677 gnd.n676 585
R1474 gnd.n676 gnd.n675 585
R1475 gnd.n6652 gnd.n6651 585
R1476 gnd.n6651 gnd.n6650 585
R1477 gnd.n680 gnd.n679 585
R1478 gnd.n6649 gnd.n680 585
R1479 gnd.n6647 gnd.n6646 585
R1480 gnd.n6648 gnd.n6647 585
R1481 gnd.n683 gnd.n682 585
R1482 gnd.n682 gnd.n681 585
R1483 gnd.n6642 gnd.n6641 585
R1484 gnd.n6641 gnd.n6640 585
R1485 gnd.n686 gnd.n685 585
R1486 gnd.n6639 gnd.n686 585
R1487 gnd.n6637 gnd.n6636 585
R1488 gnd.n6638 gnd.n6637 585
R1489 gnd.n1133 gnd.n1132 585
R1490 gnd.n4714 gnd.n1133 585
R1491 gnd.n6094 gnd.n6093 585
R1492 gnd.n6093 gnd.n6092 585
R1493 gnd.n6095 gnd.n1128 585
R1494 gnd.n4677 gnd.n1128 585
R1495 gnd.n6097 gnd.n6096 585
R1496 gnd.n6098 gnd.n6097 585
R1497 gnd.n1112 gnd.n1111 585
R1498 gnd.n4437 gnd.n1112 585
R1499 gnd.n6106 gnd.n6105 585
R1500 gnd.n6105 gnd.n6104 585
R1501 gnd.n6107 gnd.n1107 585
R1502 gnd.n4690 gnd.n1107 585
R1503 gnd.n6109 gnd.n6108 585
R1504 gnd.n6110 gnd.n6109 585
R1505 gnd.n1093 gnd.n1092 585
R1506 gnd.n4430 gnd.n1093 585
R1507 gnd.n6118 gnd.n6117 585
R1508 gnd.n6117 gnd.n6116 585
R1509 gnd.n6119 gnd.n1088 585
R1510 gnd.n4422 gnd.n1088 585
R1511 gnd.n6121 gnd.n6120 585
R1512 gnd.n6122 gnd.n6121 585
R1513 gnd.n1072 gnd.n1071 585
R1514 gnd.n4387 gnd.n1072 585
R1515 gnd.n6130 gnd.n6129 585
R1516 gnd.n6129 gnd.n6128 585
R1517 gnd.n6131 gnd.n1066 585
R1518 gnd.n4395 gnd.n1066 585
R1519 gnd.n6133 gnd.n6132 585
R1520 gnd.n6134 gnd.n6133 585
R1521 gnd.n1067 gnd.n1065 585
R1522 gnd.n4376 gnd.n1065 585
R1523 gnd.n4352 gnd.n1054 585
R1524 gnd.n6140 gnd.n1054 585
R1525 gnd.n4354 gnd.n4353 585
R1526 gnd.n4353 gnd.n1050 585
R1527 gnd.n4355 gnd.n2335 585
R1528 gnd.n4367 gnd.n2335 585
R1529 gnd.n4356 gnd.n2344 585
R1530 gnd.n2344 gnd.n2342 585
R1531 gnd.n4358 gnd.n4357 585
R1532 gnd.n4359 gnd.n4358 585
R1533 gnd.n2345 gnd.n2343 585
R1534 gnd.n2343 gnd.n2339 585
R1535 gnd.n4328 gnd.n2354 585
R1536 gnd.n4340 gnd.n2354 585
R1537 gnd.n4329 gnd.n2362 585
R1538 gnd.n2362 gnd.n2352 585
R1539 gnd.n4331 gnd.n4330 585
R1540 gnd.n4332 gnd.n4331 585
R1541 gnd.n2363 gnd.n2361 585
R1542 gnd.n2361 gnd.n2358 585
R1543 gnd.n4307 gnd.n2369 585
R1544 gnd.n4320 gnd.n2369 585
R1545 gnd.n4308 gnd.n2380 585
R1546 gnd.n2380 gnd.n2378 585
R1547 gnd.n4310 gnd.n4309 585
R1548 gnd.n4311 gnd.n4310 585
R1549 gnd.n2381 gnd.n2379 585
R1550 gnd.n2379 gnd.n2375 585
R1551 gnd.n4287 gnd.n2388 585
R1552 gnd.n4299 gnd.n2388 585
R1553 gnd.n4288 gnd.n2398 585
R1554 gnd.n2398 gnd.n2386 585
R1555 gnd.n4290 gnd.n4289 585
R1556 gnd.n4291 gnd.n4290 585
R1557 gnd.n2399 gnd.n2397 585
R1558 gnd.n2397 gnd.n2394 585
R1559 gnd.n4267 gnd.n2405 585
R1560 gnd.n4279 gnd.n2405 585
R1561 gnd.n4268 gnd.n2416 585
R1562 gnd.n2416 gnd.n2414 585
R1563 gnd.n4270 gnd.n4269 585
R1564 gnd.n4271 gnd.n4270 585
R1565 gnd.n2417 gnd.n2415 585
R1566 gnd.n2415 gnd.n2411 585
R1567 gnd.n2438 gnd.n2424 585
R1568 gnd.n4259 gnd.n2424 585
R1569 gnd.n2436 gnd.n2434 585
R1570 gnd.n2434 gnd.n2422 585
R1571 gnd.n4250 gnd.n4249 585
R1572 gnd.n4251 gnd.n4250 585
R1573 gnd.n2435 gnd.n2433 585
R1574 gnd.n2433 gnd.n2430 585
R1575 gnd.n4121 gnd.n4120 585
R1576 gnd.n4119 gnd.n4118 585
R1577 gnd.n4117 gnd.n4116 585
R1578 gnd.n4115 gnd.n4114 585
R1579 gnd.n4113 gnd.n4112 585
R1580 gnd.n4111 gnd.n4110 585
R1581 gnd.n4109 gnd.n4108 585
R1582 gnd.n4107 gnd.n4106 585
R1583 gnd.n4105 gnd.n4104 585
R1584 gnd.n4103 gnd.n4102 585
R1585 gnd.n4101 gnd.n4100 585
R1586 gnd.n4099 gnd.n4098 585
R1587 gnd.n4097 gnd.n4096 585
R1588 gnd.n4095 gnd.n4094 585
R1589 gnd.n4093 gnd.n4092 585
R1590 gnd.n4091 gnd.n4090 585
R1591 gnd.n4089 gnd.n4088 585
R1592 gnd.n4026 gnd.n4023 585
R1593 gnd.n4084 gnd.n3942 585
R1594 gnd.n4241 gnd.n3942 585
R1595 gnd.n4717 gnd.n4716 585
R1596 gnd.n4514 gnd.n2294 585
R1597 gnd.n4526 gnd.n4515 585
R1598 gnd.n4527 gnd.n4513 585
R1599 gnd.n4512 gnd.n4504 585
R1600 gnd.n4534 gnd.n4503 585
R1601 gnd.n4535 gnd.n4502 585
R1602 gnd.n4496 gnd.n4495 585
R1603 gnd.n4542 gnd.n4494 585
R1604 gnd.n4543 gnd.n4493 585
R1605 gnd.n4492 gnd.n4484 585
R1606 gnd.n4550 gnd.n4483 585
R1607 gnd.n4551 gnd.n4482 585
R1608 gnd.n4476 gnd.n4475 585
R1609 gnd.n4558 gnd.n4474 585
R1610 gnd.n4559 gnd.n4473 585
R1611 gnd.n4472 gnd.n4464 585
R1612 gnd.n4566 gnd.n4463 585
R1613 gnd.n4567 gnd.n1145 585
R1614 gnd.n6084 gnd.n1145 585
R1615 gnd.n4715 gnd.n2295 585
R1616 gnd.n4715 gnd.n4714 585
R1617 gnd.n4679 gnd.n1136 585
R1618 gnd.n6092 gnd.n1136 585
R1619 gnd.n4682 gnd.n4678 585
R1620 gnd.n4678 gnd.n4677 585
R1621 gnd.n4683 gnd.n1126 585
R1622 gnd.n6098 gnd.n1126 585
R1623 gnd.n4684 gnd.n2312 585
R1624 gnd.n4437 gnd.n2312 585
R1625 gnd.n2309 gnd.n1115 585
R1626 gnd.n6104 gnd.n1115 585
R1627 gnd.n4689 gnd.n4688 585
R1628 gnd.n4690 gnd.n4689 585
R1629 gnd.n2308 gnd.n1106 585
R1630 gnd.n6110 gnd.n1106 585
R1631 gnd.n4429 gnd.n4428 585
R1632 gnd.n4430 gnd.n4429 585
R1633 gnd.n2315 gnd.n1095 585
R1634 gnd.n6116 gnd.n1095 585
R1635 gnd.n4424 gnd.n4423 585
R1636 gnd.n4423 gnd.n4422 585
R1637 gnd.n2317 gnd.n1086 585
R1638 gnd.n6122 gnd.n1086 585
R1639 gnd.n4389 gnd.n4388 585
R1640 gnd.n4388 gnd.n4387 585
R1641 gnd.n2326 gnd.n1075 585
R1642 gnd.n6128 gnd.n1075 585
R1643 gnd.n4394 gnd.n4393 585
R1644 gnd.n4395 gnd.n4394 585
R1645 gnd.n2325 gnd.n1064 585
R1646 gnd.n6134 gnd.n1064 585
R1647 gnd.n4375 gnd.n4374 585
R1648 gnd.n4376 gnd.n4375 585
R1649 gnd.n2330 gnd.n1052 585
R1650 gnd.n6140 gnd.n1052 585
R1651 gnd.n4370 gnd.n4369 585
R1652 gnd.n4369 gnd.n1050 585
R1653 gnd.n4368 gnd.n2332 585
R1654 gnd.n4368 gnd.n4367 585
R1655 gnd.n4047 gnd.n2333 585
R1656 gnd.n2342 gnd.n2333 585
R1657 gnd.n4050 gnd.n2341 585
R1658 gnd.n4359 gnd.n2341 585
R1659 gnd.n4052 gnd.n4051 585
R1660 gnd.n4051 gnd.n2339 585
R1661 gnd.n4053 gnd.n2353 585
R1662 gnd.n4340 gnd.n2353 585
R1663 gnd.n4055 gnd.n4054 585
R1664 gnd.n4054 gnd.n2352 585
R1665 gnd.n4056 gnd.n2360 585
R1666 gnd.n4332 gnd.n2360 585
R1667 gnd.n4058 gnd.n4057 585
R1668 gnd.n4057 gnd.n2358 585
R1669 gnd.n4059 gnd.n2368 585
R1670 gnd.n4320 gnd.n2368 585
R1671 gnd.n4061 gnd.n4060 585
R1672 gnd.n4060 gnd.n2378 585
R1673 gnd.n4062 gnd.n2377 585
R1674 gnd.n4311 gnd.n2377 585
R1675 gnd.n4064 gnd.n4063 585
R1676 gnd.n4063 gnd.n2375 585
R1677 gnd.n4065 gnd.n2387 585
R1678 gnd.n4299 gnd.n2387 585
R1679 gnd.n4067 gnd.n4066 585
R1680 gnd.n4066 gnd.n2386 585
R1681 gnd.n4068 gnd.n2396 585
R1682 gnd.n4291 gnd.n2396 585
R1683 gnd.n4070 gnd.n4069 585
R1684 gnd.n4069 gnd.n2394 585
R1685 gnd.n4071 gnd.n2404 585
R1686 gnd.n4279 gnd.n2404 585
R1687 gnd.n4073 gnd.n4072 585
R1688 gnd.n4072 gnd.n2414 585
R1689 gnd.n4074 gnd.n2413 585
R1690 gnd.n4271 gnd.n2413 585
R1691 gnd.n4076 gnd.n4075 585
R1692 gnd.n4075 gnd.n2411 585
R1693 gnd.n4077 gnd.n2423 585
R1694 gnd.n4259 gnd.n2423 585
R1695 gnd.n4079 gnd.n4078 585
R1696 gnd.n4078 gnd.n2422 585
R1697 gnd.n4080 gnd.n2432 585
R1698 gnd.n4251 gnd.n2432 585
R1699 gnd.n4082 gnd.n4081 585
R1700 gnd.n4081 gnd.n2430 585
R1701 gnd.n3813 gnd.n3812 585
R1702 gnd.n3814 gnd.n3813 585
R1703 gnd.n2519 gnd.n2518 585
R1704 gnd.n2525 gnd.n2518 585
R1705 gnd.n3788 gnd.n2537 585
R1706 gnd.n2537 gnd.n2524 585
R1707 gnd.n3790 gnd.n3789 585
R1708 gnd.n3791 gnd.n3790 585
R1709 gnd.n2538 gnd.n2536 585
R1710 gnd.n2536 gnd.n2532 585
R1711 gnd.n3522 gnd.n3521 585
R1712 gnd.n3521 gnd.n3520 585
R1713 gnd.n2543 gnd.n2542 585
R1714 gnd.n3490 gnd.n2543 585
R1715 gnd.n3510 gnd.n3509 585
R1716 gnd.n3509 gnd.n3508 585
R1717 gnd.n2550 gnd.n2549 585
R1718 gnd.n3496 gnd.n2550 585
R1719 gnd.n3466 gnd.n2570 585
R1720 gnd.n2570 gnd.n2569 585
R1721 gnd.n3468 gnd.n3467 585
R1722 gnd.n3469 gnd.n3468 585
R1723 gnd.n2571 gnd.n2568 585
R1724 gnd.n2579 gnd.n2568 585
R1725 gnd.n3444 gnd.n2591 585
R1726 gnd.n2591 gnd.n2578 585
R1727 gnd.n3446 gnd.n3445 585
R1728 gnd.n3447 gnd.n3446 585
R1729 gnd.n2592 gnd.n2590 585
R1730 gnd.n2590 gnd.n2586 585
R1731 gnd.n3432 gnd.n3431 585
R1732 gnd.n3431 gnd.n3430 585
R1733 gnd.n2597 gnd.n2596 585
R1734 gnd.n2607 gnd.n2597 585
R1735 gnd.n3421 gnd.n3420 585
R1736 gnd.n3420 gnd.n3419 585
R1737 gnd.n2604 gnd.n2603 585
R1738 gnd.n3407 gnd.n2604 585
R1739 gnd.n3381 gnd.n2625 585
R1740 gnd.n2625 gnd.n2614 585
R1741 gnd.n3383 gnd.n3382 585
R1742 gnd.n3384 gnd.n3383 585
R1743 gnd.n2626 gnd.n2624 585
R1744 gnd.n2634 gnd.n2624 585
R1745 gnd.n3359 gnd.n2646 585
R1746 gnd.n2646 gnd.n2633 585
R1747 gnd.n3361 gnd.n3360 585
R1748 gnd.n3362 gnd.n3361 585
R1749 gnd.n2647 gnd.n2645 585
R1750 gnd.n2645 gnd.n2641 585
R1751 gnd.n3347 gnd.n3346 585
R1752 gnd.n3346 gnd.n3345 585
R1753 gnd.n2652 gnd.n2651 585
R1754 gnd.n2661 gnd.n2652 585
R1755 gnd.n3336 gnd.n3335 585
R1756 gnd.n3335 gnd.n3334 585
R1757 gnd.n2659 gnd.n2658 585
R1758 gnd.n3322 gnd.n2659 585
R1759 gnd.n2760 gnd.n2759 585
R1760 gnd.n2760 gnd.n2668 585
R1761 gnd.n3279 gnd.n3278 585
R1762 gnd.n3278 gnd.n3277 585
R1763 gnd.n3280 gnd.n2754 585
R1764 gnd.n2765 gnd.n2754 585
R1765 gnd.n3282 gnd.n3281 585
R1766 gnd.n3283 gnd.n3282 585
R1767 gnd.n2755 gnd.n2753 585
R1768 gnd.n2778 gnd.n2753 585
R1769 gnd.n2738 gnd.n2737 585
R1770 gnd.n2741 gnd.n2738 585
R1771 gnd.n3293 gnd.n3292 585
R1772 gnd.n3292 gnd.n3291 585
R1773 gnd.n3294 gnd.n2732 585
R1774 gnd.n3253 gnd.n2732 585
R1775 gnd.n3296 gnd.n3295 585
R1776 gnd.n3297 gnd.n3296 585
R1777 gnd.n2733 gnd.n2731 585
R1778 gnd.n2792 gnd.n2731 585
R1779 gnd.n3245 gnd.n3244 585
R1780 gnd.n3244 gnd.n3243 585
R1781 gnd.n2789 gnd.n2788 585
R1782 gnd.n3227 gnd.n2789 585
R1783 gnd.n3214 gnd.n2808 585
R1784 gnd.n2808 gnd.n2807 585
R1785 gnd.n3216 gnd.n3215 585
R1786 gnd.n3217 gnd.n3216 585
R1787 gnd.n2809 gnd.n2806 585
R1788 gnd.n2815 gnd.n2806 585
R1789 gnd.n3195 gnd.n3194 585
R1790 gnd.n3196 gnd.n3195 585
R1791 gnd.n2826 gnd.n2825 585
R1792 gnd.n2825 gnd.n2821 585
R1793 gnd.n3185 gnd.n3184 585
R1794 gnd.n3186 gnd.n3185 585
R1795 gnd.n2836 gnd.n2835 585
R1796 gnd.n2841 gnd.n2835 585
R1797 gnd.n3163 gnd.n2854 585
R1798 gnd.n2854 gnd.n2840 585
R1799 gnd.n3165 gnd.n3164 585
R1800 gnd.n3166 gnd.n3165 585
R1801 gnd.n2855 gnd.n2853 585
R1802 gnd.n2853 gnd.n2849 585
R1803 gnd.n3154 gnd.n3153 585
R1804 gnd.n3155 gnd.n3154 585
R1805 gnd.n2862 gnd.n2861 585
R1806 gnd.n2866 gnd.n2861 585
R1807 gnd.n3131 gnd.n2883 585
R1808 gnd.n2883 gnd.n2865 585
R1809 gnd.n3133 gnd.n3132 585
R1810 gnd.n3134 gnd.n3133 585
R1811 gnd.n2884 gnd.n2882 585
R1812 gnd.n2882 gnd.n2873 585
R1813 gnd.n3126 gnd.n3125 585
R1814 gnd.n3125 gnd.n3124 585
R1815 gnd.n2931 gnd.n2930 585
R1816 gnd.n2932 gnd.n2931 585
R1817 gnd.n3085 gnd.n3084 585
R1818 gnd.n3086 gnd.n3085 585
R1819 gnd.n2941 gnd.n2940 585
R1820 gnd.n2940 gnd.n2939 585
R1821 gnd.n3080 gnd.n3079 585
R1822 gnd.n3079 gnd.n3078 585
R1823 gnd.n2944 gnd.n2943 585
R1824 gnd.n2945 gnd.n2944 585
R1825 gnd.n3069 gnd.n3068 585
R1826 gnd.n3070 gnd.n3069 585
R1827 gnd.n2952 gnd.n2951 585
R1828 gnd.n3061 gnd.n2951 585
R1829 gnd.n3064 gnd.n3063 585
R1830 gnd.n3063 gnd.n3062 585
R1831 gnd.n2955 gnd.n2954 585
R1832 gnd.n2956 gnd.n2955 585
R1833 gnd.n3050 gnd.n3049 585
R1834 gnd.n3048 gnd.n2974 585
R1835 gnd.n3047 gnd.n2973 585
R1836 gnd.n3052 gnd.n2973 585
R1837 gnd.n3046 gnd.n3045 585
R1838 gnd.n3044 gnd.n3043 585
R1839 gnd.n3042 gnd.n3041 585
R1840 gnd.n3040 gnd.n3039 585
R1841 gnd.n3038 gnd.n3037 585
R1842 gnd.n3036 gnd.n3035 585
R1843 gnd.n3034 gnd.n3033 585
R1844 gnd.n3032 gnd.n3031 585
R1845 gnd.n3030 gnd.n3029 585
R1846 gnd.n3028 gnd.n3027 585
R1847 gnd.n3026 gnd.n3025 585
R1848 gnd.n3024 gnd.n3023 585
R1849 gnd.n3022 gnd.n3021 585
R1850 gnd.n3020 gnd.n3019 585
R1851 gnd.n3018 gnd.n3017 585
R1852 gnd.n3016 gnd.n3015 585
R1853 gnd.n3014 gnd.n3013 585
R1854 gnd.n3012 gnd.n3011 585
R1855 gnd.n3010 gnd.n3009 585
R1856 gnd.n3008 gnd.n3007 585
R1857 gnd.n3006 gnd.n3005 585
R1858 gnd.n3004 gnd.n3003 585
R1859 gnd.n2961 gnd.n2960 585
R1860 gnd.n3055 gnd.n3054 585
R1861 gnd.n3817 gnd.n3816 585
R1862 gnd.n3819 gnd.n3818 585
R1863 gnd.n3821 gnd.n3820 585
R1864 gnd.n3823 gnd.n3822 585
R1865 gnd.n3825 gnd.n3824 585
R1866 gnd.n3827 gnd.n3826 585
R1867 gnd.n3829 gnd.n3828 585
R1868 gnd.n3831 gnd.n3830 585
R1869 gnd.n3833 gnd.n3832 585
R1870 gnd.n3835 gnd.n3834 585
R1871 gnd.n3837 gnd.n3836 585
R1872 gnd.n3839 gnd.n3838 585
R1873 gnd.n3841 gnd.n3840 585
R1874 gnd.n3843 gnd.n3842 585
R1875 gnd.n3845 gnd.n3844 585
R1876 gnd.n3847 gnd.n3846 585
R1877 gnd.n3849 gnd.n3848 585
R1878 gnd.n3851 gnd.n3850 585
R1879 gnd.n3853 gnd.n3852 585
R1880 gnd.n3855 gnd.n3854 585
R1881 gnd.n3857 gnd.n3856 585
R1882 gnd.n3859 gnd.n3858 585
R1883 gnd.n3861 gnd.n3860 585
R1884 gnd.n3863 gnd.n3862 585
R1885 gnd.n3865 gnd.n3864 585
R1886 gnd.n3866 gnd.n2486 585
R1887 gnd.n3867 gnd.n2444 585
R1888 gnd.n3905 gnd.n2444 585
R1889 gnd.n3815 gnd.n2516 585
R1890 gnd.n3815 gnd.n3814 585
R1891 gnd.n3483 gnd.n2515 585
R1892 gnd.n2525 gnd.n2515 585
R1893 gnd.n3485 gnd.n3484 585
R1894 gnd.n3484 gnd.n2524 585
R1895 gnd.n3486 gnd.n2534 585
R1896 gnd.n3791 gnd.n2534 585
R1897 gnd.n3488 gnd.n3487 585
R1898 gnd.n3487 gnd.n2532 585
R1899 gnd.n3489 gnd.n2545 585
R1900 gnd.n3520 gnd.n2545 585
R1901 gnd.n3492 gnd.n3491 585
R1902 gnd.n3491 gnd.n3490 585
R1903 gnd.n3493 gnd.n2552 585
R1904 gnd.n3508 gnd.n2552 585
R1905 gnd.n3495 gnd.n3494 585
R1906 gnd.n3496 gnd.n3495 585
R1907 gnd.n2562 gnd.n2561 585
R1908 gnd.n2569 gnd.n2561 585
R1909 gnd.n3471 gnd.n3470 585
R1910 gnd.n3470 gnd.n3469 585
R1911 gnd.n2565 gnd.n2564 585
R1912 gnd.n2579 gnd.n2565 585
R1913 gnd.n3397 gnd.n3396 585
R1914 gnd.n3396 gnd.n2578 585
R1915 gnd.n3398 gnd.n2588 585
R1916 gnd.n3447 gnd.n2588 585
R1917 gnd.n3400 gnd.n3399 585
R1918 gnd.n3399 gnd.n2586 585
R1919 gnd.n3401 gnd.n2599 585
R1920 gnd.n3430 gnd.n2599 585
R1921 gnd.n3403 gnd.n3402 585
R1922 gnd.n3402 gnd.n2607 585
R1923 gnd.n3404 gnd.n2606 585
R1924 gnd.n3419 gnd.n2606 585
R1925 gnd.n3406 gnd.n3405 585
R1926 gnd.n3407 gnd.n3406 585
R1927 gnd.n2618 gnd.n2617 585
R1928 gnd.n2617 gnd.n2614 585
R1929 gnd.n3386 gnd.n3385 585
R1930 gnd.n3385 gnd.n3384 585
R1931 gnd.n2621 gnd.n2620 585
R1932 gnd.n2634 gnd.n2621 585
R1933 gnd.n3310 gnd.n3309 585
R1934 gnd.n3309 gnd.n2633 585
R1935 gnd.n3311 gnd.n2643 585
R1936 gnd.n3362 gnd.n2643 585
R1937 gnd.n3313 gnd.n3312 585
R1938 gnd.n3312 gnd.n2641 585
R1939 gnd.n3314 gnd.n2654 585
R1940 gnd.n3345 gnd.n2654 585
R1941 gnd.n3316 gnd.n3315 585
R1942 gnd.n3315 gnd.n2661 585
R1943 gnd.n3317 gnd.n2660 585
R1944 gnd.n3334 gnd.n2660 585
R1945 gnd.n3319 gnd.n3318 585
R1946 gnd.n3322 gnd.n3319 585
R1947 gnd.n2671 gnd.n2670 585
R1948 gnd.n2670 gnd.n2668 585
R1949 gnd.n2762 gnd.n2761 585
R1950 gnd.n3277 gnd.n2761 585
R1951 gnd.n2764 gnd.n2763 585
R1952 gnd.n2765 gnd.n2764 585
R1953 gnd.n2775 gnd.n2751 585
R1954 gnd.n3283 gnd.n2751 585
R1955 gnd.n2777 gnd.n2776 585
R1956 gnd.n2778 gnd.n2777 585
R1957 gnd.n2774 gnd.n2773 585
R1958 gnd.n2774 gnd.n2741 585
R1959 gnd.n2772 gnd.n2739 585
R1960 gnd.n3291 gnd.n2739 585
R1961 gnd.n2728 gnd.n2726 585
R1962 gnd.n3253 gnd.n2728 585
R1963 gnd.n3299 gnd.n3298 585
R1964 gnd.n3298 gnd.n3297 585
R1965 gnd.n2727 gnd.n2725 585
R1966 gnd.n2792 gnd.n2727 585
R1967 gnd.n3224 gnd.n2791 585
R1968 gnd.n3243 gnd.n2791 585
R1969 gnd.n3226 gnd.n3225 585
R1970 gnd.n3227 gnd.n3226 585
R1971 gnd.n2801 gnd.n2800 585
R1972 gnd.n2807 gnd.n2800 585
R1973 gnd.n3219 gnd.n3218 585
R1974 gnd.n3218 gnd.n3217 585
R1975 gnd.n2804 gnd.n2803 585
R1976 gnd.n2815 gnd.n2804 585
R1977 gnd.n3104 gnd.n2823 585
R1978 gnd.n3196 gnd.n2823 585
R1979 gnd.n3106 gnd.n3105 585
R1980 gnd.n3105 gnd.n2821 585
R1981 gnd.n3107 gnd.n2834 585
R1982 gnd.n3186 gnd.n2834 585
R1983 gnd.n3109 gnd.n3108 585
R1984 gnd.n3109 gnd.n2841 585
R1985 gnd.n3111 gnd.n3110 585
R1986 gnd.n3110 gnd.n2840 585
R1987 gnd.n3112 gnd.n2851 585
R1988 gnd.n3166 gnd.n2851 585
R1989 gnd.n3114 gnd.n3113 585
R1990 gnd.n3113 gnd.n2849 585
R1991 gnd.n3115 gnd.n2860 585
R1992 gnd.n3155 gnd.n2860 585
R1993 gnd.n3117 gnd.n3116 585
R1994 gnd.n3117 gnd.n2866 585
R1995 gnd.n3119 gnd.n3118 585
R1996 gnd.n3118 gnd.n2865 585
R1997 gnd.n3120 gnd.n2881 585
R1998 gnd.n3134 gnd.n2881 585
R1999 gnd.n3121 gnd.n2934 585
R2000 gnd.n2934 gnd.n2873 585
R2001 gnd.n3123 gnd.n3122 585
R2002 gnd.n3124 gnd.n3123 585
R2003 gnd.n2935 gnd.n2933 585
R2004 gnd.n2933 gnd.n2932 585
R2005 gnd.n3088 gnd.n3087 585
R2006 gnd.n3087 gnd.n3086 585
R2007 gnd.n2938 gnd.n2937 585
R2008 gnd.n2939 gnd.n2938 585
R2009 gnd.n3077 gnd.n3076 585
R2010 gnd.n3078 gnd.n3077 585
R2011 gnd.n2947 gnd.n2946 585
R2012 gnd.n2946 gnd.n2945 585
R2013 gnd.n3072 gnd.n3071 585
R2014 gnd.n3071 gnd.n3070 585
R2015 gnd.n2950 gnd.n2949 585
R2016 gnd.n3061 gnd.n2950 585
R2017 gnd.n3060 gnd.n3059 585
R2018 gnd.n3062 gnd.n3060 585
R2019 gnd.n2958 gnd.n2957 585
R2020 gnd.n2957 gnd.n2956 585
R2021 gnd.n6968 gnd.n6967 585
R2022 gnd.n6969 gnd.n6968 585
R2023 gnd.n153 gnd.n152 585
R2024 gnd.n162 gnd.n153 585
R2025 gnd.n6977 gnd.n6976 585
R2026 gnd.n6976 gnd.n6975 585
R2027 gnd.n6978 gnd.n148 585
R2028 gnd.n148 gnd.n147 585
R2029 gnd.n6980 gnd.n6979 585
R2030 gnd.n6981 gnd.n6980 585
R2031 gnd.n133 gnd.n132 585
R2032 gnd.n144 gnd.n133 585
R2033 gnd.n6989 gnd.n6988 585
R2034 gnd.n6988 gnd.n6987 585
R2035 gnd.n6990 gnd.n128 585
R2036 gnd.n128 gnd.n127 585
R2037 gnd.n6992 gnd.n6991 585
R2038 gnd.n6993 gnd.n6992 585
R2039 gnd.n113 gnd.n112 585
R2040 gnd.n124 gnd.n113 585
R2041 gnd.n7001 gnd.n7000 585
R2042 gnd.n7000 gnd.n6999 585
R2043 gnd.n7002 gnd.n108 585
R2044 gnd.n114 gnd.n108 585
R2045 gnd.n7004 gnd.n7003 585
R2046 gnd.n7005 gnd.n7004 585
R2047 gnd.n96 gnd.n95 585
R2048 gnd.n99 gnd.n96 585
R2049 gnd.n7013 gnd.n7012 585
R2050 gnd.n7012 gnd.n7011 585
R2051 gnd.n7014 gnd.n90 585
R2052 gnd.n90 gnd.n88 585
R2053 gnd.n7016 gnd.n7015 585
R2054 gnd.n7017 gnd.n7016 585
R2055 gnd.n91 gnd.n89 585
R2056 gnd.n89 gnd.n85 585
R2057 gnd.n6932 gnd.n6931 585
R2058 gnd.n6931 gnd.n70 585
R2059 gnd.n6930 gnd.n71 585
R2060 gnd.n7025 gnd.n71 585
R2061 gnd.n6929 gnd.n6928 585
R2062 gnd.n6928 gnd.n6927 585
R2063 gnd.n498 gnd.n496 585
R2064 gnd.n499 gnd.n498 585
R2065 gnd.n6920 gnd.n6919 585
R2066 gnd.n6919 gnd.n6918 585
R2067 gnd.n504 gnd.n503 585
R2068 gnd.n6910 gnd.n504 585
R2069 gnd.n6893 gnd.n6892 585
R2070 gnd.n6892 gnd.n509 585
R2071 gnd.n6894 gnd.n519 585
R2072 gnd.n6902 gnd.n519 585
R2073 gnd.n6896 gnd.n6895 585
R2074 gnd.n6897 gnd.n6896 585
R2075 gnd.n525 gnd.n524 585
R2076 gnd.n6883 gnd.n524 585
R2077 gnd.n6859 gnd.n6858 585
R2078 gnd.n6858 gnd.n6857 585
R2079 gnd.n6860 gnd.n539 585
R2080 gnd.n6875 gnd.n539 585
R2081 gnd.n6861 gnd.n551 585
R2082 gnd.n1725 gnd.n551 585
R2083 gnd.n6863 gnd.n6862 585
R2084 gnd.n6864 gnd.n6863 585
R2085 gnd.n552 gnd.n550 585
R2086 gnd.n1732 gnd.n550 585
R2087 gnd.n5605 gnd.n1720 585
R2088 gnd.n5601 gnd.n1720 585
R2089 gnd.n5607 gnd.n5606 585
R2090 gnd.n5608 gnd.n5607 585
R2091 gnd.n1703 gnd.n1702 585
R2092 gnd.n5550 gnd.n1703 585
R2093 gnd.n5616 gnd.n5615 585
R2094 gnd.n5615 gnd.n5614 585
R2095 gnd.n5617 gnd.n1696 585
R2096 gnd.n5543 gnd.n1696 585
R2097 gnd.n5619 gnd.n5618 585
R2098 gnd.n5620 gnd.n5619 585
R2099 gnd.n1697 gnd.n1695 585
R2100 gnd.n5537 gnd.n1695 585
R2101 gnd.n1679 gnd.n1673 585
R2102 gnd.n5626 gnd.n1679 585
R2103 gnd.n5631 gnd.n1671 585
R2104 gnd.n5572 gnd.n1671 585
R2105 gnd.n5633 gnd.n5632 585
R2106 gnd.n5634 gnd.n5633 585
R2107 gnd.n1670 gnd.n1510 585
R2108 gnd.n5801 gnd.n1511 585
R2109 gnd.n5800 gnd.n1512 585
R2110 gnd.n1587 gnd.n1513 585
R2111 gnd.n5793 gnd.n1519 585
R2112 gnd.n5792 gnd.n1520 585
R2113 gnd.n1590 gnd.n1521 585
R2114 gnd.n5785 gnd.n1527 585
R2115 gnd.n5784 gnd.n1528 585
R2116 gnd.n1592 gnd.n1529 585
R2117 gnd.n5777 gnd.n1535 585
R2118 gnd.n5776 gnd.n1536 585
R2119 gnd.n1595 gnd.n1537 585
R2120 gnd.n5769 gnd.n1543 585
R2121 gnd.n5768 gnd.n1544 585
R2122 gnd.n1597 gnd.n1545 585
R2123 gnd.n5761 gnd.n1553 585
R2124 gnd.n5760 gnd.n5757 585
R2125 gnd.n1556 gnd.n1554 585
R2126 gnd.n5755 gnd.n1556 585
R2127 gnd.n199 gnd.n198 585
R2128 gnd.n250 gnd.n194 585
R2129 gnd.n252 gnd.n251 585
R2130 gnd.n254 gnd.n192 585
R2131 gnd.n256 gnd.n255 585
R2132 gnd.n257 gnd.n187 585
R2133 gnd.n259 gnd.n258 585
R2134 gnd.n261 gnd.n185 585
R2135 gnd.n263 gnd.n262 585
R2136 gnd.n264 gnd.n180 585
R2137 gnd.n266 gnd.n265 585
R2138 gnd.n268 gnd.n178 585
R2139 gnd.n270 gnd.n269 585
R2140 gnd.n271 gnd.n173 585
R2141 gnd.n273 gnd.n272 585
R2142 gnd.n275 gnd.n171 585
R2143 gnd.n277 gnd.n276 585
R2144 gnd.n278 gnd.n169 585
R2145 gnd.n279 gnd.n166 585
R2146 gnd.n166 gnd.n165 585
R2147 gnd.n246 gnd.n164 585
R2148 gnd.n6969 gnd.n164 585
R2149 gnd.n245 gnd.n244 585
R2150 gnd.n244 gnd.n162 585
R2151 gnd.n243 gnd.n155 585
R2152 gnd.n6975 gnd.n155 585
R2153 gnd.n204 gnd.n203 585
R2154 gnd.n203 gnd.n147 585
R2155 gnd.n239 gnd.n146 585
R2156 gnd.n6981 gnd.n146 585
R2157 gnd.n238 gnd.n237 585
R2158 gnd.n237 gnd.n144 585
R2159 gnd.n236 gnd.n135 585
R2160 gnd.n6987 gnd.n135 585
R2161 gnd.n207 gnd.n206 585
R2162 gnd.n206 gnd.n127 585
R2163 gnd.n232 gnd.n126 585
R2164 gnd.n6993 gnd.n126 585
R2165 gnd.n231 gnd.n230 585
R2166 gnd.n230 gnd.n124 585
R2167 gnd.n229 gnd.n116 585
R2168 gnd.n6999 gnd.n116 585
R2169 gnd.n210 gnd.n209 585
R2170 gnd.n209 gnd.n114 585
R2171 gnd.n225 gnd.n107 585
R2172 gnd.n7005 gnd.n107 585
R2173 gnd.n224 gnd.n223 585
R2174 gnd.n223 gnd.n99 585
R2175 gnd.n222 gnd.n98 585
R2176 gnd.n7011 gnd.n98 585
R2177 gnd.n213 gnd.n212 585
R2178 gnd.n212 gnd.n88 585
R2179 gnd.n218 gnd.n87 585
R2180 gnd.n7017 gnd.n87 585
R2181 gnd.n217 gnd.n216 585
R2182 gnd.n216 gnd.n85 585
R2183 gnd.n68 gnd.n67 585
R2184 gnd.n70 gnd.n68 585
R2185 gnd.n7027 gnd.n7026 585
R2186 gnd.n7026 gnd.n7025 585
R2187 gnd.n7028 gnd.n66 585
R2188 gnd.n6927 gnd.n66 585
R2189 gnd.n506 gnd.n64 585
R2190 gnd.n506 gnd.n499 585
R2191 gnd.n513 gnd.n507 585
R2192 gnd.n6918 gnd.n507 585
R2193 gnd.n6909 gnd.n6908 585
R2194 gnd.n6910 gnd.n6909 585
R2195 gnd.n512 gnd.n511 585
R2196 gnd.n511 gnd.n509 585
R2197 gnd.n6904 gnd.n6903 585
R2198 gnd.n6903 gnd.n6902 585
R2199 gnd.n516 gnd.n515 585
R2200 gnd.n6897 gnd.n516 585
R2201 gnd.n6882 gnd.n6881 585
R2202 gnd.n6883 gnd.n6882 585
R2203 gnd.n532 gnd.n531 585
R2204 gnd.n6857 gnd.n531 585
R2205 gnd.n6877 gnd.n6876 585
R2206 gnd.n6876 gnd.n6875 585
R2207 gnd.n535 gnd.n534 585
R2208 gnd.n1725 gnd.n535 585
R2209 gnd.n5554 gnd.n548 585
R2210 gnd.n6864 gnd.n548 585
R2211 gnd.n5553 gnd.n5552 585
R2212 gnd.n5552 gnd.n1732 585
R2213 gnd.n5558 gnd.n1731 585
R2214 gnd.n5601 gnd.n1731 585
R2215 gnd.n5559 gnd.n1718 585
R2216 gnd.n5608 gnd.n1718 585
R2217 gnd.n5560 gnd.n5551 585
R2218 gnd.n5551 gnd.n5550 585
R2219 gnd.n5540 gnd.n1706 585
R2220 gnd.n5614 gnd.n1706 585
R2221 gnd.n5564 gnd.n5539 585
R2222 gnd.n5543 gnd.n5539 585
R2223 gnd.n5565 gnd.n1693 585
R2224 gnd.n5620 gnd.n1693 585
R2225 gnd.n5566 gnd.n5538 585
R2226 gnd.n5538 gnd.n5537 585
R2227 gnd.n1745 gnd.n1677 585
R2228 gnd.n5626 gnd.n1677 585
R2229 gnd.n5571 gnd.n5570 585
R2230 gnd.n5572 gnd.n5571 585
R2231 gnd.n1744 gnd.n1668 585
R2232 gnd.n5634 gnd.n1668 585
R2233 gnd.n3800 gnd.n2466 585
R2234 gnd.n2466 gnd.n2443 585
R2235 gnd.n3801 gnd.n2527 585
R2236 gnd.n2527 gnd.n2517 585
R2237 gnd.n3803 gnd.n3802 585
R2238 gnd.n3804 gnd.n3803 585
R2239 gnd.n2528 gnd.n2526 585
R2240 gnd.n2535 gnd.n2526 585
R2241 gnd.n3794 gnd.n3793 585
R2242 gnd.n3793 gnd.n3792 585
R2243 gnd.n2531 gnd.n2530 585
R2244 gnd.n3519 gnd.n2531 585
R2245 gnd.n3504 gnd.n2554 585
R2246 gnd.n2554 gnd.n2544 585
R2247 gnd.n3506 gnd.n3505 585
R2248 gnd.n3507 gnd.n3506 585
R2249 gnd.n2555 gnd.n2553 585
R2250 gnd.n2553 gnd.n2551 585
R2251 gnd.n3499 gnd.n3498 585
R2252 gnd.n3498 gnd.n3497 585
R2253 gnd.n2558 gnd.n2557 585
R2254 gnd.n2567 gnd.n2558 585
R2255 gnd.n3455 gnd.n2581 585
R2256 gnd.n2581 gnd.n2566 585
R2257 gnd.n3457 gnd.n3456 585
R2258 gnd.n3458 gnd.n3457 585
R2259 gnd.n2582 gnd.n2580 585
R2260 gnd.n2589 gnd.n2580 585
R2261 gnd.n3450 gnd.n3449 585
R2262 gnd.n3449 gnd.n3448 585
R2263 gnd.n2585 gnd.n2584 585
R2264 gnd.n3429 gnd.n2585 585
R2265 gnd.n3415 gnd.n2609 585
R2266 gnd.n2609 gnd.n2598 585
R2267 gnd.n3417 gnd.n3416 585
R2268 gnd.n3418 gnd.n3417 585
R2269 gnd.n2610 gnd.n2608 585
R2270 gnd.n2608 gnd.n2605 585
R2271 gnd.n3410 gnd.n3409 585
R2272 gnd.n3409 gnd.n3408 585
R2273 gnd.n2613 gnd.n2612 585
R2274 gnd.n2623 gnd.n2613 585
R2275 gnd.n3370 gnd.n2636 585
R2276 gnd.n2636 gnd.n2622 585
R2277 gnd.n3372 gnd.n3371 585
R2278 gnd.n3373 gnd.n3372 585
R2279 gnd.n2637 gnd.n2635 585
R2280 gnd.n2644 gnd.n2635 585
R2281 gnd.n3365 gnd.n3364 585
R2282 gnd.n3364 gnd.n3363 585
R2283 gnd.n2640 gnd.n2639 585
R2284 gnd.n3344 gnd.n2640 585
R2285 gnd.n3330 gnd.n2663 585
R2286 gnd.n2663 gnd.n2653 585
R2287 gnd.n3332 gnd.n3331 585
R2288 gnd.n3333 gnd.n3332 585
R2289 gnd.n2664 gnd.n2662 585
R2290 gnd.n3321 gnd.n2662 585
R2291 gnd.n3325 gnd.n3324 585
R2292 gnd.n3324 gnd.n3323 585
R2293 gnd.n2667 gnd.n2666 585
R2294 gnd.n3276 gnd.n2667 585
R2295 gnd.n2769 gnd.n2768 585
R2296 gnd.n2770 gnd.n2769 585
R2297 gnd.n2749 gnd.n2748 585
R2298 gnd.n2752 gnd.n2749 585
R2299 gnd.n3286 gnd.n3285 585
R2300 gnd.n3285 gnd.n3284 585
R2301 gnd.n3287 gnd.n2743 585
R2302 gnd.n2779 gnd.n2743 585
R2303 gnd.n3289 gnd.n3288 585
R2304 gnd.n3290 gnd.n3289 585
R2305 gnd.n2744 gnd.n2742 585
R2306 gnd.n3254 gnd.n2742 585
R2307 gnd.n3238 gnd.n3237 585
R2308 gnd.n3237 gnd.n2730 585
R2309 gnd.n3239 gnd.n2794 585
R2310 gnd.n2794 gnd.n2729 585
R2311 gnd.n3241 gnd.n3240 585
R2312 gnd.n3242 gnd.n3241 585
R2313 gnd.n2795 gnd.n2793 585
R2314 gnd.n2793 gnd.n2790 585
R2315 gnd.n3230 gnd.n3229 585
R2316 gnd.n3229 gnd.n3228 585
R2317 gnd.n2798 gnd.n2797 585
R2318 gnd.n2805 gnd.n2798 585
R2319 gnd.n3204 gnd.n3203 585
R2320 gnd.n3205 gnd.n3204 585
R2321 gnd.n2817 gnd.n2816 585
R2322 gnd.n2824 gnd.n2816 585
R2323 gnd.n3199 gnd.n3198 585
R2324 gnd.n3198 gnd.n3197 585
R2325 gnd.n2820 gnd.n2819 585
R2326 gnd.n3187 gnd.n2820 585
R2327 gnd.n3174 gnd.n2844 585
R2328 gnd.n2844 gnd.n2843 585
R2329 gnd.n3176 gnd.n3175 585
R2330 gnd.n3177 gnd.n3176 585
R2331 gnd.n2845 gnd.n2842 585
R2332 gnd.n2852 gnd.n2842 585
R2333 gnd.n3169 gnd.n3168 585
R2334 gnd.n3168 gnd.n3167 585
R2335 gnd.n2848 gnd.n2847 585
R2336 gnd.n3156 gnd.n2848 585
R2337 gnd.n3143 gnd.n2869 585
R2338 gnd.n2869 gnd.n2868 585
R2339 gnd.n3145 gnd.n3144 585
R2340 gnd.n3146 gnd.n3145 585
R2341 gnd.n3139 gnd.n2867 585
R2342 gnd.n3138 gnd.n3137 585
R2343 gnd.n2872 gnd.n2871 585
R2344 gnd.n3135 gnd.n2872 585
R2345 gnd.n2894 gnd.n2893 585
R2346 gnd.n2897 gnd.n2896 585
R2347 gnd.n2895 gnd.n2890 585
R2348 gnd.n2902 gnd.n2901 585
R2349 gnd.n2904 gnd.n2903 585
R2350 gnd.n2907 gnd.n2906 585
R2351 gnd.n2905 gnd.n2888 585
R2352 gnd.n2912 gnd.n2911 585
R2353 gnd.n2914 gnd.n2913 585
R2354 gnd.n2917 gnd.n2916 585
R2355 gnd.n2915 gnd.n2886 585
R2356 gnd.n2922 gnd.n2921 585
R2357 gnd.n2926 gnd.n2923 585
R2358 gnd.n2927 gnd.n2864 585
R2359 gnd.n3806 gnd.n2481 585
R2360 gnd.n3873 gnd.n3872 585
R2361 gnd.n3875 gnd.n3874 585
R2362 gnd.n3877 gnd.n3876 585
R2363 gnd.n3879 gnd.n3878 585
R2364 gnd.n3881 gnd.n3880 585
R2365 gnd.n3883 gnd.n3882 585
R2366 gnd.n3885 gnd.n3884 585
R2367 gnd.n3887 gnd.n3886 585
R2368 gnd.n3889 gnd.n3888 585
R2369 gnd.n3891 gnd.n3890 585
R2370 gnd.n3893 gnd.n3892 585
R2371 gnd.n3895 gnd.n3894 585
R2372 gnd.n3898 gnd.n3897 585
R2373 gnd.n3896 gnd.n2469 585
R2374 gnd.n3902 gnd.n2467 585
R2375 gnd.n3904 gnd.n3903 585
R2376 gnd.n3905 gnd.n3904 585
R2377 gnd.n3807 gnd.n2522 585
R2378 gnd.n3807 gnd.n2443 585
R2379 gnd.n3809 gnd.n3808 585
R2380 gnd.n3808 gnd.n2517 585
R2381 gnd.n3805 gnd.n2521 585
R2382 gnd.n3805 gnd.n3804 585
R2383 gnd.n3784 gnd.n2523 585
R2384 gnd.n2535 gnd.n2523 585
R2385 gnd.n3783 gnd.n2533 585
R2386 gnd.n3792 gnd.n2533 585
R2387 gnd.n3517 gnd.n2540 585
R2388 gnd.n3519 gnd.n3517 585
R2389 gnd.n3516 gnd.n3515 585
R2390 gnd.n3516 gnd.n2544 585
R2391 gnd.n3514 gnd.n2546 585
R2392 gnd.n3507 gnd.n2546 585
R2393 gnd.n2559 gnd.n2547 585
R2394 gnd.n2559 gnd.n2551 585
R2395 gnd.n3463 gnd.n2560 585
R2396 gnd.n3497 gnd.n2560 585
R2397 gnd.n3462 gnd.n3461 585
R2398 gnd.n3461 gnd.n2567 585
R2399 gnd.n3460 gnd.n2575 585
R2400 gnd.n3460 gnd.n2566 585
R2401 gnd.n3459 gnd.n2577 585
R2402 gnd.n3459 gnd.n3458 585
R2403 gnd.n3438 gnd.n2576 585
R2404 gnd.n2589 gnd.n2576 585
R2405 gnd.n3437 gnd.n2587 585
R2406 gnd.n3448 gnd.n2587 585
R2407 gnd.n3428 gnd.n2594 585
R2408 gnd.n3429 gnd.n3428 585
R2409 gnd.n3427 gnd.n3426 585
R2410 gnd.n3427 gnd.n2598 585
R2411 gnd.n3425 gnd.n2600 585
R2412 gnd.n3418 gnd.n2600 585
R2413 gnd.n2615 gnd.n2601 585
R2414 gnd.n2615 gnd.n2605 585
R2415 gnd.n3378 gnd.n2616 585
R2416 gnd.n3408 gnd.n2616 585
R2417 gnd.n3377 gnd.n3376 585
R2418 gnd.n3376 gnd.n2623 585
R2419 gnd.n3375 gnd.n2630 585
R2420 gnd.n3375 gnd.n2622 585
R2421 gnd.n3374 gnd.n2632 585
R2422 gnd.n3374 gnd.n3373 585
R2423 gnd.n3353 gnd.n2631 585
R2424 gnd.n2644 gnd.n2631 585
R2425 gnd.n3352 gnd.n2642 585
R2426 gnd.n3363 gnd.n2642 585
R2427 gnd.n3343 gnd.n2649 585
R2428 gnd.n3344 gnd.n3343 585
R2429 gnd.n3342 gnd.n3341 585
R2430 gnd.n3342 gnd.n2653 585
R2431 gnd.n3340 gnd.n2655 585
R2432 gnd.n3333 gnd.n2655 585
R2433 gnd.n3320 gnd.n2656 585
R2434 gnd.n3321 gnd.n3320 585
R2435 gnd.n3273 gnd.n2669 585
R2436 gnd.n3323 gnd.n2669 585
R2437 gnd.n3275 gnd.n3274 585
R2438 gnd.n3276 gnd.n3275 585
R2439 gnd.n3268 gnd.n2771 585
R2440 gnd.n2771 gnd.n2770 585
R2441 gnd.n3266 gnd.n3265 585
R2442 gnd.n3265 gnd.n2752 585
R2443 gnd.n3263 gnd.n2750 585
R2444 gnd.n3284 gnd.n2750 585
R2445 gnd.n2781 gnd.n2780 585
R2446 gnd.n2780 gnd.n2779 585
R2447 gnd.n3257 gnd.n2740 585
R2448 gnd.n3290 gnd.n2740 585
R2449 gnd.n3256 gnd.n3255 585
R2450 gnd.n3255 gnd.n3254 585
R2451 gnd.n3252 gnd.n2783 585
R2452 gnd.n3252 gnd.n2730 585
R2453 gnd.n3251 gnd.n3250 585
R2454 gnd.n3251 gnd.n2729 585
R2455 gnd.n2786 gnd.n2785 585
R2456 gnd.n3242 gnd.n2785 585
R2457 gnd.n3210 gnd.n3209 585
R2458 gnd.n3209 gnd.n2790 585
R2459 gnd.n3211 gnd.n2799 585
R2460 gnd.n3228 gnd.n2799 585
R2461 gnd.n3208 gnd.n3207 585
R2462 gnd.n3207 gnd.n2805 585
R2463 gnd.n3206 gnd.n2813 585
R2464 gnd.n3206 gnd.n3205 585
R2465 gnd.n3191 gnd.n2814 585
R2466 gnd.n2824 gnd.n2814 585
R2467 gnd.n3190 gnd.n2822 585
R2468 gnd.n3197 gnd.n2822 585
R2469 gnd.n3189 gnd.n3188 585
R2470 gnd.n3188 gnd.n3187 585
R2471 gnd.n2833 gnd.n2830 585
R2472 gnd.n2843 gnd.n2833 585
R2473 gnd.n3179 gnd.n3178 585
R2474 gnd.n3178 gnd.n3177 585
R2475 gnd.n2839 gnd.n2838 585
R2476 gnd.n2852 gnd.n2839 585
R2477 gnd.n3159 gnd.n2850 585
R2478 gnd.n3167 gnd.n2850 585
R2479 gnd.n3158 gnd.n3157 585
R2480 gnd.n3157 gnd.n3156 585
R2481 gnd.n2859 gnd.n2857 585
R2482 gnd.n2868 gnd.n2859 585
R2483 gnd.n3148 gnd.n3147 585
R2484 gnd.n3147 gnd.n3146 585
R2485 gnd.n5478 gnd.n1796 585
R2486 gnd.n5478 gnd.n5477 585
R2487 gnd.n5480 gnd.n5479 585
R2488 gnd.n5479 gnd.n1784 585
R2489 gnd.n5481 gnd.n1794 585
R2490 gnd.n5404 gnd.n1794 585
R2491 gnd.n5483 gnd.n5482 585
R2492 gnd.n5484 gnd.n5483 585
R2493 gnd.n1795 gnd.n1793 585
R2494 gnd.n1793 gnd.n1790 585
R2495 gnd.n1947 gnd.n1924 585
R2496 gnd.n5396 gnd.n1924 585
R2497 gnd.n1949 gnd.n1948 585
R2498 gnd.n5367 gnd.n1949 585
R2499 gnd.n5370 gnd.n1946 585
R2500 gnd.n5370 gnd.n5369 585
R2501 gnd.n5372 gnd.n5371 585
R2502 gnd.n5371 gnd.n1931 585
R2503 gnd.n5373 gnd.n1944 585
R2504 gnd.n5360 gnd.n1944 585
R2505 gnd.n5375 gnd.n5374 585
R2506 gnd.n5376 gnd.n5375 585
R2507 gnd.n1945 gnd.n1943 585
R2508 gnd.n1943 gnd.n1939 585
R2509 gnd.n5354 gnd.n5353 585
R2510 gnd.n5355 gnd.n5354 585
R2511 gnd.n5352 gnd.n1954 585
R2512 gnd.n1960 gnd.n1954 585
R2513 gnd.n5351 gnd.n5350 585
R2514 gnd.n5350 gnd.n5349 585
R2515 gnd.n1956 gnd.n1955 585
R2516 gnd.n1957 gnd.n1956 585
R2517 gnd.n5338 gnd.n5337 585
R2518 gnd.n5339 gnd.n5338 585
R2519 gnd.n5336 gnd.n1970 585
R2520 gnd.n1970 gnd.n1967 585
R2521 gnd.n5335 gnd.n5334 585
R2522 gnd.n5334 gnd.n5333 585
R2523 gnd.n1972 gnd.n1971 585
R2524 gnd.n1979 gnd.n1972 585
R2525 gnd.n5320 gnd.n5319 585
R2526 gnd.n5321 gnd.n5320 585
R2527 gnd.n5318 gnd.n1982 585
R2528 gnd.n1982 gnd.n1978 585
R2529 gnd.n5317 gnd.n5316 585
R2530 gnd.n5316 gnd.n5315 585
R2531 gnd.n1984 gnd.n1983 585
R2532 gnd.n1995 gnd.n1984 585
R2533 gnd.n5302 gnd.n5301 585
R2534 gnd.n5303 gnd.n5302 585
R2535 gnd.n5300 gnd.n1996 585
R2536 gnd.n5294 gnd.n1996 585
R2537 gnd.n5299 gnd.n5298 585
R2538 gnd.n5298 gnd.n5297 585
R2539 gnd.n1998 gnd.n1997 585
R2540 gnd.n5284 gnd.n1998 585
R2541 gnd.n2024 gnd.n2023 585
R2542 gnd.n2024 gnd.n2003 585
R2543 gnd.n5263 gnd.n5262 585
R2544 gnd.n5262 gnd.n5261 585
R2545 gnd.n5264 gnd.n2011 585
R2546 gnd.n5275 gnd.n2011 585
R2547 gnd.n5265 gnd.n2021 585
R2548 gnd.n2021 gnd.n2010 585
R2549 gnd.n5267 gnd.n5266 585
R2550 gnd.n5268 gnd.n5267 585
R2551 gnd.n2022 gnd.n2020 585
R2552 gnd.n2032 gnd.n2020 585
R2553 gnd.n5203 gnd.n5202 585
R2554 gnd.n5203 gnd.n2033 585
R2555 gnd.n5205 gnd.n5204 585
R2556 gnd.n5204 gnd.n2031 585
R2557 gnd.n5206 gnd.n2046 585
R2558 gnd.n2046 gnd.n2044 585
R2559 gnd.n5208 gnd.n5207 585
R2560 gnd.n5209 gnd.n5208 585
R2561 gnd.n5201 gnd.n2045 585
R2562 gnd.n2045 gnd.n2040 585
R2563 gnd.n5200 gnd.n5199 585
R2564 gnd.n5199 gnd.n5198 585
R2565 gnd.n2048 gnd.n2047 585
R2566 gnd.n2049 gnd.n2048 585
R2567 gnd.n5168 gnd.n5167 585
R2568 gnd.n5168 gnd.n2058 585
R2569 gnd.n5170 gnd.n5169 585
R2570 gnd.n5169 gnd.n2057 585
R2571 gnd.n5171 gnd.n2071 585
R2572 gnd.n5156 gnd.n2071 585
R2573 gnd.n5173 gnd.n5172 585
R2574 gnd.n5174 gnd.n5173 585
R2575 gnd.n5166 gnd.n2070 585
R2576 gnd.n5162 gnd.n2070 585
R2577 gnd.n5165 gnd.n5164 585
R2578 gnd.n5164 gnd.n5163 585
R2579 gnd.n2073 gnd.n2072 585
R2580 gnd.n5136 gnd.n2073 585
R2581 gnd.n5122 gnd.n5121 585
R2582 gnd.n5121 gnd.n5120 585
R2583 gnd.n5123 gnd.n2090 585
R2584 gnd.n5119 gnd.n2090 585
R2585 gnd.n5125 gnd.n5124 585
R2586 gnd.n5126 gnd.n5125 585
R2587 gnd.n2091 gnd.n2089 585
R2588 gnd.n2089 gnd.n2084 585
R2589 gnd.n5111 gnd.n5110 585
R2590 gnd.n5112 gnd.n5111 585
R2591 gnd.n5109 gnd.n2095 585
R2592 gnd.n2102 gnd.n2095 585
R2593 gnd.n5108 gnd.n5107 585
R2594 gnd.n5107 gnd.n5106 585
R2595 gnd.n2097 gnd.n2096 585
R2596 gnd.n2099 gnd.n2097 585
R2597 gnd.n5095 gnd.n5094 585
R2598 gnd.n5096 gnd.n5095 585
R2599 gnd.n5093 gnd.n2111 585
R2600 gnd.n2111 gnd.n2108 585
R2601 gnd.n5092 gnd.n5091 585
R2602 gnd.n5091 gnd.n5090 585
R2603 gnd.n2113 gnd.n2112 585
R2604 gnd.n5017 gnd.n2113 585
R2605 gnd.n5043 gnd.n5042 585
R2606 gnd.n5043 gnd.n2122 585
R2607 gnd.n5045 gnd.n5044 585
R2608 gnd.n5044 gnd.n2121 585
R2609 gnd.n5046 gnd.n2135 585
R2610 gnd.n5031 gnd.n2135 585
R2611 gnd.n5048 gnd.n5047 585
R2612 gnd.n5049 gnd.n5048 585
R2613 gnd.n5041 gnd.n2134 585
R2614 gnd.n2134 gnd.n2130 585
R2615 gnd.n5040 gnd.n5039 585
R2616 gnd.n5039 gnd.n5038 585
R2617 gnd.n2137 gnd.n2136 585
R2618 gnd.n4908 gnd.n2137 585
R2619 gnd.n5010 gnd.n5009 585
R2620 gnd.n5011 gnd.n5010 585
R2621 gnd.n5008 gnd.n2145 585
R2622 gnd.n2145 gnd.n2142 585
R2623 gnd.n5007 gnd.n5006 585
R2624 gnd.n5006 gnd.n5005 585
R2625 gnd.n2147 gnd.n2146 585
R2626 gnd.n2158 gnd.n2147 585
R2627 gnd.n4992 gnd.n4991 585
R2628 gnd.n4993 gnd.n4992 585
R2629 gnd.n4990 gnd.n2159 585
R2630 gnd.n4984 gnd.n2159 585
R2631 gnd.n4989 gnd.n4988 585
R2632 gnd.n4988 gnd.n4987 585
R2633 gnd.n2161 gnd.n2160 585
R2634 gnd.n2162 gnd.n2161 585
R2635 gnd.n4972 gnd.n4971 585
R2636 gnd.n4973 gnd.n4972 585
R2637 gnd.n4970 gnd.n2169 585
R2638 gnd.n4966 gnd.n2169 585
R2639 gnd.n4969 gnd.n4968 585
R2640 gnd.n4968 gnd.n4967 585
R2641 gnd.n2171 gnd.n2170 585
R2642 gnd.n4930 gnd.n2171 585
R2643 gnd.n4958 gnd.n4957 585
R2644 gnd.n4959 gnd.n4958 585
R2645 gnd.n4956 gnd.n2177 585
R2646 gnd.n2177 gnd.n2176 585
R2647 gnd.n4955 gnd.n4954 585
R2648 gnd.n4954 gnd.n4953 585
R2649 gnd.n2179 gnd.n2178 585
R2650 gnd.n2184 gnd.n2179 585
R2651 gnd.n4946 gnd.n4945 585
R2652 gnd.n4947 gnd.n4946 585
R2653 gnd.n4944 gnd.n2186 585
R2654 gnd.n2191 gnd.n2186 585
R2655 gnd.n4943 gnd.n4942 585
R2656 gnd.n4942 gnd.n4941 585
R2657 gnd.n2188 gnd.n2187 585
R2658 gnd.n4852 gnd.n2188 585
R2659 gnd.n4871 gnd.n4870 585
R2660 gnd.n4871 gnd.n2223 585
R2661 gnd.n4873 gnd.n4872 585
R2662 gnd.n4872 gnd.n2222 585
R2663 gnd.n4874 gnd.n2234 585
R2664 gnd.n2234 gnd.n2232 585
R2665 gnd.n4876 gnd.n4875 585
R2666 gnd.n4877 gnd.n4876 585
R2667 gnd.n4869 gnd.n2233 585
R2668 gnd.n4864 gnd.n2233 585
R2669 gnd.n4868 gnd.n4867 585
R2670 gnd.n4867 gnd.n4866 585
R2671 gnd.n2236 gnd.n2235 585
R2672 gnd.n4846 gnd.n2236 585
R2673 gnd.n4799 gnd.n4798 585
R2674 gnd.n4798 gnd.n2241 585
R2675 gnd.n4801 gnd.n4800 585
R2676 gnd.n4801 gnd.n2243 585
R2677 gnd.n4816 gnd.n4797 585
R2678 gnd.n4816 gnd.n4815 585
R2679 gnd.n4818 gnd.n4817 585
R2680 gnd.n4817 gnd.n1394 585
R2681 gnd.n4819 gnd.n4796 585
R2682 gnd.n4796 gnd.n1392 585
R2683 gnd.n4821 gnd.n4820 585
R2684 gnd.n4822 gnd.n4821 585
R2685 gnd.n1376 gnd.n1375 585
R2686 gnd.n1380 gnd.n1376 585
R2687 gnd.n5942 gnd.n5941 585
R2688 gnd.n5941 gnd.n5940 585
R2689 gnd.n5943 gnd.n1373 585
R2690 gnd.n1377 gnd.n1373 585
R2691 gnd.n5945 gnd.n5944 585
R2692 gnd.n5946 gnd.n5945 585
R2693 gnd.n1374 gnd.n1372 585
R2694 gnd.n1372 gnd.n1292 585
R2695 gnd.n4773 gnd.n1290 585
R2696 gnd.n5952 gnd.n1290 585
R2697 gnd.n4775 gnd.n4774 585
R2698 gnd.n4776 gnd.n4775 585
R2699 gnd.n4772 gnd.n4771 585
R2700 gnd.n4771 gnd.n1280 585
R2701 gnd.n1275 gnd.n1274 585
R2702 gnd.n5959 gnd.n1275 585
R2703 gnd.n5962 gnd.n5961 585
R2704 gnd.n5961 gnd.n5960 585
R2705 gnd.n5963 gnd.n1253 585
R2706 gnd.n1361 gnd.n1253 585
R2707 gnd.n6028 gnd.n6027 585
R2708 gnd.n6026 gnd.n1252 585
R2709 gnd.n6025 gnd.n1251 585
R2710 gnd.n6030 gnd.n1251 585
R2711 gnd.n6024 gnd.n6023 585
R2712 gnd.n6022 gnd.n6021 585
R2713 gnd.n6020 gnd.n6019 585
R2714 gnd.n6018 gnd.n6017 585
R2715 gnd.n6016 gnd.n6015 585
R2716 gnd.n6014 gnd.n6013 585
R2717 gnd.n6012 gnd.n6011 585
R2718 gnd.n6010 gnd.n6009 585
R2719 gnd.n6008 gnd.n6007 585
R2720 gnd.n6006 gnd.n6005 585
R2721 gnd.n6004 gnd.n6003 585
R2722 gnd.n6002 gnd.n6001 585
R2723 gnd.n6000 gnd.n5999 585
R2724 gnd.n5998 gnd.n5997 585
R2725 gnd.n5996 gnd.n5995 585
R2726 gnd.n5994 gnd.n5993 585
R2727 gnd.n5992 gnd.n5991 585
R2728 gnd.n5990 gnd.n5989 585
R2729 gnd.n5988 gnd.n5987 585
R2730 gnd.n5986 gnd.n5985 585
R2731 gnd.n5984 gnd.n5983 585
R2732 gnd.n5982 gnd.n5981 585
R2733 gnd.n5980 gnd.n5979 585
R2734 gnd.n5978 gnd.n5977 585
R2735 gnd.n5976 gnd.n5975 585
R2736 gnd.n5974 gnd.n5973 585
R2737 gnd.n5972 gnd.n5971 585
R2738 gnd.n5970 gnd.n5969 585
R2739 gnd.n5968 gnd.n1215 585
R2740 gnd.n6033 gnd.n6032 585
R2741 gnd.n1217 gnd.n1214 585
R2742 gnd.n1299 gnd.n1298 585
R2743 gnd.n1301 gnd.n1300 585
R2744 gnd.n1304 gnd.n1303 585
R2745 gnd.n1306 gnd.n1305 585
R2746 gnd.n1308 gnd.n1307 585
R2747 gnd.n1310 gnd.n1309 585
R2748 gnd.n1312 gnd.n1311 585
R2749 gnd.n1314 gnd.n1313 585
R2750 gnd.n1316 gnd.n1315 585
R2751 gnd.n1318 gnd.n1317 585
R2752 gnd.n1320 gnd.n1319 585
R2753 gnd.n1322 gnd.n1321 585
R2754 gnd.n1324 gnd.n1323 585
R2755 gnd.n1326 gnd.n1325 585
R2756 gnd.n1328 gnd.n1327 585
R2757 gnd.n1330 gnd.n1329 585
R2758 gnd.n1332 gnd.n1331 585
R2759 gnd.n1334 gnd.n1333 585
R2760 gnd.n1336 gnd.n1335 585
R2761 gnd.n1338 gnd.n1337 585
R2762 gnd.n1340 gnd.n1339 585
R2763 gnd.n1342 gnd.n1341 585
R2764 gnd.n1344 gnd.n1343 585
R2765 gnd.n1346 gnd.n1345 585
R2766 gnd.n1348 gnd.n1347 585
R2767 gnd.n1350 gnd.n1349 585
R2768 gnd.n1352 gnd.n1351 585
R2769 gnd.n1354 gnd.n1353 585
R2770 gnd.n1356 gnd.n1355 585
R2771 gnd.n1358 gnd.n1357 585
R2772 gnd.n1360 gnd.n1359 585
R2773 gnd.n5410 gnd.n5409 585
R2774 gnd.n5412 gnd.n5411 585
R2775 gnd.n5414 gnd.n5413 585
R2776 gnd.n5416 gnd.n5415 585
R2777 gnd.n5418 gnd.n5417 585
R2778 gnd.n5420 gnd.n5419 585
R2779 gnd.n5422 gnd.n5421 585
R2780 gnd.n5424 gnd.n5423 585
R2781 gnd.n5426 gnd.n5425 585
R2782 gnd.n5428 gnd.n5427 585
R2783 gnd.n5430 gnd.n5429 585
R2784 gnd.n5432 gnd.n5431 585
R2785 gnd.n5434 gnd.n5433 585
R2786 gnd.n5436 gnd.n5435 585
R2787 gnd.n5438 gnd.n5437 585
R2788 gnd.n5440 gnd.n5439 585
R2789 gnd.n5442 gnd.n5441 585
R2790 gnd.n5444 gnd.n5443 585
R2791 gnd.n5446 gnd.n5445 585
R2792 gnd.n5448 gnd.n5447 585
R2793 gnd.n5450 gnd.n5449 585
R2794 gnd.n5452 gnd.n5451 585
R2795 gnd.n5454 gnd.n5453 585
R2796 gnd.n5456 gnd.n5455 585
R2797 gnd.n5458 gnd.n5457 585
R2798 gnd.n5460 gnd.n5459 585
R2799 gnd.n5462 gnd.n5461 585
R2800 gnd.n5464 gnd.n5463 585
R2801 gnd.n5466 gnd.n5465 585
R2802 gnd.n5469 gnd.n5468 585
R2803 gnd.n5471 gnd.n5470 585
R2804 gnd.n5473 gnd.n5472 585
R2805 gnd.n5475 gnd.n5474 585
R2806 gnd.n1901 gnd.n1631 585
R2807 gnd.n1900 gnd.n1899 585
R2808 gnd.n1898 gnd.n1897 585
R2809 gnd.n1896 gnd.n1895 585
R2810 gnd.n1893 gnd.n1892 585
R2811 gnd.n1891 gnd.n1890 585
R2812 gnd.n1889 gnd.n1888 585
R2813 gnd.n1887 gnd.n1886 585
R2814 gnd.n1885 gnd.n1884 585
R2815 gnd.n1883 gnd.n1882 585
R2816 gnd.n1881 gnd.n1880 585
R2817 gnd.n1879 gnd.n1878 585
R2818 gnd.n1877 gnd.n1876 585
R2819 gnd.n1875 gnd.n1874 585
R2820 gnd.n1873 gnd.n1872 585
R2821 gnd.n1871 gnd.n1870 585
R2822 gnd.n1869 gnd.n1868 585
R2823 gnd.n1867 gnd.n1866 585
R2824 gnd.n1865 gnd.n1864 585
R2825 gnd.n1863 gnd.n1862 585
R2826 gnd.n1861 gnd.n1860 585
R2827 gnd.n1859 gnd.n1858 585
R2828 gnd.n1857 gnd.n1856 585
R2829 gnd.n1855 gnd.n1854 585
R2830 gnd.n1853 gnd.n1852 585
R2831 gnd.n1851 gnd.n1850 585
R2832 gnd.n1849 gnd.n1848 585
R2833 gnd.n1847 gnd.n1846 585
R2834 gnd.n1845 gnd.n1844 585
R2835 gnd.n1843 gnd.n1842 585
R2836 gnd.n1841 gnd.n1840 585
R2837 gnd.n1839 gnd.n1838 585
R2838 gnd.n1837 gnd.n1797 585
R2839 gnd.n5408 gnd.n1798 585
R2840 gnd.n5477 gnd.n1798 585
R2841 gnd.n5407 gnd.n5406 585
R2842 gnd.n5406 gnd.n1784 585
R2843 gnd.n5405 gnd.n5401 585
R2844 gnd.n5405 gnd.n5404 585
R2845 gnd.n5400 gnd.n1792 585
R2846 gnd.n5484 gnd.n1792 585
R2847 gnd.n5399 gnd.n5398 585
R2848 gnd.n5398 gnd.n1790 585
R2849 gnd.n5397 gnd.n1922 585
R2850 gnd.n5397 gnd.n5396 585
R2851 gnd.n5364 gnd.n1923 585
R2852 gnd.n5367 gnd.n1923 585
R2853 gnd.n5366 gnd.n5365 585
R2854 gnd.n5369 gnd.n5366 585
R2855 gnd.n5363 gnd.n1950 585
R2856 gnd.n1950 gnd.n1931 585
R2857 gnd.n5362 gnd.n5361 585
R2858 gnd.n5361 gnd.n5360 585
R2859 gnd.n5359 gnd.n1941 585
R2860 gnd.n5376 gnd.n1941 585
R2861 gnd.n5358 gnd.n5357 585
R2862 gnd.n5357 gnd.n1939 585
R2863 gnd.n5356 gnd.n1951 585
R2864 gnd.n5356 gnd.n5355 585
R2865 gnd.n5325 gnd.n1952 585
R2866 gnd.n1960 gnd.n1952 585
R2867 gnd.n5326 gnd.n1958 585
R2868 gnd.n5349 gnd.n1958 585
R2869 gnd.n5328 gnd.n5327 585
R2870 gnd.n5327 gnd.n1957 585
R2871 gnd.n5329 gnd.n1969 585
R2872 gnd.n5339 gnd.n1969 585
R2873 gnd.n5330 gnd.n1975 585
R2874 gnd.n1975 gnd.n1967 585
R2875 gnd.n5332 gnd.n5331 585
R2876 gnd.n5333 gnd.n5332 585
R2877 gnd.n5324 gnd.n1974 585
R2878 gnd.n1979 gnd.n1974 585
R2879 gnd.n5323 gnd.n5322 585
R2880 gnd.n5322 gnd.n5321 585
R2881 gnd.n1977 gnd.n1976 585
R2882 gnd.n1978 gnd.n1977 585
R2883 gnd.n5288 gnd.n1985 585
R2884 gnd.n5315 gnd.n1985 585
R2885 gnd.n5290 gnd.n5289 585
R2886 gnd.n5289 gnd.n1995 585
R2887 gnd.n5291 gnd.n1994 585
R2888 gnd.n5303 gnd.n1994 585
R2889 gnd.n5293 gnd.n5292 585
R2890 gnd.n5294 gnd.n5293 585
R2891 gnd.n5287 gnd.n1999 585
R2892 gnd.n5297 gnd.n1999 585
R2893 gnd.n5286 gnd.n5285 585
R2894 gnd.n5285 gnd.n5284 585
R2895 gnd.n2002 gnd.n2001 585
R2896 gnd.n2003 gnd.n2002 585
R2897 gnd.n5272 gnd.n2014 585
R2898 gnd.n5261 gnd.n2014 585
R2899 gnd.n5274 gnd.n5273 585
R2900 gnd.n5275 gnd.n5274 585
R2901 gnd.n5271 gnd.n2013 585
R2902 gnd.n2013 gnd.n2010 585
R2903 gnd.n5270 gnd.n5269 585
R2904 gnd.n5269 gnd.n5268 585
R2905 gnd.n2016 gnd.n2015 585
R2906 gnd.n2032 gnd.n2016 585
R2907 gnd.n5144 gnd.n5143 585
R2908 gnd.n5144 gnd.n2033 585
R2909 gnd.n5145 gnd.n5142 585
R2910 gnd.n5145 gnd.n2031 585
R2911 gnd.n5147 gnd.n5146 585
R2912 gnd.n5146 gnd.n2044 585
R2913 gnd.n5148 gnd.n2042 585
R2914 gnd.n5209 gnd.n2042 585
R2915 gnd.n5150 gnd.n5149 585
R2916 gnd.n5149 gnd.n2040 585
R2917 gnd.n5151 gnd.n2050 585
R2918 gnd.n5198 gnd.n2050 585
R2919 gnd.n5152 gnd.n5141 585
R2920 gnd.n5141 gnd.n2049 585
R2921 gnd.n5154 gnd.n5153 585
R2922 gnd.n5154 gnd.n2058 585
R2923 gnd.n5155 gnd.n5140 585
R2924 gnd.n5155 gnd.n2057 585
R2925 gnd.n5158 gnd.n5157 585
R2926 gnd.n5157 gnd.n5156 585
R2927 gnd.n5159 gnd.n2067 585
R2928 gnd.n5174 gnd.n2067 585
R2929 gnd.n5161 gnd.n5160 585
R2930 gnd.n5162 gnd.n5161 585
R2931 gnd.n5139 gnd.n2075 585
R2932 gnd.n5163 gnd.n2075 585
R2933 gnd.n5138 gnd.n5137 585
R2934 gnd.n5137 gnd.n5136 585
R2935 gnd.n2077 gnd.n2076 585
R2936 gnd.n5120 gnd.n2077 585
R2937 gnd.n5118 gnd.n5117 585
R2938 gnd.n5119 gnd.n5118 585
R2939 gnd.n5116 gnd.n2086 585
R2940 gnd.n5126 gnd.n2086 585
R2941 gnd.n5115 gnd.n5114 585
R2942 gnd.n5114 gnd.n2084 585
R2943 gnd.n5113 gnd.n2092 585
R2944 gnd.n5113 gnd.n5112 585
R2945 gnd.n5019 gnd.n2093 585
R2946 gnd.n2102 gnd.n2093 585
R2947 gnd.n5020 gnd.n2100 585
R2948 gnd.n5106 gnd.n2100 585
R2949 gnd.n5022 gnd.n5021 585
R2950 gnd.n5021 gnd.n2099 585
R2951 gnd.n5023 gnd.n2110 585
R2952 gnd.n5096 gnd.n2110 585
R2953 gnd.n5025 gnd.n5024 585
R2954 gnd.n5024 gnd.n2108 585
R2955 gnd.n5026 gnd.n2114 585
R2956 gnd.n5090 gnd.n2114 585
R2957 gnd.n5027 gnd.n5018 585
R2958 gnd.n5018 gnd.n5017 585
R2959 gnd.n5029 gnd.n5028 585
R2960 gnd.n5029 gnd.n2122 585
R2961 gnd.n5030 gnd.n5015 585
R2962 gnd.n5030 gnd.n2121 585
R2963 gnd.n5033 gnd.n5032 585
R2964 gnd.n5032 gnd.n5031 585
R2965 gnd.n5034 gnd.n2132 585
R2966 gnd.n5049 gnd.n2132 585
R2967 gnd.n5035 gnd.n2139 585
R2968 gnd.n2139 gnd.n2130 585
R2969 gnd.n5037 gnd.n5036 585
R2970 gnd.n5038 gnd.n5037 585
R2971 gnd.n5014 gnd.n2138 585
R2972 gnd.n4908 gnd.n2138 585
R2973 gnd.n5013 gnd.n5012 585
R2974 gnd.n5012 gnd.n5011 585
R2975 gnd.n2141 gnd.n2140 585
R2976 gnd.n2142 gnd.n2141 585
R2977 gnd.n4978 gnd.n2148 585
R2978 gnd.n5005 gnd.n2148 585
R2979 gnd.n4980 gnd.n4979 585
R2980 gnd.n4979 gnd.n2158 585
R2981 gnd.n4981 gnd.n2157 585
R2982 gnd.n4993 gnd.n2157 585
R2983 gnd.n4983 gnd.n4982 585
R2984 gnd.n4984 gnd.n4983 585
R2985 gnd.n4977 gnd.n2163 585
R2986 gnd.n4987 gnd.n2163 585
R2987 gnd.n4976 gnd.n4975 585
R2988 gnd.n4975 gnd.n2162 585
R2989 gnd.n4974 gnd.n2165 585
R2990 gnd.n4974 gnd.n4973 585
R2991 gnd.n4963 gnd.n2166 585
R2992 gnd.n4966 gnd.n2166 585
R2993 gnd.n4965 gnd.n4964 585
R2994 gnd.n4967 gnd.n4965 585
R2995 gnd.n4962 gnd.n2173 585
R2996 gnd.n4930 gnd.n2173 585
R2997 gnd.n4961 gnd.n4960 585
R2998 gnd.n4960 gnd.n4959 585
R2999 gnd.n2175 gnd.n2174 585
R3000 gnd.n2176 gnd.n2175 585
R3001 gnd.n4952 gnd.n4951 585
R3002 gnd.n4953 gnd.n4952 585
R3003 gnd.n4950 gnd.n2181 585
R3004 gnd.n2184 gnd.n2181 585
R3005 gnd.n4949 gnd.n4948 585
R3006 gnd.n4948 gnd.n4947 585
R3007 gnd.n2183 gnd.n2182 585
R3008 gnd.n2191 gnd.n2183 585
R3009 gnd.n4854 gnd.n2189 585
R3010 gnd.n4941 gnd.n2189 585
R3011 gnd.n4855 gnd.n4853 585
R3012 gnd.n4853 gnd.n4852 585
R3013 gnd.n4857 gnd.n4856 585
R3014 gnd.n4857 gnd.n2223 585
R3015 gnd.n4858 gnd.n4850 585
R3016 gnd.n4858 gnd.n2222 585
R3017 gnd.n4860 gnd.n4859 585
R3018 gnd.n4859 gnd.n2232 585
R3019 gnd.n4861 gnd.n2230 585
R3020 gnd.n4877 gnd.n2230 585
R3021 gnd.n4863 gnd.n4862 585
R3022 gnd.n4864 gnd.n4863 585
R3023 gnd.n4849 gnd.n2237 585
R3024 gnd.n4866 gnd.n2237 585
R3025 gnd.n4848 gnd.n4847 585
R3026 gnd.n4847 gnd.n4846 585
R3027 gnd.n2240 gnd.n2239 585
R3028 gnd.n2241 gnd.n2240 585
R3029 gnd.n4812 gnd.n4804 585
R3030 gnd.n4804 gnd.n2243 585
R3031 gnd.n4814 gnd.n4813 585
R3032 gnd.n4815 gnd.n4814 585
R3033 gnd.n4811 gnd.n4803 585
R3034 gnd.n4803 gnd.n1394 585
R3035 gnd.n4810 gnd.n4809 585
R3036 gnd.n4809 gnd.n1392 585
R3037 gnd.n4808 gnd.n4795 585
R3038 gnd.n4822 gnd.n4795 585
R3039 gnd.n4807 gnd.n4806 585
R3040 gnd.n4806 gnd.n1380 585
R3041 gnd.n4805 gnd.n1378 585
R3042 gnd.n5940 gnd.n1378 585
R3043 gnd.n1370 gnd.n1369 585
R3044 gnd.n1377 gnd.n1370 585
R3045 gnd.n5948 gnd.n5947 585
R3046 gnd.n5947 gnd.n5946 585
R3047 gnd.n5949 gnd.n1295 585
R3048 gnd.n1295 gnd.n1292 585
R3049 gnd.n5951 gnd.n5950 585
R3050 gnd.n5952 gnd.n5951 585
R3051 gnd.n1368 gnd.n1294 585
R3052 gnd.n4776 gnd.n1294 585
R3053 gnd.n1367 gnd.n1366 585
R3054 gnd.n1366 gnd.n1280 585
R3055 gnd.n1365 gnd.n1278 585
R3056 gnd.n5959 gnd.n1278 585
R3057 gnd.n1364 gnd.n1277 585
R3058 gnd.n5960 gnd.n1277 585
R3059 gnd.n1363 gnd.n1362 585
R3060 gnd.n1362 gnd.n1361 585
R3061 gnd.n6089 gnd.n1138 585
R3062 gnd.n4714 gnd.n1138 585
R3063 gnd.n6091 gnd.n6090 585
R3064 gnd.n6092 gnd.n6091 585
R3065 gnd.n1123 gnd.n1122 585
R3066 gnd.n4677 gnd.n1123 585
R3067 gnd.n6100 gnd.n6099 585
R3068 gnd.n6099 gnd.n6098 585
R3069 gnd.n6101 gnd.n1117 585
R3070 gnd.n4437 gnd.n1117 585
R3071 gnd.n6103 gnd.n6102 585
R3072 gnd.n6104 gnd.n6103 585
R3073 gnd.n1103 gnd.n1102 585
R3074 gnd.n4690 gnd.n1103 585
R3075 gnd.n6112 gnd.n6111 585
R3076 gnd.n6111 gnd.n6110 585
R3077 gnd.n6113 gnd.n1097 585
R3078 gnd.n4430 gnd.n1097 585
R3079 gnd.n6115 gnd.n6114 585
R3080 gnd.n6116 gnd.n6115 585
R3081 gnd.n1083 gnd.n1082 585
R3082 gnd.n4422 gnd.n1083 585
R3083 gnd.n6124 gnd.n6123 585
R3084 gnd.n6123 gnd.n6122 585
R3085 gnd.n6125 gnd.n1077 585
R3086 gnd.n4387 gnd.n1077 585
R3087 gnd.n6127 gnd.n6126 585
R3088 gnd.n6128 gnd.n6127 585
R3089 gnd.n1061 gnd.n1060 585
R3090 gnd.n4395 gnd.n1061 585
R3091 gnd.n6136 gnd.n6135 585
R3092 gnd.n6135 gnd.n6134 585
R3093 gnd.n6137 gnd.n1056 585
R3094 gnd.n4376 gnd.n1056 585
R3095 gnd.n6139 gnd.n6138 585
R3096 gnd.n6140 gnd.n6139 585
R3097 gnd.n4364 gnd.n1055 585
R3098 gnd.n1055 gnd.n1050 585
R3099 gnd.n4366 gnd.n4365 585
R3100 gnd.n4367 gnd.n4366 585
R3101 gnd.n4362 gnd.n2336 585
R3102 gnd.n2342 gnd.n2336 585
R3103 gnd.n4361 gnd.n4360 585
R3104 gnd.n4360 gnd.n4359 585
R3105 gnd.n4337 gnd.n2338 585
R3106 gnd.n2339 gnd.n2338 585
R3107 gnd.n4339 gnd.n4338 585
R3108 gnd.n4340 gnd.n4339 585
R3109 gnd.n4335 gnd.n2355 585
R3110 gnd.n2355 gnd.n2352 585
R3111 gnd.n4334 gnd.n4333 585
R3112 gnd.n4333 gnd.n4332 585
R3113 gnd.n4317 gnd.n2357 585
R3114 gnd.n2358 gnd.n2357 585
R3115 gnd.n4319 gnd.n4318 585
R3116 gnd.n4320 gnd.n4319 585
R3117 gnd.n2371 gnd.n2370 585
R3118 gnd.n2378 gnd.n2370 585
R3119 gnd.n4313 gnd.n4312 585
R3120 gnd.n4312 gnd.n4311 585
R3121 gnd.n2374 gnd.n2373 585
R3122 gnd.n2375 gnd.n2374 585
R3123 gnd.n4298 gnd.n4297 585
R3124 gnd.n4299 gnd.n4298 585
R3125 gnd.n2390 gnd.n2389 585
R3126 gnd.n2389 gnd.n2386 585
R3127 gnd.n4293 gnd.n4292 585
R3128 gnd.n4292 gnd.n4291 585
R3129 gnd.n2393 gnd.n2392 585
R3130 gnd.n2394 gnd.n2393 585
R3131 gnd.n4278 gnd.n4277 585
R3132 gnd.n4279 gnd.n4278 585
R3133 gnd.n2407 gnd.n2406 585
R3134 gnd.n2414 gnd.n2406 585
R3135 gnd.n4273 gnd.n4272 585
R3136 gnd.n4272 gnd.n4271 585
R3137 gnd.n2410 gnd.n2409 585
R3138 gnd.n2411 gnd.n2410 585
R3139 gnd.n4258 gnd.n4257 585
R3140 gnd.n4259 gnd.n4258 585
R3141 gnd.n2426 gnd.n2425 585
R3142 gnd.n2425 gnd.n2422 585
R3143 gnd.n4253 gnd.n4252 585
R3144 gnd.n4252 gnd.n4251 585
R3145 gnd.n2429 gnd.n2428 585
R3146 gnd.n2430 gnd.n2429 585
R3147 gnd.n4239 gnd.n4238 585
R3148 gnd.n4237 gnd.n3944 585
R3149 gnd.n4236 gnd.n3943 585
R3150 gnd.n4241 gnd.n3943 585
R3151 gnd.n4235 gnd.n4234 585
R3152 gnd.n4233 gnd.n4232 585
R3153 gnd.n4231 gnd.n4230 585
R3154 gnd.n4229 gnd.n4228 585
R3155 gnd.n4227 gnd.n4226 585
R3156 gnd.n4225 gnd.n4224 585
R3157 gnd.n4223 gnd.n4222 585
R3158 gnd.n4221 gnd.n4220 585
R3159 gnd.n4219 gnd.n4218 585
R3160 gnd.n4217 gnd.n4216 585
R3161 gnd.n4215 gnd.n4214 585
R3162 gnd.n4213 gnd.n4212 585
R3163 gnd.n4211 gnd.n4210 585
R3164 gnd.n4209 gnd.n4208 585
R3165 gnd.n4207 gnd.n4206 585
R3166 gnd.n4204 gnd.n4203 585
R3167 gnd.n4202 gnd.n4201 585
R3168 gnd.n4200 gnd.n4199 585
R3169 gnd.n4198 gnd.n4197 585
R3170 gnd.n4196 gnd.n4195 585
R3171 gnd.n4194 gnd.n4193 585
R3172 gnd.n4192 gnd.n4191 585
R3173 gnd.n4190 gnd.n4189 585
R3174 gnd.n4188 gnd.n4187 585
R3175 gnd.n4186 gnd.n4185 585
R3176 gnd.n4184 gnd.n4183 585
R3177 gnd.n4182 gnd.n4181 585
R3178 gnd.n4180 gnd.n4179 585
R3179 gnd.n4178 gnd.n4177 585
R3180 gnd.n4176 gnd.n4175 585
R3181 gnd.n4174 gnd.n4173 585
R3182 gnd.n4172 gnd.n4171 585
R3183 gnd.n4170 gnd.n4169 585
R3184 gnd.n4168 gnd.n4167 585
R3185 gnd.n4166 gnd.n4165 585
R3186 gnd.n4164 gnd.n4163 585
R3187 gnd.n4162 gnd.n4161 585
R3188 gnd.n4160 gnd.n4159 585
R3189 gnd.n4158 gnd.n4157 585
R3190 gnd.n4156 gnd.n4155 585
R3191 gnd.n4154 gnd.n4153 585
R3192 gnd.n4152 gnd.n4151 585
R3193 gnd.n4150 gnd.n4149 585
R3194 gnd.n4148 gnd.n4147 585
R3195 gnd.n4146 gnd.n4145 585
R3196 gnd.n4144 gnd.n4143 585
R3197 gnd.n4142 gnd.n4141 585
R3198 gnd.n4140 gnd.n4139 585
R3199 gnd.n4138 gnd.n4137 585
R3200 gnd.n4136 gnd.n4135 585
R3201 gnd.n4134 gnd.n4133 585
R3202 gnd.n4132 gnd.n4131 585
R3203 gnd.n4130 gnd.n4129 585
R3204 gnd.n4128 gnd.n4127 585
R3205 gnd.n4126 gnd.n2442 585
R3206 gnd.n4243 gnd.n2441 585
R3207 gnd.n4669 gnd.n4668 585
R3208 gnd.n4667 gnd.n4578 585
R3209 gnd.n4666 gnd.n4665 585
R3210 gnd.n4659 gnd.n4579 585
R3211 gnd.n4661 gnd.n4660 585
R3212 gnd.n4658 gnd.n4657 585
R3213 gnd.n4656 gnd.n4655 585
R3214 gnd.n4649 gnd.n4581 585
R3215 gnd.n4651 gnd.n4650 585
R3216 gnd.n4648 gnd.n4647 585
R3217 gnd.n4646 gnd.n4645 585
R3218 gnd.n4639 gnd.n4583 585
R3219 gnd.n4641 gnd.n4640 585
R3220 gnd.n4638 gnd.n4637 585
R3221 gnd.n4636 gnd.n4635 585
R3222 gnd.n4629 gnd.n4585 585
R3223 gnd.n4631 gnd.n4630 585
R3224 gnd.n4628 gnd.n4627 585
R3225 gnd.n4626 gnd.n4625 585
R3226 gnd.n4619 gnd.n4587 585
R3227 gnd.n4621 gnd.n4620 585
R3228 gnd.n4618 gnd.n4591 585
R3229 gnd.n4617 gnd.n4616 585
R3230 gnd.n4610 gnd.n4592 585
R3231 gnd.n4612 gnd.n4611 585
R3232 gnd.n4609 gnd.n4608 585
R3233 gnd.n4607 gnd.n4606 585
R3234 gnd.n4600 gnd.n4594 585
R3235 gnd.n4602 gnd.n4601 585
R3236 gnd.n4599 gnd.n4598 585
R3237 gnd.n4597 gnd.n1211 585
R3238 gnd.n6036 gnd.n6035 585
R3239 gnd.n6038 gnd.n6037 585
R3240 gnd.n6040 gnd.n6039 585
R3241 gnd.n6042 gnd.n6041 585
R3242 gnd.n6044 gnd.n6043 585
R3243 gnd.n6046 gnd.n6045 585
R3244 gnd.n6048 gnd.n6047 585
R3245 gnd.n6050 gnd.n6049 585
R3246 gnd.n6053 gnd.n6052 585
R3247 gnd.n6055 gnd.n6054 585
R3248 gnd.n6057 gnd.n6056 585
R3249 gnd.n6059 gnd.n6058 585
R3250 gnd.n6061 gnd.n6060 585
R3251 gnd.n6063 gnd.n6062 585
R3252 gnd.n6065 gnd.n6064 585
R3253 gnd.n6067 gnd.n6066 585
R3254 gnd.n6069 gnd.n6068 585
R3255 gnd.n6071 gnd.n6070 585
R3256 gnd.n6073 gnd.n6072 585
R3257 gnd.n6075 gnd.n6074 585
R3258 gnd.n6077 gnd.n6076 585
R3259 gnd.n6079 gnd.n6078 585
R3260 gnd.n6080 gnd.n1184 585
R3261 gnd.n6082 gnd.n6081 585
R3262 gnd.n1143 gnd.n1142 585
R3263 gnd.n6086 gnd.n6085 585
R3264 gnd.n6085 gnd.n6084 585
R3265 gnd.n4673 gnd.n2296 585
R3266 gnd.n4714 gnd.n2296 585
R3267 gnd.n4674 gnd.n1135 585
R3268 gnd.n6092 gnd.n1135 585
R3269 gnd.n4676 gnd.n4675 585
R3270 gnd.n4677 gnd.n4676 585
R3271 gnd.n4440 gnd.n1125 585
R3272 gnd.n6098 gnd.n1125 585
R3273 gnd.n4439 gnd.n4438 585
R3274 gnd.n4438 gnd.n4437 585
R3275 gnd.n4435 gnd.n1114 585
R3276 gnd.n6104 gnd.n1114 585
R3277 gnd.n4434 gnd.n2307 585
R3278 gnd.n4690 gnd.n2307 585
R3279 gnd.n4433 gnd.n1105 585
R3280 gnd.n6110 gnd.n1105 585
R3281 gnd.n4432 gnd.n4431 585
R3282 gnd.n4431 gnd.n4430 585
R3283 gnd.n2313 gnd.n1094 585
R3284 gnd.n6116 gnd.n1094 585
R3285 gnd.n4383 gnd.n2318 585
R3286 gnd.n4422 gnd.n2318 585
R3287 gnd.n4384 gnd.n1085 585
R3288 gnd.n6122 gnd.n1085 585
R3289 gnd.n4386 gnd.n4385 585
R3290 gnd.n4387 gnd.n4386 585
R3291 gnd.n4381 gnd.n1074 585
R3292 gnd.n6128 gnd.n1074 585
R3293 gnd.n4380 gnd.n2324 585
R3294 gnd.n4395 gnd.n2324 585
R3295 gnd.n4379 gnd.n1063 585
R3296 gnd.n6134 gnd.n1063 585
R3297 gnd.n4378 gnd.n4377 585
R3298 gnd.n4377 gnd.n4376 585
R3299 gnd.n2328 gnd.n1051 585
R3300 gnd.n6140 gnd.n1051 585
R3301 gnd.n4349 gnd.n4348 585
R3302 gnd.n4348 gnd.n1050 585
R3303 gnd.n4347 gnd.n2334 585
R3304 gnd.n4367 gnd.n2334 585
R3305 gnd.n4346 gnd.n4345 585
R3306 gnd.n4345 gnd.n2342 585
R3307 gnd.n4344 gnd.n2340 585
R3308 gnd.n4359 gnd.n2340 585
R3309 gnd.n4343 gnd.n4342 585
R3310 gnd.n4342 gnd.n2339 585
R3311 gnd.n4341 gnd.n2349 585
R3312 gnd.n4341 gnd.n4340 585
R3313 gnd.n4325 gnd.n2351 585
R3314 gnd.n2352 gnd.n2351 585
R3315 gnd.n4324 gnd.n2359 585
R3316 gnd.n4332 gnd.n2359 585
R3317 gnd.n4323 gnd.n4322 585
R3318 gnd.n4322 gnd.n2358 585
R3319 gnd.n4321 gnd.n2365 585
R3320 gnd.n4321 gnd.n4320 585
R3321 gnd.n4304 gnd.n2367 585
R3322 gnd.n2378 gnd.n2367 585
R3323 gnd.n4303 gnd.n2376 585
R3324 gnd.n4311 gnd.n2376 585
R3325 gnd.n4302 gnd.n4301 585
R3326 gnd.n4301 gnd.n2375 585
R3327 gnd.n4300 gnd.n2383 585
R3328 gnd.n4300 gnd.n4299 585
R3329 gnd.n4284 gnd.n2385 585
R3330 gnd.n2386 gnd.n2385 585
R3331 gnd.n4283 gnd.n2395 585
R3332 gnd.n4291 gnd.n2395 585
R3333 gnd.n4282 gnd.n4281 585
R3334 gnd.n4281 gnd.n2394 585
R3335 gnd.n4280 gnd.n2401 585
R3336 gnd.n4280 gnd.n4279 585
R3337 gnd.n4264 gnd.n2403 585
R3338 gnd.n2414 gnd.n2403 585
R3339 gnd.n4263 gnd.n2412 585
R3340 gnd.n4271 gnd.n2412 585
R3341 gnd.n4262 gnd.n4261 585
R3342 gnd.n4261 gnd.n2411 585
R3343 gnd.n4260 gnd.n2419 585
R3344 gnd.n4260 gnd.n4259 585
R3345 gnd.n4246 gnd.n2421 585
R3346 gnd.n2422 gnd.n2421 585
R3347 gnd.n4247 gnd.n2431 585
R3348 gnd.n4251 gnd.n2431 585
R3349 gnd.n4245 gnd.n4244 585
R3350 gnd.n4244 gnd.n2430 585
R3351 gnd.n6971 gnd.n6970 585
R3352 gnd.n6970 gnd.n6969 585
R3353 gnd.n6972 gnd.n156 585
R3354 gnd.n162 gnd.n156 585
R3355 gnd.n6974 gnd.n6973 585
R3356 gnd.n6975 gnd.n6974 585
R3357 gnd.n143 gnd.n142 585
R3358 gnd.n147 gnd.n143 585
R3359 gnd.n6983 gnd.n6982 585
R3360 gnd.n6982 gnd.n6981 585
R3361 gnd.n6984 gnd.n137 585
R3362 gnd.n144 gnd.n137 585
R3363 gnd.n6986 gnd.n6985 585
R3364 gnd.n6987 gnd.n6986 585
R3365 gnd.n123 gnd.n122 585
R3366 gnd.n127 gnd.n123 585
R3367 gnd.n6995 gnd.n6994 585
R3368 gnd.n6994 gnd.n6993 585
R3369 gnd.n6996 gnd.n117 585
R3370 gnd.n124 gnd.n117 585
R3371 gnd.n6998 gnd.n6997 585
R3372 gnd.n6999 gnd.n6998 585
R3373 gnd.n105 gnd.n104 585
R3374 gnd.n114 gnd.n105 585
R3375 gnd.n7007 gnd.n7006 585
R3376 gnd.n7006 gnd.n7005 585
R3377 gnd.n7008 gnd.n100 585
R3378 gnd.n100 gnd.n99 585
R3379 gnd.n7010 gnd.n7009 585
R3380 gnd.n7011 gnd.n7010 585
R3381 gnd.n84 gnd.n82 585
R3382 gnd.n88 gnd.n84 585
R3383 gnd.n7019 gnd.n7018 585
R3384 gnd.n7018 gnd.n7017 585
R3385 gnd.n83 gnd.n75 585
R3386 gnd.n85 gnd.n83 585
R3387 gnd.n7022 gnd.n73 585
R3388 gnd.n73 gnd.n70 585
R3389 gnd.n7024 gnd.n7023 585
R3390 gnd.n7025 gnd.n7024 585
R3391 gnd.n6912 gnd.n72 585
R3392 gnd.n6927 gnd.n72 585
R3393 gnd.n6914 gnd.n6913 585
R3394 gnd.n6914 gnd.n499 585
R3395 gnd.n6917 gnd.n6916 585
R3396 gnd.n6918 gnd.n6917 585
R3397 gnd.n6915 gnd.n6911 585
R3398 gnd.n6911 gnd.n6910 585
R3399 gnd.n6899 gnd.n508 585
R3400 gnd.n509 gnd.n508 585
R3401 gnd.n6901 gnd.n6900 585
R3402 gnd.n6902 gnd.n6901 585
R3403 gnd.n6898 gnd.n521 585
R3404 gnd.n6898 gnd.n6897 585
R3405 gnd.n6871 gnd.n520 585
R3406 gnd.n6883 gnd.n520 585
R3407 gnd.n6872 gnd.n541 585
R3408 gnd.n6857 gnd.n541 585
R3409 gnd.n6874 gnd.n6873 585
R3410 gnd.n6875 gnd.n6874 585
R3411 gnd.n542 gnd.n540 585
R3412 gnd.n1725 gnd.n540 585
R3413 gnd.n6866 gnd.n6865 585
R3414 gnd.n6865 gnd.n6864 585
R3415 gnd.n545 gnd.n544 585
R3416 gnd.n1732 gnd.n545 585
R3417 gnd.n1715 gnd.n1714 585
R3418 gnd.n5601 gnd.n1715 585
R3419 gnd.n5610 gnd.n5609 585
R3420 gnd.n5609 gnd.n5608 585
R3421 gnd.n5611 gnd.n1708 585
R3422 gnd.n5550 gnd.n1708 585
R3423 gnd.n5613 gnd.n5612 585
R3424 gnd.n5614 gnd.n5613 585
R3425 gnd.n1690 gnd.n1689 585
R3426 gnd.n5543 gnd.n1690 585
R3427 gnd.n5622 gnd.n5621 585
R3428 gnd.n5621 gnd.n5620 585
R3429 gnd.n5623 gnd.n1681 585
R3430 gnd.n5537 gnd.n1681 585
R3431 gnd.n5625 gnd.n5624 585
R3432 gnd.n5626 gnd.n5625 585
R3433 gnd.n1682 gnd.n1680 585
R3434 gnd.n5572 gnd.n1680 585
R3435 gnd.n1683 gnd.n1602 585
R3436 gnd.n5634 gnd.n1602 585
R3437 gnd.n5753 gnd.n5752 585
R3438 gnd.n5751 gnd.n1601 585
R3439 gnd.n5750 gnd.n1600 585
R3440 gnd.n5755 gnd.n1600 585
R3441 gnd.n5749 gnd.n5748 585
R3442 gnd.n5747 gnd.n5746 585
R3443 gnd.n5745 gnd.n5744 585
R3444 gnd.n5743 gnd.n5742 585
R3445 gnd.n5741 gnd.n5740 585
R3446 gnd.n5739 gnd.n5738 585
R3447 gnd.n5737 gnd.n5736 585
R3448 gnd.n5735 gnd.n5734 585
R3449 gnd.n5733 gnd.n5732 585
R3450 gnd.n5731 gnd.n5730 585
R3451 gnd.n5729 gnd.n5728 585
R3452 gnd.n5727 gnd.n5726 585
R3453 gnd.n5725 gnd.n5724 585
R3454 gnd.n5723 gnd.n5722 585
R3455 gnd.n5721 gnd.n5720 585
R3456 gnd.n5718 gnd.n5717 585
R3457 gnd.n5716 gnd.n5715 585
R3458 gnd.n5714 gnd.n5713 585
R3459 gnd.n5712 gnd.n5711 585
R3460 gnd.n5710 gnd.n5709 585
R3461 gnd.n5708 gnd.n5707 585
R3462 gnd.n5706 gnd.n5705 585
R3463 gnd.n5704 gnd.n5703 585
R3464 gnd.n5701 gnd.n5700 585
R3465 gnd.n5699 gnd.n5698 585
R3466 gnd.n5697 gnd.n5696 585
R3467 gnd.n5695 gnd.n5694 585
R3468 gnd.n5693 gnd.n5692 585
R3469 gnd.n5691 gnd.n5690 585
R3470 gnd.n5689 gnd.n5688 585
R3471 gnd.n5687 gnd.n5686 585
R3472 gnd.n5685 gnd.n5684 585
R3473 gnd.n5683 gnd.n5682 585
R3474 gnd.n5681 gnd.n5680 585
R3475 gnd.n5679 gnd.n5678 585
R3476 gnd.n5677 gnd.n5676 585
R3477 gnd.n5675 gnd.n5674 585
R3478 gnd.n5673 gnd.n5672 585
R3479 gnd.n5671 gnd.n5670 585
R3480 gnd.n5669 gnd.n5668 585
R3481 gnd.n5667 gnd.n5666 585
R3482 gnd.n5665 gnd.n5664 585
R3483 gnd.n5663 gnd.n5662 585
R3484 gnd.n5661 gnd.n5660 585
R3485 gnd.n5659 gnd.n5658 585
R3486 gnd.n5657 gnd.n5656 585
R3487 gnd.n5655 gnd.n5654 585
R3488 gnd.n5653 gnd.n5652 585
R3489 gnd.n5651 gnd.n5650 585
R3490 gnd.n5649 gnd.n5648 585
R3491 gnd.n5647 gnd.n5646 585
R3492 gnd.n5645 gnd.n5644 585
R3493 gnd.n5643 gnd.n5642 585
R3494 gnd.n5637 gnd.n5636 585
R3495 gnd.n491 gnd.n490 585
R3496 gnd.n488 gnd.n284 585
R3497 gnd.n487 gnd.n486 585
R3498 gnd.n480 gnd.n286 585
R3499 gnd.n482 gnd.n481 585
R3500 gnd.n478 gnd.n288 585
R3501 gnd.n477 gnd.n476 585
R3502 gnd.n470 gnd.n290 585
R3503 gnd.n472 gnd.n471 585
R3504 gnd.n468 gnd.n292 585
R3505 gnd.n467 gnd.n466 585
R3506 gnd.n460 gnd.n294 585
R3507 gnd.n462 gnd.n461 585
R3508 gnd.n458 gnd.n296 585
R3509 gnd.n457 gnd.n456 585
R3510 gnd.n450 gnd.n298 585
R3511 gnd.n452 gnd.n451 585
R3512 gnd.n448 gnd.n300 585
R3513 gnd.n447 gnd.n446 585
R3514 gnd.n440 gnd.n302 585
R3515 gnd.n442 gnd.n441 585
R3516 gnd.n438 gnd.n306 585
R3517 gnd.n437 gnd.n436 585
R3518 gnd.n430 gnd.n308 585
R3519 gnd.n432 gnd.n431 585
R3520 gnd.n428 gnd.n310 585
R3521 gnd.n427 gnd.n426 585
R3522 gnd.n420 gnd.n312 585
R3523 gnd.n422 gnd.n421 585
R3524 gnd.n418 gnd.n314 585
R3525 gnd.n417 gnd.n416 585
R3526 gnd.n410 gnd.n316 585
R3527 gnd.n412 gnd.n411 585
R3528 gnd.n408 gnd.n318 585
R3529 gnd.n407 gnd.n406 585
R3530 gnd.n400 gnd.n320 585
R3531 gnd.n402 gnd.n401 585
R3532 gnd.n398 gnd.n322 585
R3533 gnd.n397 gnd.n396 585
R3534 gnd.n390 gnd.n324 585
R3535 gnd.n392 gnd.n391 585
R3536 gnd.n388 gnd.n387 585
R3537 gnd.n386 gnd.n329 585
R3538 gnd.n380 gnd.n330 585
R3539 gnd.n382 gnd.n381 585
R3540 gnd.n377 gnd.n332 585
R3541 gnd.n376 gnd.n375 585
R3542 gnd.n369 gnd.n334 585
R3543 gnd.n371 gnd.n370 585
R3544 gnd.n367 gnd.n336 585
R3545 gnd.n366 gnd.n365 585
R3546 gnd.n359 gnd.n338 585
R3547 gnd.n361 gnd.n360 585
R3548 gnd.n357 gnd.n340 585
R3549 gnd.n356 gnd.n355 585
R3550 gnd.n349 gnd.n342 585
R3551 gnd.n351 gnd.n350 585
R3552 gnd.n347 gnd.n346 585
R3553 gnd.n345 gnd.n161 585
R3554 gnd.n165 gnd.n161 585
R3555 gnd.n6965 gnd.n163 585
R3556 gnd.n6969 gnd.n163 585
R3557 gnd.n6964 gnd.n6963 585
R3558 gnd.n6963 gnd.n162 585
R3559 gnd.n6962 gnd.n154 585
R3560 gnd.n6975 gnd.n154 585
R3561 gnd.n6961 gnd.n6960 585
R3562 gnd.n6960 gnd.n147 585
R3563 gnd.n6959 gnd.n145 585
R3564 gnd.n6981 gnd.n145 585
R3565 gnd.n6958 gnd.n6957 585
R3566 gnd.n6957 gnd.n144 585
R3567 gnd.n6955 gnd.n134 585
R3568 gnd.n6987 gnd.n134 585
R3569 gnd.n6954 gnd.n6953 585
R3570 gnd.n6953 gnd.n127 585
R3571 gnd.n6952 gnd.n125 585
R3572 gnd.n6993 gnd.n125 585
R3573 gnd.n6951 gnd.n6950 585
R3574 gnd.n6950 gnd.n124 585
R3575 gnd.n6948 gnd.n115 585
R3576 gnd.n6999 gnd.n115 585
R3577 gnd.n6947 gnd.n6946 585
R3578 gnd.n6946 gnd.n114 585
R3579 gnd.n6945 gnd.n106 585
R3580 gnd.n7005 gnd.n106 585
R3581 gnd.n6944 gnd.n6943 585
R3582 gnd.n6943 gnd.n99 585
R3583 gnd.n6941 gnd.n97 585
R3584 gnd.n7011 gnd.n97 585
R3585 gnd.n6940 gnd.n6939 585
R3586 gnd.n6939 gnd.n88 585
R3587 gnd.n6938 gnd.n86 585
R3588 gnd.n7017 gnd.n86 585
R3589 gnd.n6937 gnd.n6936 585
R3590 gnd.n6936 gnd.n85 585
R3591 gnd.n6935 gnd.n494 585
R3592 gnd.n6935 gnd.n70 585
R3593 gnd.n6924 gnd.n69 585
R3594 gnd.n7025 gnd.n69 585
R3595 gnd.n6926 gnd.n6925 585
R3596 gnd.n6927 gnd.n6926 585
R3597 gnd.n6923 gnd.n500 585
R3598 gnd.n500 gnd.n499 585
R3599 gnd.n505 gnd.n501 585
R3600 gnd.n6918 gnd.n505 585
R3601 gnd.n6888 gnd.n510 585
R3602 gnd.n6910 gnd.n510 585
R3603 gnd.n6890 gnd.n6889 585
R3604 gnd.n6889 gnd.n509 585
R3605 gnd.n6887 gnd.n518 585
R3606 gnd.n6902 gnd.n518 585
R3607 gnd.n6886 gnd.n523 585
R3608 gnd.n6897 gnd.n523 585
R3609 gnd.n6885 gnd.n6884 585
R3610 gnd.n6884 gnd.n6883 585
R3611 gnd.n530 gnd.n528 585
R3612 gnd.n6857 gnd.n530 585
R3613 gnd.n1724 gnd.n537 585
R3614 gnd.n6875 gnd.n537 585
R3615 gnd.n1727 gnd.n1726 585
R3616 gnd.n1726 gnd.n1725 585
R3617 gnd.n1728 gnd.n547 585
R3618 gnd.n6864 gnd.n547 585
R3619 gnd.n1730 gnd.n1729 585
R3620 gnd.n1732 gnd.n1730 585
R3621 gnd.n5603 gnd.n5602 585
R3622 gnd.n5602 gnd.n5601 585
R3623 gnd.n1723 gnd.n1717 585
R3624 gnd.n5608 gnd.n1717 585
R3625 gnd.n5549 gnd.n5548 585
R3626 gnd.n5550 gnd.n5549 585
R3627 gnd.n5546 gnd.n1705 585
R3628 gnd.n5614 gnd.n1705 585
R3629 gnd.n5545 gnd.n5544 585
R3630 gnd.n5544 gnd.n5543 585
R3631 gnd.n5542 gnd.n1692 585
R3632 gnd.n5620 gnd.n1692 585
R3633 gnd.n1676 gnd.n1675 585
R3634 gnd.n5537 gnd.n1676 585
R3635 gnd.n5628 gnd.n5627 585
R3636 gnd.n5627 gnd.n5626 585
R3637 gnd.n5629 gnd.n1665 585
R3638 gnd.n5572 gnd.n1665 585
R3639 gnd.n5635 gnd.n1666 585
R3640 gnd.n5635 gnd.n5634 585
R3641 gnd.n6143 gnd.n6142 585
R3642 gnd.n6142 gnd.n6141 585
R3643 gnd.n6849 gnd.n6847 585
R3644 gnd.n6849 gnd.n6848 585
R3645 gnd.n6852 gnd.n6850 585
R3646 gnd.n6850 gnd.n517 585
R3647 gnd.n6853 gnd.n558 585
R3648 gnd.n558 gnd.n522 585
R3649 gnd.n6855 gnd.n6854 585
R3650 gnd.n6856 gnd.n6855 585
R3651 gnd.n559 gnd.n557 585
R3652 gnd.n557 gnd.n538 585
R3653 gnd.n5594 gnd.n5593 585
R3654 gnd.n5594 gnd.n536 585
R3655 gnd.n5596 gnd.n5595 585
R3656 gnd.n5595 gnd.n549 585
R3657 gnd.n5597 gnd.n1734 585
R3658 gnd.n1734 gnd.n546 585
R3659 gnd.n5599 gnd.n5598 585
R3660 gnd.n5600 gnd.n5599 585
R3661 gnd.n1735 gnd.n1733 585
R3662 gnd.n1733 gnd.n1719 585
R3663 gnd.n5585 gnd.n5584 585
R3664 gnd.n5584 gnd.n1716 585
R3665 gnd.n5583 gnd.n1737 585
R3666 gnd.n5583 gnd.n1707 585
R3667 gnd.n5582 gnd.n5581 585
R3668 gnd.n5582 gnd.n1704 585
R3669 gnd.n1739 gnd.n1738 585
R3670 gnd.n1738 gnd.n1694 585
R3671 gnd.n5577 gnd.n5576 585
R3672 gnd.n5576 gnd.n1691 585
R3673 gnd.n5575 gnd.n1741 585
R3674 gnd.n5575 gnd.n1678 585
R3675 gnd.n5574 gnd.n1743 585
R3676 gnd.n5574 gnd.n5573 585
R3677 gnd.n5519 gnd.n1742 585
R3678 gnd.n1742 gnd.n1669 585
R3679 gnd.n5521 gnd.n5520 585
R3680 gnd.n5521 gnd.n1667 585
R3681 gnd.n5522 gnd.n5514 585
R3682 gnd.n5522 gnd.n1599 585
R3683 gnd.n5524 gnd.n5523 585
R3684 gnd.n5523 gnd.n1557 585
R3685 gnd.n5525 gnd.n1774 585
R3686 gnd.n1774 gnd.n1772 585
R3687 gnd.n5527 gnd.n5526 585
R3688 gnd.n5528 gnd.n5527 585
R3689 gnd.n1775 gnd.n1773 585
R3690 gnd.n1773 gnd.n1490 585
R3691 gnd.n5508 gnd.n1489 585
R3692 gnd.n5823 gnd.n1489 585
R3693 gnd.n5507 gnd.n5506 585
R3694 gnd.n5506 gnd.n1488 585
R3695 gnd.n5505 gnd.n1777 585
R3696 gnd.n5505 gnd.n5504 585
R3697 gnd.n5493 gnd.n1778 585
R3698 gnd.n5476 gnd.n1778 585
R3699 gnd.n5495 gnd.n5494 585
R3700 gnd.n5496 gnd.n5495 585
R3701 gnd.n1786 gnd.n1785 585
R3702 gnd.n5403 gnd.n1785 585
R3703 gnd.n5487 gnd.n5486 585
R3704 gnd.n5486 gnd.n5485 585
R3705 gnd.n1789 gnd.n1788 585
R3706 gnd.n5396 gnd.n1789 585
R3707 gnd.n5384 gnd.n1934 585
R3708 gnd.n5368 gnd.n1934 585
R3709 gnd.n5386 gnd.n5385 585
R3710 gnd.n5387 gnd.n5386 585
R3711 gnd.n1935 gnd.n1933 585
R3712 gnd.n1942 gnd.n1933 585
R3713 gnd.n5379 gnd.n5378 585
R3714 gnd.n5378 gnd.n5377 585
R3715 gnd.n1938 gnd.n1937 585
R3716 gnd.n1953 gnd.n1938 585
R3717 gnd.n5347 gnd.n5346 585
R3718 gnd.n5348 gnd.n5347 585
R3719 gnd.n1963 gnd.n1962 585
R3720 gnd.n5234 gnd.n1962 585
R3721 gnd.n5342 gnd.n5341 585
R3722 gnd.n5341 gnd.n5340 585
R3723 gnd.n1966 gnd.n1965 585
R3724 gnd.n1973 gnd.n1966 585
R3725 gnd.n5311 gnd.n1988 585
R3726 gnd.n1988 gnd.n1981 585
R3727 gnd.n5313 gnd.n5312 585
R3728 gnd.n5314 gnd.n5313 585
R3729 gnd.n1989 gnd.n1987 585
R3730 gnd.n1987 gnd.t45 585
R3731 gnd.n5306 gnd.n5305 585
R3732 gnd.n5305 gnd.n5304 585
R3733 gnd.n1992 gnd.n1991 585
R3734 gnd.n5296 gnd.n1992 585
R3735 gnd.n5282 gnd.n5281 585
R3736 gnd.n5283 gnd.n5282 585
R3737 gnd.n2006 gnd.n2005 585
R3738 gnd.n5260 gnd.n2005 585
R3739 gnd.n5277 gnd.n5276 585
R3740 gnd.n5276 gnd.n5275 585
R3741 gnd.n2009 gnd.n2008 585
R3742 gnd.n2019 gnd.n2009 585
R3743 gnd.n5218 gnd.n2035 585
R3744 gnd.n2035 gnd.n2017 585
R3745 gnd.n5220 gnd.n5219 585
R3746 gnd.n5221 gnd.n5220 585
R3747 gnd.n2036 gnd.n2034 585
R3748 gnd.n2043 gnd.n2034 585
R3749 gnd.n5213 gnd.n5212 585
R3750 gnd.n5212 gnd.n5211 585
R3751 gnd.n2039 gnd.n2038 585
R3752 gnd.n5197 gnd.n2039 585
R3753 gnd.n5182 gnd.n2061 585
R3754 gnd.n2061 gnd.n2060 585
R3755 gnd.n5184 gnd.n5183 585
R3756 gnd.n5185 gnd.n5184 585
R3757 gnd.n2062 gnd.n2059 585
R3758 gnd.n2069 gnd.n2059 585
R3759 gnd.n5177 gnd.n5176 585
R3760 gnd.n5176 gnd.n5175 585
R3761 gnd.n2065 gnd.n2064 585
R3762 gnd.n2074 gnd.n2065 585
R3763 gnd.n5134 gnd.n5133 585
R3764 gnd.n5135 gnd.n5134 585
R3765 gnd.n2080 gnd.n2079 585
R3766 gnd.n2088 gnd.n2079 585
R3767 gnd.n5129 gnd.n5128 585
R3768 gnd.n5128 gnd.n5127 585
R3769 gnd.n2083 gnd.n2082 585
R3770 gnd.n2094 gnd.n2083 585
R3771 gnd.n5104 gnd.n5103 585
R3772 gnd.n5105 gnd.n5104 585
R3773 gnd.n2104 gnd.n2103 585
R3774 gnd.n2103 gnd.n2099 585
R3775 gnd.n5099 gnd.n5098 585
R3776 gnd.n5098 gnd.n5097 585
R3777 gnd.n2107 gnd.n2106 585
R3778 gnd.n5089 gnd.n2107 585
R3779 gnd.n5057 gnd.n2125 585
R3780 gnd.n5016 gnd.n2125 585
R3781 gnd.n5059 gnd.n5058 585
R3782 gnd.n5060 gnd.n5059 585
R3783 gnd.n2126 gnd.n2124 585
R3784 gnd.n2133 gnd.n2124 585
R3785 gnd.n5052 gnd.n5051 585
R3786 gnd.n5051 gnd.n5050 585
R3787 gnd.n2129 gnd.n2128 585
R3788 gnd.n4909 gnd.n2129 585
R3789 gnd.n5001 gnd.n2151 585
R3790 gnd.n2151 gnd.n2144 585
R3791 gnd.n5003 gnd.n5002 585
R3792 gnd.n5004 gnd.n5003 585
R3793 gnd.n2152 gnd.n2150 585
R3794 gnd.n4905 gnd.n2150 585
R3795 gnd.n4996 gnd.n4995 585
R3796 gnd.n4995 gnd.n4994 585
R3797 gnd.n2155 gnd.n2154 585
R3798 gnd.n4986 gnd.n2155 585
R3799 gnd.n2207 gnd.n2206 585
R3800 gnd.n2207 gnd.n2168 585
R3801 gnd.n2209 gnd.n2208 585
R3802 gnd.n2208 gnd.n2167 585
R3803 gnd.n2210 gnd.n2200 585
R3804 gnd.n2200 gnd.n2172 585
R3805 gnd.n4933 gnd.n2211 585
R3806 gnd.n4933 gnd.n4932 585
R3807 gnd.n4934 gnd.n2199 585
R3808 gnd.n4934 gnd.n2176 585
R3809 gnd.n4936 gnd.n4935 585
R3810 gnd.n4935 gnd.n2180 585
R3811 gnd.n4937 gnd.n2194 585
R3812 gnd.n2194 gnd.n2185 585
R3813 gnd.n4939 gnd.n4938 585
R3814 gnd.n4940 gnd.n4939 585
R3815 gnd.n2195 gnd.n2193 585
R3816 gnd.n4851 gnd.n2193 585
R3817 gnd.n4887 gnd.n4886 585
R3818 gnd.t6 gnd.n4887 585
R3819 gnd.n2225 gnd.n2224 585
R3820 gnd.n2231 gnd.n2224 585
R3821 gnd.n4881 gnd.n4880 585
R3822 gnd.n4880 gnd.n4879 585
R3823 gnd.n2228 gnd.n2227 585
R3824 gnd.n4865 gnd.n2228 585
R3825 gnd.n4844 gnd.n4843 585
R3826 gnd.n4845 gnd.n4844 585
R3827 gnd.n4839 gnd.n4838 585
R3828 gnd.n4838 gnd.n4837 585
R3829 gnd.n1391 gnd.n1390 585
R3830 gnd.n4802 gnd.n1391 585
R3831 gnd.n5935 gnd.n5934 585
R3832 gnd.n5934 gnd.n5933 585
R3833 gnd.n5936 gnd.n1383 585
R3834 gnd.n4823 gnd.n1383 585
R3835 gnd.n5938 gnd.n5937 585
R3836 gnd.n5939 gnd.n5938 585
R3837 gnd.n1384 gnd.n1382 585
R3838 gnd.n1382 gnd.n1371 585
R3839 gnd.n1289 gnd.n1288 585
R3840 gnd.n4788 gnd.n1289 585
R3841 gnd.n5954 gnd.n5953 585
R3842 gnd.n5953 gnd.n5952 585
R3843 gnd.n5955 gnd.n1283 585
R3844 gnd.n4777 gnd.n1283 585
R3845 gnd.n5957 gnd.n5956 585
R3846 gnd.n5958 gnd.n5957 585
R3847 gnd.n1284 gnd.n1282 585
R3848 gnd.n1282 gnd.n1276 585
R3849 gnd.n4749 gnd.n4748 585
R3850 gnd.n4749 gnd.n1250 585
R3851 gnd.n4751 gnd.n4750 585
R3852 gnd.n4750 gnd.n1218 585
R3853 gnd.n4752 gnd.n2268 585
R3854 gnd.n2268 gnd.n2265 585
R3855 gnd.n4754 gnd.n4753 585
R3856 gnd.n4755 gnd.n4754 585
R3857 gnd.n2269 gnd.n2267 585
R3858 gnd.n2267 gnd.n2264 585
R3859 gnd.n4740 gnd.n4739 585
R3860 gnd.n4739 gnd.n4738 585
R3861 gnd.n2272 gnd.n2271 585
R3862 gnd.n2273 gnd.n2272 585
R3863 gnd.n4709 gnd.n4708 585
R3864 gnd.n4708 gnd.n1155 585
R3865 gnd.n4710 gnd.n2298 585
R3866 gnd.n2298 gnd.n1144 585
R3867 gnd.n4712 gnd.n4711 585
R3868 gnd.n4713 gnd.n4712 585
R3869 gnd.n2299 gnd.n2297 585
R3870 gnd.n2297 gnd.n1137 585
R3871 gnd.n4702 gnd.n4701 585
R3872 gnd.n4701 gnd.n1134 585
R3873 gnd.n4700 gnd.n2301 585
R3874 gnd.n4700 gnd.n1127 585
R3875 gnd.n4699 gnd.n4698 585
R3876 gnd.n4699 gnd.n1124 585
R3877 gnd.n2303 gnd.n2302 585
R3878 gnd.n2302 gnd.n1116 585
R3879 gnd.n4694 gnd.n4693 585
R3880 gnd.n4693 gnd.n1113 585
R3881 gnd.n4692 gnd.n2305 585
R3882 gnd.n4692 gnd.n4691 585
R3883 gnd.n4417 gnd.n2306 585
R3884 gnd.n2306 gnd.n1104 585
R3885 gnd.n4418 gnd.n2320 585
R3886 gnd.n2320 gnd.n1096 585
R3887 gnd.n4420 gnd.n4419 585
R3888 gnd.n4421 gnd.n4420 585
R3889 gnd.n2321 gnd.n2319 585
R3890 gnd.n2319 gnd.n1087 585
R3891 gnd.n4411 gnd.n4410 585
R3892 gnd.n4410 gnd.n1084 585
R3893 gnd.n4409 gnd.n2323 585
R3894 gnd.n4409 gnd.n1076 585
R3895 gnd.n4408 gnd.n4407 585
R3896 gnd.n4408 gnd.n1073 585
R3897 gnd.n4398 gnd.n4397 585
R3898 gnd.n4397 gnd.n4396 585
R3899 gnd.n4403 gnd.n4402 585
R3900 gnd.n4402 gnd.n1062 585
R3901 gnd.n4401 gnd.n1049 585
R3902 gnd.n1053 gnd.n1049 585
R3903 gnd.n5822 gnd.n5821 585
R3904 gnd.n5823 gnd.n5822 585
R3905 gnd.n1493 gnd.n1491 585
R3906 gnd.n1491 gnd.n1488 585
R3907 gnd.n5503 gnd.n5502 585
R3908 gnd.n5504 gnd.n5503 585
R3909 gnd.n1780 gnd.n1779 585
R3910 gnd.n5476 gnd.n1779 585
R3911 gnd.n5498 gnd.n5497 585
R3912 gnd.n5497 gnd.n5496 585
R3913 gnd.n1783 gnd.n1782 585
R3914 gnd.n5403 gnd.n1783 585
R3915 gnd.n1927 gnd.n1791 585
R3916 gnd.n5485 gnd.n1791 585
R3917 gnd.n5395 gnd.n5394 585
R3918 gnd.n5396 gnd.n5395 585
R3919 gnd.n1926 gnd.n1925 585
R3920 gnd.n5368 gnd.n1925 585
R3921 gnd.n5389 gnd.n5388 585
R3922 gnd.n5388 gnd.n5387 585
R3923 gnd.n1930 gnd.n1929 585
R3924 gnd.n1942 gnd.n1930 585
R3925 gnd.n5240 gnd.n1940 585
R3926 gnd.n5377 gnd.n1940 585
R3927 gnd.n5241 gnd.n5238 585
R3928 gnd.n5238 gnd.n1953 585
R3929 gnd.n5242 gnd.n1959 585
R3930 gnd.n5348 gnd.n1959 585
R3931 gnd.n5236 gnd.n5235 585
R3932 gnd.n5235 gnd.n5234 585
R3933 gnd.n5246 gnd.n1968 585
R3934 gnd.n5340 gnd.n1968 585
R3935 gnd.n5247 gnd.n5233 585
R3936 gnd.n5233 gnd.n1973 585
R3937 gnd.n5248 gnd.n5232 585
R3938 gnd.n5232 gnd.n1981 585
R3939 gnd.n5230 gnd.n1986 585
R3940 gnd.n5314 gnd.n1986 585
R3941 gnd.n5252 gnd.n5229 585
R3942 gnd.n5229 gnd.t45 585
R3943 gnd.n5253 gnd.n1993 585
R3944 gnd.n5304 gnd.n1993 585
R3945 gnd.n5254 gnd.n2000 585
R3946 gnd.n5296 gnd.n2000 585
R3947 gnd.n2026 gnd.n2004 585
R3948 gnd.n5283 gnd.n2004 585
R3949 gnd.n5259 gnd.n5258 585
R3950 gnd.n5260 gnd.n5259 585
R3951 gnd.n2025 gnd.n2012 585
R3952 gnd.n5275 gnd.n2012 585
R3953 gnd.n5225 gnd.n5224 585
R3954 gnd.n5224 gnd.n2019 585
R3955 gnd.n5223 gnd.n2028 585
R3956 gnd.n5223 gnd.n2017 585
R3957 gnd.n5222 gnd.n2030 585
R3958 gnd.n5222 gnd.n5221 585
R3959 gnd.n5191 gnd.n2029 585
R3960 gnd.n2043 gnd.n2029 585
R3961 gnd.n2053 gnd.n2041 585
R3962 gnd.n5211 gnd.n2041 585
R3963 gnd.n5196 gnd.n5195 585
R3964 gnd.n5197 gnd.n5196 585
R3965 gnd.n2052 gnd.n2051 585
R3966 gnd.n2060 gnd.n2051 585
R3967 gnd.n5187 gnd.n5186 585
R3968 gnd.n5186 gnd.n5185 585
R3969 gnd.n2056 gnd.n2055 585
R3970 gnd.n2069 gnd.n2056 585
R3971 gnd.n5072 gnd.n2066 585
R3972 gnd.n5175 gnd.n2066 585
R3973 gnd.n5075 gnd.n5071 585
R3974 gnd.n5071 gnd.n2074 585
R3975 gnd.n5076 gnd.n2078 585
R3976 gnd.n5135 gnd.n2078 585
R3977 gnd.n5077 gnd.n5070 585
R3978 gnd.n5070 gnd.n2088 585
R3979 gnd.n5068 gnd.n2085 585
R3980 gnd.n5127 gnd.n2085 585
R3981 gnd.n5081 gnd.n5067 585
R3982 gnd.n5067 gnd.n2094 585
R3983 gnd.n5082 gnd.n2101 585
R3984 gnd.n5105 gnd.n2101 585
R3985 gnd.n5083 gnd.n5066 585
R3986 gnd.n5066 gnd.n2099 585
R3987 gnd.n2117 gnd.n2109 585
R3988 gnd.n5097 gnd.n2109 585
R3989 gnd.n5088 gnd.n5087 585
R3990 gnd.n5089 gnd.n5088 585
R3991 gnd.n2116 gnd.n2115 585
R3992 gnd.n5016 gnd.n2115 585
R3993 gnd.n5062 gnd.n5061 585
R3994 gnd.n5061 gnd.n5060 585
R3995 gnd.n2120 gnd.n2119 585
R3996 gnd.n2133 gnd.n2120 585
R3997 gnd.n4912 gnd.n2131 585
R3998 gnd.n5050 gnd.n2131 585
R3999 gnd.n4911 gnd.n4910 585
R4000 gnd.n4910 gnd.n4909 585
R4001 gnd.n4916 gnd.n4907 585
R4002 gnd.n4907 gnd.n2144 585
R4003 gnd.n4917 gnd.n2149 585
R4004 gnd.n5004 gnd.n2149 585
R4005 gnd.n4918 gnd.n4906 585
R4006 gnd.n4906 gnd.n4905 585
R4007 gnd.n4903 gnd.n2156 585
R4008 gnd.n4994 gnd.n2156 585
R4009 gnd.n4922 gnd.n2164 585
R4010 gnd.n4986 gnd.n2164 585
R4011 gnd.n4923 gnd.n4902 585
R4012 gnd.n4902 gnd.n2168 585
R4013 gnd.n4924 gnd.n4901 585
R4014 gnd.n4901 gnd.n2167 585
R4015 gnd.n2215 gnd.n2213 585
R4016 gnd.n2213 gnd.n2172 585
R4017 gnd.n4929 gnd.n4928 585
R4018 gnd.n4932 gnd.n4929 585
R4019 gnd.n2214 gnd.n2212 585
R4020 gnd.n2212 gnd.n2176 585
R4021 gnd.n4897 gnd.n4896 585
R4022 gnd.n4896 gnd.n2180 585
R4023 gnd.n4895 gnd.n4894 585
R4024 gnd.n4895 gnd.n2185 585
R4025 gnd.n4893 gnd.n2190 585
R4026 gnd.n4940 gnd.n2190 585
R4027 gnd.n2221 gnd.n2217 585
R4028 gnd.n4851 gnd.n2221 585
R4029 gnd.n4889 gnd.n4888 585
R4030 gnd.n4888 gnd.t6 585
R4031 gnd.n2220 gnd.n2219 585
R4032 gnd.n2231 gnd.n2220 585
R4033 gnd.n4830 gnd.n2229 585
R4034 gnd.n4879 gnd.n2229 585
R4035 gnd.n4831 gnd.n2238 585
R4036 gnd.n4865 gnd.n2238 585
R4037 gnd.n2246 gnd.n2242 585
R4038 gnd.n4845 gnd.n2242 585
R4039 gnd.n4836 gnd.n4835 585
R4040 gnd.n4837 gnd.n4836 585
R4041 gnd.n2245 gnd.n2244 585
R4042 gnd.n4802 gnd.n2244 585
R4043 gnd.n4826 gnd.n1393 585
R4044 gnd.n5933 gnd.n1393 585
R4045 gnd.n4825 gnd.n4824 585
R4046 gnd.n4824 gnd.n4823 585
R4047 gnd.n4794 gnd.n1379 585
R4048 gnd.n5939 gnd.n1379 585
R4049 gnd.n2251 gnd.n2248 585
R4050 gnd.n2251 gnd.n1371 585
R4051 gnd.n4790 gnd.n4789 585
R4052 gnd.n4789 gnd.n4788 585
R4053 gnd.n2250 gnd.n1291 585
R4054 gnd.n5952 gnd.n1291 585
R4055 gnd.n4770 gnd.n4769 585
R4056 gnd.n4777 gnd.n4770 585
R4057 gnd.n2257 gnd.n1279 585
R4058 gnd.n5958 gnd.n1279 585
R4059 gnd.n4765 gnd.n4764 585
R4060 gnd.n4764 gnd.n1276 585
R4061 gnd.n4763 gnd.n2259 585
R4062 gnd.n4763 gnd.n1250 585
R4063 gnd.n4762 gnd.n4761 585
R4064 gnd.n4762 gnd.n1218 585
R4065 gnd.n2261 gnd.n2260 585
R4066 gnd.n2265 gnd.n2260 585
R4067 gnd.n4757 gnd.n4756 585
R4068 gnd.n4756 gnd.n4755 585
R4069 gnd.n4447 gnd.n2263 585
R4070 gnd.n4449 gnd.n4448 585
R4071 gnd.n4451 gnd.n4450 585
R4072 gnd.n4444 gnd.n4443 585
R4073 gnd.n4455 gnd.n4445 585
R4074 gnd.n4457 gnd.n4456 585
R4075 gnd.n4572 gnd.n4458 585
R4076 gnd.n4571 gnd.n4459 585
R4077 gnd.n4570 gnd.n4460 585
R4078 gnd.n4466 gnd.n4461 585
R4079 gnd.n4563 gnd.n4467 585
R4080 gnd.n4562 gnd.n4468 585
R4081 gnd.n4470 gnd.n4469 585
R4082 gnd.n4555 gnd.n4478 585
R4083 gnd.n4554 gnd.n4479 585
R4084 gnd.n4486 gnd.n4480 585
R4085 gnd.n4547 gnd.n4487 585
R4086 gnd.n4546 gnd.n4488 585
R4087 gnd.n4490 gnd.n4489 585
R4088 gnd.n4539 gnd.n4498 585
R4089 gnd.n4538 gnd.n4499 585
R4090 gnd.n4506 gnd.n4500 585
R4091 gnd.n4531 gnd.n4507 585
R4092 gnd.n4530 gnd.n4508 585
R4093 gnd.n4510 gnd.n4509 585
R4094 gnd.n4523 gnd.n4520 585
R4095 gnd.n4522 gnd.n4521 585
R4096 gnd.n2289 gnd.n2288 585
R4097 gnd.n4737 gnd.n4736 585
R4098 gnd.n4738 gnd.n4737 585
R4099 gnd.n5825 gnd.n5824 585
R4100 gnd.n5824 gnd.n5823 585
R4101 gnd.n1486 gnd.n1484 585
R4102 gnd.n1488 gnd.n1486 585
R4103 gnd.n5829 gnd.n1483 585
R4104 gnd.n5504 gnd.n1483 585
R4105 gnd.n5830 gnd.n1482 585
R4106 gnd.n5476 gnd.n1482 585
R4107 gnd.n5831 gnd.n1481 585
R4108 gnd.n5496 gnd.n1481 585
R4109 gnd.n5402 gnd.n1479 585
R4110 gnd.n5403 gnd.n5402 585
R4111 gnd.n5835 gnd.n1478 585
R4112 gnd.n5485 gnd.n1478 585
R4113 gnd.n5836 gnd.n1477 585
R4114 gnd.n5396 gnd.n1477 585
R4115 gnd.n5837 gnd.n1476 585
R4116 gnd.n5368 gnd.n1476 585
R4117 gnd.n1932 gnd.n1474 585
R4118 gnd.n5387 gnd.n1932 585
R4119 gnd.n5841 gnd.n1473 585
R4120 gnd.n1942 gnd.n1473 585
R4121 gnd.n5842 gnd.n1472 585
R4122 gnd.n5377 gnd.n1472 585
R4123 gnd.n5843 gnd.n1471 585
R4124 gnd.n1953 gnd.n1471 585
R4125 gnd.n1961 gnd.n1469 585
R4126 gnd.n5348 gnd.n1961 585
R4127 gnd.n5847 gnd.n1468 585
R4128 gnd.n5234 gnd.n1468 585
R4129 gnd.n5848 gnd.n1467 585
R4130 gnd.n5340 gnd.n1467 585
R4131 gnd.n5849 gnd.n1466 585
R4132 gnd.n1973 gnd.n1466 585
R4133 gnd.n1980 gnd.n1464 585
R4134 gnd.n1981 gnd.n1980 585
R4135 gnd.n5853 gnd.n1463 585
R4136 gnd.n5314 gnd.n1463 585
R4137 gnd.n5854 gnd.n1462 585
R4138 gnd.t45 gnd.n1462 585
R4139 gnd.n5855 gnd.n1461 585
R4140 gnd.n5304 gnd.n1461 585
R4141 gnd.n5295 gnd.n1459 585
R4142 gnd.n5296 gnd.n5295 585
R4143 gnd.n5859 gnd.n1458 585
R4144 gnd.n5283 gnd.n1458 585
R4145 gnd.n5860 gnd.n1457 585
R4146 gnd.n5260 gnd.n1457 585
R4147 gnd.n5861 gnd.n1456 585
R4148 gnd.n5275 gnd.n1456 585
R4149 gnd.n2018 gnd.n1454 585
R4150 gnd.n2019 gnd.n2018 585
R4151 gnd.n5865 gnd.n1453 585
R4152 gnd.n2017 gnd.n1453 585
R4153 gnd.n5866 gnd.n1452 585
R4154 gnd.n5221 gnd.n1452 585
R4155 gnd.n5867 gnd.n1451 585
R4156 gnd.n2043 gnd.n1451 585
R4157 gnd.n5210 gnd.n1449 585
R4158 gnd.n5211 gnd.n5210 585
R4159 gnd.n5871 gnd.n1448 585
R4160 gnd.n5197 gnd.n1448 585
R4161 gnd.n5872 gnd.n1447 585
R4162 gnd.n2060 gnd.n1447 585
R4163 gnd.n5873 gnd.n1446 585
R4164 gnd.n5185 gnd.n1446 585
R4165 gnd.n2068 gnd.n1444 585
R4166 gnd.n2069 gnd.n2068 585
R4167 gnd.n5877 gnd.n1443 585
R4168 gnd.n5175 gnd.n1443 585
R4169 gnd.n5878 gnd.n1442 585
R4170 gnd.n2074 gnd.n1442 585
R4171 gnd.n5879 gnd.n1441 585
R4172 gnd.n5135 gnd.n1441 585
R4173 gnd.n2087 gnd.n1439 585
R4174 gnd.n2088 gnd.n2087 585
R4175 gnd.n5883 gnd.n1438 585
R4176 gnd.n5127 gnd.n1438 585
R4177 gnd.n5884 gnd.n1437 585
R4178 gnd.n2094 gnd.n1437 585
R4179 gnd.n5885 gnd.n1436 585
R4180 gnd.n5105 gnd.n1436 585
R4181 gnd.n2098 gnd.n1434 585
R4182 gnd.n2099 gnd.n2098 585
R4183 gnd.n5889 gnd.n1433 585
R4184 gnd.n5097 gnd.n1433 585
R4185 gnd.n5890 gnd.n1432 585
R4186 gnd.n5089 gnd.n1432 585
R4187 gnd.n5891 gnd.n1431 585
R4188 gnd.n5016 gnd.n1431 585
R4189 gnd.n2123 gnd.n1429 585
R4190 gnd.n5060 gnd.n2123 585
R4191 gnd.n5895 gnd.n1428 585
R4192 gnd.n2133 gnd.n1428 585
R4193 gnd.n5896 gnd.n1427 585
R4194 gnd.n5050 gnd.n1427 585
R4195 gnd.n5897 gnd.n1426 585
R4196 gnd.n4909 gnd.n1426 585
R4197 gnd.n2143 gnd.n1424 585
R4198 gnd.n2144 gnd.n2143 585
R4199 gnd.n5901 gnd.n1423 585
R4200 gnd.n5004 gnd.n1423 585
R4201 gnd.n5902 gnd.n1422 585
R4202 gnd.n4905 gnd.n1422 585
R4203 gnd.n5903 gnd.n1421 585
R4204 gnd.n4994 gnd.n1421 585
R4205 gnd.n4985 gnd.n1419 585
R4206 gnd.n4986 gnd.n4985 585
R4207 gnd.n5907 gnd.n1418 585
R4208 gnd.n2168 gnd.n1418 585
R4209 gnd.n5908 gnd.n1417 585
R4210 gnd.n2167 gnd.n1417 585
R4211 gnd.n5909 gnd.n1416 585
R4212 gnd.n2172 gnd.n1416 585
R4213 gnd.n4931 gnd.n1414 585
R4214 gnd.n4932 gnd.n4931 585
R4215 gnd.n5913 gnd.n1413 585
R4216 gnd.n2176 gnd.n1413 585
R4217 gnd.n5914 gnd.n1412 585
R4218 gnd.n2180 gnd.n1412 585
R4219 gnd.n5915 gnd.n1411 585
R4220 gnd.n2185 gnd.n1411 585
R4221 gnd.n2192 gnd.n1409 585
R4222 gnd.n4940 gnd.n2192 585
R4223 gnd.n5919 gnd.n1408 585
R4224 gnd.n4851 gnd.n1408 585
R4225 gnd.n5920 gnd.n1407 585
R4226 gnd.t6 gnd.n1407 585
R4227 gnd.n5921 gnd.n1406 585
R4228 gnd.n2231 gnd.n1406 585
R4229 gnd.n4878 gnd.n1404 585
R4230 gnd.n4879 gnd.n4878 585
R4231 gnd.n5925 gnd.n1403 585
R4232 gnd.n4865 gnd.n1403 585
R4233 gnd.n5926 gnd.n1402 585
R4234 gnd.n4845 gnd.n1402 585
R4235 gnd.n5927 gnd.n1401 585
R4236 gnd.n4837 gnd.n1401 585
R4237 gnd.n1398 gnd.n1396 585
R4238 gnd.n4802 gnd.n1396 585
R4239 gnd.n5932 gnd.n5931 585
R4240 gnd.n5933 gnd.n5932 585
R4241 gnd.n1397 gnd.n1395 585
R4242 gnd.n4823 gnd.n1395 585
R4243 gnd.n4782 gnd.n1381 585
R4244 gnd.n5939 gnd.n1381 585
R4245 gnd.n2254 gnd.n2252 585
R4246 gnd.n2252 gnd.n1371 585
R4247 gnd.n4787 gnd.n4786 585
R4248 gnd.n4788 gnd.n4787 585
R4249 gnd.n2253 gnd.n1293 585
R4250 gnd.n5952 gnd.n1293 585
R4251 gnd.n4779 gnd.n4778 585
R4252 gnd.n4778 gnd.n4777 585
R4253 gnd.n2256 gnd.n1281 585
R4254 gnd.n5958 gnd.n1281 585
R4255 gnd.n4727 gnd.n4726 585
R4256 gnd.n4726 gnd.n1276 585
R4257 gnd.n4725 gnd.n4724 585
R4258 gnd.n4725 gnd.n1250 585
R4259 gnd.n4731 gnd.n4723 585
R4260 gnd.n4723 gnd.n1218 585
R4261 gnd.n4732 gnd.n4722 585
R4262 gnd.n4722 gnd.n2265 585
R4263 gnd.n4733 gnd.n2266 585
R4264 gnd.n4755 gnd.n2266 585
R4265 gnd.n5764 gnd.n1548 585
R4266 gnd.n5765 gnd.n1547 585
R4267 gnd.n1767 gnd.n1541 585
R4268 gnd.n5772 gnd.n1540 585
R4269 gnd.n5773 gnd.n1539 585
R4270 gnd.n1764 gnd.n1533 585
R4271 gnd.n5780 gnd.n1532 585
R4272 gnd.n5781 gnd.n1531 585
R4273 gnd.n1762 gnd.n1525 585
R4274 gnd.n5788 gnd.n1524 585
R4275 gnd.n5789 gnd.n1523 585
R4276 gnd.n1759 gnd.n1517 585
R4277 gnd.n5796 gnd.n1516 585
R4278 gnd.n5797 gnd.n1515 585
R4279 gnd.n1757 gnd.n1508 585
R4280 gnd.n5804 gnd.n1507 585
R4281 gnd.n5805 gnd.n1506 585
R4282 gnd.n1754 gnd.n1503 585
R4283 gnd.n5810 gnd.n1502 585
R4284 gnd.n5811 gnd.n1501 585
R4285 gnd.n5812 gnd.n1500 585
R4286 gnd.n1751 gnd.n1498 585
R4287 gnd.n5816 gnd.n1497 585
R4288 gnd.n5817 gnd.n1496 585
R4289 gnd.n5818 gnd.n1492 585
R4290 gnd.n5531 gnd.n1487 585
R4291 gnd.n5528 gnd.n1487 585
R4292 gnd.n5532 gnd.n5530 585
R4293 gnd.n1749 gnd.n1748 585
R4294 gnd.n1770 gnd.n1769 585
R4295 gnd.n5478 gnd.n1797 506.916
R4296 gnd.n5409 gnd.n1798 506.916
R4297 gnd.n1362 gnd.n1360 506.916
R4298 gnd.n6028 gnd.n1253 506.916
R4299 gnd.n1296 gnd.t167 389.64
R4300 gnd.n1920 gnd.t91 389.64
R4301 gnd.n5965 gnd.t101 389.64
R4302 gnd.n1815 gnd.t142 389.64
R4303 gnd.n6309 gnd.n878 371.755
R4304 gnd.n4517 gnd.t132 371.625
R4305 gnd.n5758 gnd.t154 371.625
R4306 gnd.n2292 gnd.t174 371.625
R4307 gnd.n1621 gnd.t151 371.625
R4308 gnd.n1644 gnd.t139 371.625
R4309 gnd.n5638 gnd.t81 371.625
R4310 gnd.n282 gnd.t88 371.625
R4311 gnd.n304 gnd.t77 371.625
R4312 gnd.n326 gnd.t145 371.625
R4313 gnd.n200 gnd.t161 371.625
R4314 gnd.n3963 gnd.t116 371.625
R4315 gnd.n3985 gnd.t98 371.625
R4316 gnd.n4006 gnd.t122 371.625
R4317 gnd.n4024 gnd.t73 371.625
R4318 gnd.n1201 gnd.t164 371.625
R4319 gnd.n4576 gnd.t105 371.625
R4320 gnd.n4589 gnd.t129 371.625
R4321 gnd.n1549 gnd.t112 371.625
R4322 gnd.n2924 gnd.t125 323.425
R4323 gnd.n2482 gnd.t157 323.425
R4324 gnd.n3773 gnd.n3747 289.615
R4325 gnd.n3741 gnd.n3715 289.615
R4326 gnd.n3709 gnd.n3683 289.615
R4327 gnd.n3678 gnd.n3652 289.615
R4328 gnd.n3646 gnd.n3620 289.615
R4329 gnd.n3614 gnd.n3588 289.615
R4330 gnd.n3582 gnd.n3556 289.615
R4331 gnd.n3551 gnd.n3525 289.615
R4332 gnd.n2998 gnd.t180 279.217
R4333 gnd.n2508 gnd.t170 279.217
R4334 gnd.n1260 gnd.t138 260.649
R4335 gnd.n1828 gnd.t150 260.649
R4336 gnd.n6030 gnd.n6029 256.663
R4337 gnd.n6030 gnd.n1219 256.663
R4338 gnd.n6030 gnd.n1220 256.663
R4339 gnd.n6030 gnd.n1221 256.663
R4340 gnd.n6030 gnd.n1222 256.663
R4341 gnd.n6030 gnd.n1223 256.663
R4342 gnd.n6030 gnd.n1224 256.663
R4343 gnd.n6030 gnd.n1225 256.663
R4344 gnd.n6030 gnd.n1226 256.663
R4345 gnd.n6030 gnd.n1227 256.663
R4346 gnd.n6030 gnd.n1228 256.663
R4347 gnd.n6030 gnd.n1229 256.663
R4348 gnd.n6030 gnd.n1230 256.663
R4349 gnd.n6030 gnd.n1231 256.663
R4350 gnd.n6030 gnd.n1232 256.663
R4351 gnd.n6030 gnd.n1233 256.663
R4352 gnd.n6033 gnd.n1216 256.663
R4353 gnd.n6031 gnd.n6030 256.663
R4354 gnd.n6030 gnd.n1234 256.663
R4355 gnd.n6030 gnd.n1235 256.663
R4356 gnd.n6030 gnd.n1236 256.663
R4357 gnd.n6030 gnd.n1237 256.663
R4358 gnd.n6030 gnd.n1238 256.663
R4359 gnd.n6030 gnd.n1239 256.663
R4360 gnd.n6030 gnd.n1240 256.663
R4361 gnd.n6030 gnd.n1241 256.663
R4362 gnd.n6030 gnd.n1242 256.663
R4363 gnd.n6030 gnd.n1243 256.663
R4364 gnd.n6030 gnd.n1244 256.663
R4365 gnd.n6030 gnd.n1245 256.663
R4366 gnd.n6030 gnd.n1246 256.663
R4367 gnd.n6030 gnd.n1247 256.663
R4368 gnd.n6030 gnd.n1248 256.663
R4369 gnd.n6030 gnd.n1249 256.663
R4370 gnd.n5475 gnd.n1903 256.663
R4371 gnd.n5475 gnd.n1904 256.663
R4372 gnd.n5475 gnd.n1905 256.663
R4373 gnd.n5475 gnd.n1906 256.663
R4374 gnd.n5475 gnd.n1907 256.663
R4375 gnd.n5475 gnd.n1908 256.663
R4376 gnd.n5475 gnd.n1909 256.663
R4377 gnd.n5475 gnd.n1910 256.663
R4378 gnd.n5475 gnd.n1911 256.663
R4379 gnd.n5475 gnd.n1912 256.663
R4380 gnd.n5475 gnd.n1913 256.663
R4381 gnd.n5475 gnd.n1914 256.663
R4382 gnd.n5475 gnd.n1915 256.663
R4383 gnd.n5475 gnd.n1916 256.663
R4384 gnd.n5475 gnd.n1917 256.663
R4385 gnd.n5475 gnd.n1918 256.663
R4386 gnd.n1919 gnd.n1631 256.663
R4387 gnd.n5475 gnd.n1902 256.663
R4388 gnd.n5475 gnd.n1814 256.663
R4389 gnd.n5475 gnd.n1813 256.663
R4390 gnd.n5475 gnd.n1812 256.663
R4391 gnd.n5475 gnd.n1811 256.663
R4392 gnd.n5475 gnd.n1810 256.663
R4393 gnd.n5475 gnd.n1809 256.663
R4394 gnd.n5475 gnd.n1808 256.663
R4395 gnd.n5475 gnd.n1807 256.663
R4396 gnd.n5475 gnd.n1806 256.663
R4397 gnd.n5475 gnd.n1805 256.663
R4398 gnd.n5475 gnd.n1804 256.663
R4399 gnd.n5475 gnd.n1803 256.663
R4400 gnd.n5475 gnd.n1802 256.663
R4401 gnd.n5475 gnd.n1801 256.663
R4402 gnd.n5475 gnd.n1800 256.663
R4403 gnd.n5475 gnd.n1799 256.663
R4404 gnd.n4241 gnd.n3933 242.672
R4405 gnd.n4241 gnd.n3934 242.672
R4406 gnd.n4241 gnd.n3935 242.672
R4407 gnd.n4241 gnd.n3936 242.672
R4408 gnd.n4241 gnd.n3937 242.672
R4409 gnd.n4241 gnd.n3938 242.672
R4410 gnd.n4241 gnd.n3939 242.672
R4411 gnd.n4241 gnd.n3940 242.672
R4412 gnd.n4241 gnd.n3941 242.672
R4413 gnd.n6084 gnd.n1154 242.672
R4414 gnd.n6084 gnd.n1153 242.672
R4415 gnd.n6084 gnd.n1152 242.672
R4416 gnd.n6084 gnd.n1151 242.672
R4417 gnd.n6084 gnd.n1150 242.672
R4418 gnd.n6084 gnd.n1149 242.672
R4419 gnd.n6084 gnd.n1148 242.672
R4420 gnd.n6084 gnd.n1147 242.672
R4421 gnd.n6084 gnd.n1146 242.672
R4422 gnd.n3052 gnd.n3051 242.672
R4423 gnd.n3052 gnd.n2962 242.672
R4424 gnd.n3052 gnd.n2963 242.672
R4425 gnd.n3052 gnd.n2964 242.672
R4426 gnd.n3052 gnd.n2965 242.672
R4427 gnd.n3052 gnd.n2966 242.672
R4428 gnd.n3052 gnd.n2967 242.672
R4429 gnd.n3052 gnd.n2968 242.672
R4430 gnd.n3052 gnd.n2969 242.672
R4431 gnd.n3052 gnd.n2970 242.672
R4432 gnd.n3052 gnd.n2971 242.672
R4433 gnd.n3052 gnd.n2972 242.672
R4434 gnd.n3053 gnd.n3052 242.672
R4435 gnd.n3905 gnd.n2457 242.672
R4436 gnd.n3905 gnd.n2456 242.672
R4437 gnd.n3905 gnd.n2455 242.672
R4438 gnd.n3905 gnd.n2454 242.672
R4439 gnd.n3905 gnd.n2453 242.672
R4440 gnd.n3905 gnd.n2452 242.672
R4441 gnd.n3905 gnd.n2451 242.672
R4442 gnd.n3905 gnd.n2450 242.672
R4443 gnd.n3905 gnd.n2449 242.672
R4444 gnd.n3905 gnd.n2448 242.672
R4445 gnd.n3905 gnd.n2447 242.672
R4446 gnd.n3905 gnd.n2446 242.672
R4447 gnd.n3905 gnd.n2445 242.672
R4448 gnd.n5755 gnd.n1586 242.672
R4449 gnd.n5755 gnd.n1588 242.672
R4450 gnd.n5755 gnd.n1589 242.672
R4451 gnd.n5755 gnd.n1591 242.672
R4452 gnd.n5755 gnd.n1593 242.672
R4453 gnd.n5755 gnd.n1594 242.672
R4454 gnd.n5755 gnd.n1596 242.672
R4455 gnd.n5755 gnd.n1598 242.672
R4456 gnd.n5756 gnd.n5755 242.672
R4457 gnd.n197 gnd.n165 242.672
R4458 gnd.n253 gnd.n165 242.672
R4459 gnd.n193 gnd.n165 242.672
R4460 gnd.n260 gnd.n165 242.672
R4461 gnd.n186 gnd.n165 242.672
R4462 gnd.n267 gnd.n165 242.672
R4463 gnd.n179 gnd.n165 242.672
R4464 gnd.n274 gnd.n165 242.672
R4465 gnd.n172 gnd.n165 242.672
R4466 gnd.n3136 gnd.n3135 242.672
R4467 gnd.n3135 gnd.n2874 242.672
R4468 gnd.n3135 gnd.n2875 242.672
R4469 gnd.n3135 gnd.n2876 242.672
R4470 gnd.n3135 gnd.n2877 242.672
R4471 gnd.n3135 gnd.n2878 242.672
R4472 gnd.n3135 gnd.n2879 242.672
R4473 gnd.n3135 gnd.n2880 242.672
R4474 gnd.n3905 gnd.n2458 242.672
R4475 gnd.n3905 gnd.n2459 242.672
R4476 gnd.n3905 gnd.n2460 242.672
R4477 gnd.n3905 gnd.n2461 242.672
R4478 gnd.n3905 gnd.n2462 242.672
R4479 gnd.n3905 gnd.n2463 242.672
R4480 gnd.n3905 gnd.n2464 242.672
R4481 gnd.n3905 gnd.n2465 242.672
R4482 gnd.n4241 gnd.n4240 242.672
R4483 gnd.n4241 gnd.n3906 242.672
R4484 gnd.n4241 gnd.n3907 242.672
R4485 gnd.n4241 gnd.n3908 242.672
R4486 gnd.n4241 gnd.n3909 242.672
R4487 gnd.n4241 gnd.n3910 242.672
R4488 gnd.n4241 gnd.n3911 242.672
R4489 gnd.n4241 gnd.n3912 242.672
R4490 gnd.n4241 gnd.n3913 242.672
R4491 gnd.n4241 gnd.n3914 242.672
R4492 gnd.n4241 gnd.n3915 242.672
R4493 gnd.n4241 gnd.n3916 242.672
R4494 gnd.n4241 gnd.n3917 242.672
R4495 gnd.n4241 gnd.n3918 242.672
R4496 gnd.n4241 gnd.n3919 242.672
R4497 gnd.n4241 gnd.n3920 242.672
R4498 gnd.n4241 gnd.n3921 242.672
R4499 gnd.n4241 gnd.n3922 242.672
R4500 gnd.n4241 gnd.n3923 242.672
R4501 gnd.n4241 gnd.n3924 242.672
R4502 gnd.n4241 gnd.n3925 242.672
R4503 gnd.n4241 gnd.n3926 242.672
R4504 gnd.n4241 gnd.n3927 242.672
R4505 gnd.n4241 gnd.n3928 242.672
R4506 gnd.n4241 gnd.n3929 242.672
R4507 gnd.n4241 gnd.n3930 242.672
R4508 gnd.n4241 gnd.n3931 242.672
R4509 gnd.n4241 gnd.n3932 242.672
R4510 gnd.n4242 gnd.n4241 242.672
R4511 gnd.n6084 gnd.n1156 242.672
R4512 gnd.n6084 gnd.n1157 242.672
R4513 gnd.n6084 gnd.n1158 242.672
R4514 gnd.n6084 gnd.n1159 242.672
R4515 gnd.n6084 gnd.n1160 242.672
R4516 gnd.n6084 gnd.n1161 242.672
R4517 gnd.n6084 gnd.n1162 242.672
R4518 gnd.n6084 gnd.n1163 242.672
R4519 gnd.n6084 gnd.n1164 242.672
R4520 gnd.n6084 gnd.n1165 242.672
R4521 gnd.n6084 gnd.n1166 242.672
R4522 gnd.n6084 gnd.n1167 242.672
R4523 gnd.n6084 gnd.n1168 242.672
R4524 gnd.n6084 gnd.n1169 242.672
R4525 gnd.n6084 gnd.n1170 242.672
R4526 gnd.n6084 gnd.n1171 242.672
R4527 gnd.n6034 gnd.n1212 242.672
R4528 gnd.n6084 gnd.n1172 242.672
R4529 gnd.n6084 gnd.n1173 242.672
R4530 gnd.n6084 gnd.n1174 242.672
R4531 gnd.n6084 gnd.n1175 242.672
R4532 gnd.n6084 gnd.n1176 242.672
R4533 gnd.n6084 gnd.n1177 242.672
R4534 gnd.n6084 gnd.n1178 242.672
R4535 gnd.n6084 gnd.n1179 242.672
R4536 gnd.n6084 gnd.n1180 242.672
R4537 gnd.n6084 gnd.n1181 242.672
R4538 gnd.n6084 gnd.n1182 242.672
R4539 gnd.n6084 gnd.n1183 242.672
R4540 gnd.n6084 gnd.n6083 242.672
R4541 gnd.n5755 gnd.n5754 242.672
R4542 gnd.n5755 gnd.n1558 242.672
R4543 gnd.n5755 gnd.n1559 242.672
R4544 gnd.n5755 gnd.n1560 242.672
R4545 gnd.n5755 gnd.n1561 242.672
R4546 gnd.n5755 gnd.n1562 242.672
R4547 gnd.n5755 gnd.n1563 242.672
R4548 gnd.n5755 gnd.n1564 242.672
R4549 gnd.n5755 gnd.n1565 242.672
R4550 gnd.n5755 gnd.n1566 242.672
R4551 gnd.n5755 gnd.n1567 242.672
R4552 gnd.n5755 gnd.n1568 242.672
R4553 gnd.n5755 gnd.n1569 242.672
R4554 gnd.n5702 gnd.n1632 242.672
R4555 gnd.n5755 gnd.n1570 242.672
R4556 gnd.n5755 gnd.n1571 242.672
R4557 gnd.n5755 gnd.n1572 242.672
R4558 gnd.n5755 gnd.n1573 242.672
R4559 gnd.n5755 gnd.n1574 242.672
R4560 gnd.n5755 gnd.n1575 242.672
R4561 gnd.n5755 gnd.n1576 242.672
R4562 gnd.n5755 gnd.n1577 242.672
R4563 gnd.n5755 gnd.n1578 242.672
R4564 gnd.n5755 gnd.n1579 242.672
R4565 gnd.n5755 gnd.n1580 242.672
R4566 gnd.n5755 gnd.n1581 242.672
R4567 gnd.n5755 gnd.n1582 242.672
R4568 gnd.n5755 gnd.n1583 242.672
R4569 gnd.n5755 gnd.n1584 242.672
R4570 gnd.n5755 gnd.n1585 242.672
R4571 gnd.n489 gnd.n165 242.672
R4572 gnd.n285 gnd.n165 242.672
R4573 gnd.n479 gnd.n165 242.672
R4574 gnd.n289 gnd.n165 242.672
R4575 gnd.n469 gnd.n165 242.672
R4576 gnd.n293 gnd.n165 242.672
R4577 gnd.n459 gnd.n165 242.672
R4578 gnd.n297 gnd.n165 242.672
R4579 gnd.n449 gnd.n165 242.672
R4580 gnd.n301 gnd.n165 242.672
R4581 gnd.n439 gnd.n165 242.672
R4582 gnd.n307 gnd.n165 242.672
R4583 gnd.n429 gnd.n165 242.672
R4584 gnd.n311 gnd.n165 242.672
R4585 gnd.n419 gnd.n165 242.672
R4586 gnd.n315 gnd.n165 242.672
R4587 gnd.n409 gnd.n165 242.672
R4588 gnd.n319 gnd.n165 242.672
R4589 gnd.n399 gnd.n165 242.672
R4590 gnd.n323 gnd.n165 242.672
R4591 gnd.n389 gnd.n165 242.672
R4592 gnd.n379 gnd.n165 242.672
R4593 gnd.n378 gnd.n165 242.672
R4594 gnd.n333 gnd.n165 242.672
R4595 gnd.n368 gnd.n165 242.672
R4596 gnd.n337 gnd.n165 242.672
R4597 gnd.n358 gnd.n165 242.672
R4598 gnd.n341 gnd.n165 242.672
R4599 gnd.n348 gnd.n165 242.672
R4600 gnd.n4738 gnd.n2274 242.672
R4601 gnd.n4738 gnd.n2275 242.672
R4602 gnd.n4738 gnd.n2276 242.672
R4603 gnd.n4738 gnd.n2277 242.672
R4604 gnd.n4738 gnd.n2278 242.672
R4605 gnd.n4738 gnd.n2279 242.672
R4606 gnd.n4738 gnd.n2280 242.672
R4607 gnd.n4738 gnd.n2281 242.672
R4608 gnd.n4738 gnd.n2282 242.672
R4609 gnd.n4738 gnd.n2283 242.672
R4610 gnd.n4738 gnd.n2284 242.672
R4611 gnd.n4738 gnd.n2285 242.672
R4612 gnd.n4738 gnd.n2286 242.672
R4613 gnd.n4738 gnd.n2287 242.672
R4614 gnd.n5528 gnd.n1771 242.672
R4615 gnd.n5528 gnd.n1768 242.672
R4616 gnd.n5528 gnd.n1766 242.672
R4617 gnd.n5528 gnd.n1765 242.672
R4618 gnd.n5528 gnd.n1763 242.672
R4619 gnd.n5528 gnd.n1761 242.672
R4620 gnd.n5528 gnd.n1760 242.672
R4621 gnd.n5528 gnd.n1758 242.672
R4622 gnd.n5528 gnd.n1756 242.672
R4623 gnd.n5528 gnd.n1755 242.672
R4624 gnd.n5528 gnd.n1753 242.672
R4625 gnd.n5528 gnd.n1752 242.672
R4626 gnd.n5528 gnd.n1750 242.672
R4627 gnd.n5529 gnd.n5528 242.672
R4628 gnd.n347 gnd.n161 240.244
R4629 gnd.n350 gnd.n349 240.244
R4630 gnd.n357 gnd.n356 240.244
R4631 gnd.n360 gnd.n359 240.244
R4632 gnd.n367 gnd.n366 240.244
R4633 gnd.n370 gnd.n369 240.244
R4634 gnd.n377 gnd.n376 240.244
R4635 gnd.n381 gnd.n380 240.244
R4636 gnd.n388 gnd.n329 240.244
R4637 gnd.n391 gnd.n390 240.244
R4638 gnd.n398 gnd.n397 240.244
R4639 gnd.n401 gnd.n400 240.244
R4640 gnd.n408 gnd.n407 240.244
R4641 gnd.n411 gnd.n410 240.244
R4642 gnd.n418 gnd.n417 240.244
R4643 gnd.n421 gnd.n420 240.244
R4644 gnd.n428 gnd.n427 240.244
R4645 gnd.n431 gnd.n430 240.244
R4646 gnd.n438 gnd.n437 240.244
R4647 gnd.n441 gnd.n440 240.244
R4648 gnd.n448 gnd.n447 240.244
R4649 gnd.n451 gnd.n450 240.244
R4650 gnd.n458 gnd.n457 240.244
R4651 gnd.n461 gnd.n460 240.244
R4652 gnd.n468 gnd.n467 240.244
R4653 gnd.n471 gnd.n470 240.244
R4654 gnd.n478 gnd.n477 240.244
R4655 gnd.n481 gnd.n480 240.244
R4656 gnd.n488 gnd.n487 240.244
R4657 gnd.n5635 gnd.n1665 240.244
R4658 gnd.n5627 gnd.n1665 240.244
R4659 gnd.n5627 gnd.n1676 240.244
R4660 gnd.n1692 gnd.n1676 240.244
R4661 gnd.n5544 gnd.n1692 240.244
R4662 gnd.n5544 gnd.n1705 240.244
R4663 gnd.n5549 gnd.n1705 240.244
R4664 gnd.n5549 gnd.n1717 240.244
R4665 gnd.n5602 gnd.n1717 240.244
R4666 gnd.n5602 gnd.n1730 240.244
R4667 gnd.n1730 gnd.n547 240.244
R4668 gnd.n1726 gnd.n547 240.244
R4669 gnd.n1726 gnd.n537 240.244
R4670 gnd.n537 gnd.n530 240.244
R4671 gnd.n6884 gnd.n530 240.244
R4672 gnd.n6884 gnd.n523 240.244
R4673 gnd.n523 gnd.n518 240.244
R4674 gnd.n6889 gnd.n518 240.244
R4675 gnd.n6889 gnd.n510 240.244
R4676 gnd.n510 gnd.n505 240.244
R4677 gnd.n505 gnd.n500 240.244
R4678 gnd.n6926 gnd.n500 240.244
R4679 gnd.n6926 gnd.n69 240.244
R4680 gnd.n6935 gnd.n69 240.244
R4681 gnd.n6936 gnd.n6935 240.244
R4682 gnd.n6936 gnd.n86 240.244
R4683 gnd.n6939 gnd.n86 240.244
R4684 gnd.n6939 gnd.n97 240.244
R4685 gnd.n6943 gnd.n97 240.244
R4686 gnd.n6943 gnd.n106 240.244
R4687 gnd.n6946 gnd.n106 240.244
R4688 gnd.n6946 gnd.n115 240.244
R4689 gnd.n6950 gnd.n115 240.244
R4690 gnd.n6950 gnd.n125 240.244
R4691 gnd.n6953 gnd.n125 240.244
R4692 gnd.n6953 gnd.n134 240.244
R4693 gnd.n6957 gnd.n134 240.244
R4694 gnd.n6957 gnd.n145 240.244
R4695 gnd.n6960 gnd.n145 240.244
R4696 gnd.n6960 gnd.n154 240.244
R4697 gnd.n6963 gnd.n154 240.244
R4698 gnd.n6963 gnd.n163 240.244
R4699 gnd.n1601 gnd.n1600 240.244
R4700 gnd.n5748 gnd.n1600 240.244
R4701 gnd.n5746 gnd.n5745 240.244
R4702 gnd.n5742 gnd.n5741 240.244
R4703 gnd.n5738 gnd.n5737 240.244
R4704 gnd.n5734 gnd.n5733 240.244
R4705 gnd.n5730 gnd.n5729 240.244
R4706 gnd.n5726 gnd.n5725 240.244
R4707 gnd.n5722 gnd.n5721 240.244
R4708 gnd.n5717 gnd.n5716 240.244
R4709 gnd.n5713 gnd.n5712 240.244
R4710 gnd.n5709 gnd.n5708 240.244
R4711 gnd.n5705 gnd.n5704 240.244
R4712 gnd.n5700 gnd.n5699 240.244
R4713 gnd.n5696 gnd.n5695 240.244
R4714 gnd.n5692 gnd.n5691 240.244
R4715 gnd.n5688 gnd.n5687 240.244
R4716 gnd.n5684 gnd.n5683 240.244
R4717 gnd.n5680 gnd.n5679 240.244
R4718 gnd.n5676 gnd.n5675 240.244
R4719 gnd.n5672 gnd.n5671 240.244
R4720 gnd.n5668 gnd.n5667 240.244
R4721 gnd.n5664 gnd.n5663 240.244
R4722 gnd.n5660 gnd.n5659 240.244
R4723 gnd.n5656 gnd.n5655 240.244
R4724 gnd.n5652 gnd.n5651 240.244
R4725 gnd.n5648 gnd.n5647 240.244
R4726 gnd.n5644 gnd.n5643 240.244
R4727 gnd.n1680 gnd.n1602 240.244
R4728 gnd.n5625 gnd.n1680 240.244
R4729 gnd.n5625 gnd.n1681 240.244
R4730 gnd.n5621 gnd.n1681 240.244
R4731 gnd.n5621 gnd.n1690 240.244
R4732 gnd.n5613 gnd.n1690 240.244
R4733 gnd.n5613 gnd.n1708 240.244
R4734 gnd.n5609 gnd.n1708 240.244
R4735 gnd.n5609 gnd.n1715 240.244
R4736 gnd.n1715 gnd.n545 240.244
R4737 gnd.n6865 gnd.n545 240.244
R4738 gnd.n6865 gnd.n540 240.244
R4739 gnd.n6874 gnd.n540 240.244
R4740 gnd.n6874 gnd.n541 240.244
R4741 gnd.n541 gnd.n520 240.244
R4742 gnd.n6898 gnd.n520 240.244
R4743 gnd.n6901 gnd.n6898 240.244
R4744 gnd.n6901 gnd.n508 240.244
R4745 gnd.n6911 gnd.n508 240.244
R4746 gnd.n6917 gnd.n6911 240.244
R4747 gnd.n6917 gnd.n6914 240.244
R4748 gnd.n6914 gnd.n72 240.244
R4749 gnd.n7024 gnd.n72 240.244
R4750 gnd.n7024 gnd.n73 240.244
R4751 gnd.n83 gnd.n73 240.244
R4752 gnd.n7018 gnd.n83 240.244
R4753 gnd.n7018 gnd.n84 240.244
R4754 gnd.n7010 gnd.n84 240.244
R4755 gnd.n7010 gnd.n100 240.244
R4756 gnd.n7006 gnd.n100 240.244
R4757 gnd.n7006 gnd.n105 240.244
R4758 gnd.n6998 gnd.n105 240.244
R4759 gnd.n6998 gnd.n117 240.244
R4760 gnd.n6994 gnd.n117 240.244
R4761 gnd.n6994 gnd.n123 240.244
R4762 gnd.n6986 gnd.n123 240.244
R4763 gnd.n6986 gnd.n137 240.244
R4764 gnd.n6982 gnd.n137 240.244
R4765 gnd.n6982 gnd.n143 240.244
R4766 gnd.n6974 gnd.n143 240.244
R4767 gnd.n6974 gnd.n156 240.244
R4768 gnd.n6970 gnd.n156 240.244
R4769 gnd.n6085 gnd.n1143 240.244
R4770 gnd.n6082 gnd.n1184 240.244
R4771 gnd.n6078 gnd.n6077 240.244
R4772 gnd.n6074 gnd.n6073 240.244
R4773 gnd.n6070 gnd.n6069 240.244
R4774 gnd.n6066 gnd.n6065 240.244
R4775 gnd.n6062 gnd.n6061 240.244
R4776 gnd.n6058 gnd.n6057 240.244
R4777 gnd.n6054 gnd.n6053 240.244
R4778 gnd.n6049 gnd.n6048 240.244
R4779 gnd.n6045 gnd.n6044 240.244
R4780 gnd.n6041 gnd.n6040 240.244
R4781 gnd.n6037 gnd.n6036 240.244
R4782 gnd.n4598 gnd.n4597 240.244
R4783 gnd.n4601 gnd.n4600 240.244
R4784 gnd.n4608 gnd.n4607 240.244
R4785 gnd.n4611 gnd.n4610 240.244
R4786 gnd.n4616 gnd.n4591 240.244
R4787 gnd.n4620 gnd.n4619 240.244
R4788 gnd.n4627 gnd.n4626 240.244
R4789 gnd.n4630 gnd.n4629 240.244
R4790 gnd.n4637 gnd.n4636 240.244
R4791 gnd.n4640 gnd.n4639 240.244
R4792 gnd.n4647 gnd.n4646 240.244
R4793 gnd.n4650 gnd.n4649 240.244
R4794 gnd.n4657 gnd.n4656 240.244
R4795 gnd.n4660 gnd.n4659 240.244
R4796 gnd.n4665 gnd.n4578 240.244
R4797 gnd.n4244 gnd.n2431 240.244
R4798 gnd.n2431 gnd.n2421 240.244
R4799 gnd.n4260 gnd.n2421 240.244
R4800 gnd.n4261 gnd.n4260 240.244
R4801 gnd.n4261 gnd.n2412 240.244
R4802 gnd.n2412 gnd.n2403 240.244
R4803 gnd.n4280 gnd.n2403 240.244
R4804 gnd.n4281 gnd.n4280 240.244
R4805 gnd.n4281 gnd.n2395 240.244
R4806 gnd.n2395 gnd.n2385 240.244
R4807 gnd.n4300 gnd.n2385 240.244
R4808 gnd.n4301 gnd.n4300 240.244
R4809 gnd.n4301 gnd.n2376 240.244
R4810 gnd.n2376 gnd.n2367 240.244
R4811 gnd.n4321 gnd.n2367 240.244
R4812 gnd.n4322 gnd.n4321 240.244
R4813 gnd.n4322 gnd.n2359 240.244
R4814 gnd.n2359 gnd.n2351 240.244
R4815 gnd.n4341 gnd.n2351 240.244
R4816 gnd.n4342 gnd.n4341 240.244
R4817 gnd.n4342 gnd.n2340 240.244
R4818 gnd.n4345 gnd.n2340 240.244
R4819 gnd.n4345 gnd.n2334 240.244
R4820 gnd.n4348 gnd.n2334 240.244
R4821 gnd.n4348 gnd.n1051 240.244
R4822 gnd.n4377 gnd.n1051 240.244
R4823 gnd.n4377 gnd.n1063 240.244
R4824 gnd.n2324 gnd.n1063 240.244
R4825 gnd.n2324 gnd.n1074 240.244
R4826 gnd.n4386 gnd.n1074 240.244
R4827 gnd.n4386 gnd.n1085 240.244
R4828 gnd.n2318 gnd.n1085 240.244
R4829 gnd.n2318 gnd.n1094 240.244
R4830 gnd.n4431 gnd.n1094 240.244
R4831 gnd.n4431 gnd.n1105 240.244
R4832 gnd.n2307 gnd.n1105 240.244
R4833 gnd.n2307 gnd.n1114 240.244
R4834 gnd.n4438 gnd.n1114 240.244
R4835 gnd.n4438 gnd.n1125 240.244
R4836 gnd.n4676 gnd.n1125 240.244
R4837 gnd.n4676 gnd.n1135 240.244
R4838 gnd.n2296 gnd.n1135 240.244
R4839 gnd.n3944 gnd.n3943 240.244
R4840 gnd.n4234 gnd.n3943 240.244
R4841 gnd.n4232 gnd.n4231 240.244
R4842 gnd.n4228 gnd.n4227 240.244
R4843 gnd.n4224 gnd.n4223 240.244
R4844 gnd.n4220 gnd.n4219 240.244
R4845 gnd.n4216 gnd.n4215 240.244
R4846 gnd.n4212 gnd.n4211 240.244
R4847 gnd.n4208 gnd.n4207 240.244
R4848 gnd.n4203 gnd.n4202 240.244
R4849 gnd.n4199 gnd.n4198 240.244
R4850 gnd.n4195 gnd.n4194 240.244
R4851 gnd.n4191 gnd.n4190 240.244
R4852 gnd.n4187 gnd.n4186 240.244
R4853 gnd.n4183 gnd.n4182 240.244
R4854 gnd.n4179 gnd.n4178 240.244
R4855 gnd.n4175 gnd.n4174 240.244
R4856 gnd.n4171 gnd.n4170 240.244
R4857 gnd.n4167 gnd.n4166 240.244
R4858 gnd.n4163 gnd.n4162 240.244
R4859 gnd.n4159 gnd.n4158 240.244
R4860 gnd.n4155 gnd.n4154 240.244
R4861 gnd.n4151 gnd.n4150 240.244
R4862 gnd.n4147 gnd.n4146 240.244
R4863 gnd.n4143 gnd.n4142 240.244
R4864 gnd.n4139 gnd.n4138 240.244
R4865 gnd.n4135 gnd.n4134 240.244
R4866 gnd.n4131 gnd.n4130 240.244
R4867 gnd.n4127 gnd.n2442 240.244
R4868 gnd.n4252 gnd.n2429 240.244
R4869 gnd.n4252 gnd.n2425 240.244
R4870 gnd.n4258 gnd.n2425 240.244
R4871 gnd.n4258 gnd.n2410 240.244
R4872 gnd.n4272 gnd.n2410 240.244
R4873 gnd.n4272 gnd.n2406 240.244
R4874 gnd.n4278 gnd.n2406 240.244
R4875 gnd.n4278 gnd.n2393 240.244
R4876 gnd.n4292 gnd.n2393 240.244
R4877 gnd.n4292 gnd.n2389 240.244
R4878 gnd.n4298 gnd.n2389 240.244
R4879 gnd.n4298 gnd.n2374 240.244
R4880 gnd.n4312 gnd.n2374 240.244
R4881 gnd.n4312 gnd.n2370 240.244
R4882 gnd.n4319 gnd.n2370 240.244
R4883 gnd.n4319 gnd.n2357 240.244
R4884 gnd.n4333 gnd.n2357 240.244
R4885 gnd.n4333 gnd.n2355 240.244
R4886 gnd.n4339 gnd.n2355 240.244
R4887 gnd.n4339 gnd.n2338 240.244
R4888 gnd.n4360 gnd.n2338 240.244
R4889 gnd.n4360 gnd.n2336 240.244
R4890 gnd.n4366 gnd.n2336 240.244
R4891 gnd.n4366 gnd.n1055 240.244
R4892 gnd.n6139 gnd.n1055 240.244
R4893 gnd.n6139 gnd.n1056 240.244
R4894 gnd.n6135 gnd.n1056 240.244
R4895 gnd.n6135 gnd.n1061 240.244
R4896 gnd.n6127 gnd.n1061 240.244
R4897 gnd.n6127 gnd.n1077 240.244
R4898 gnd.n6123 gnd.n1077 240.244
R4899 gnd.n6123 gnd.n1083 240.244
R4900 gnd.n6115 gnd.n1083 240.244
R4901 gnd.n6115 gnd.n1097 240.244
R4902 gnd.n6111 gnd.n1097 240.244
R4903 gnd.n6111 gnd.n1103 240.244
R4904 gnd.n6103 gnd.n1103 240.244
R4905 gnd.n6103 gnd.n1117 240.244
R4906 gnd.n6099 gnd.n1117 240.244
R4907 gnd.n6099 gnd.n1123 240.244
R4908 gnd.n6091 gnd.n1123 240.244
R4909 gnd.n6091 gnd.n1138 240.244
R4910 gnd.n3904 gnd.n2467 240.244
R4911 gnd.n3897 gnd.n3896 240.244
R4912 gnd.n3894 gnd.n3893 240.244
R4913 gnd.n3890 gnd.n3889 240.244
R4914 gnd.n3886 gnd.n3885 240.244
R4915 gnd.n3882 gnd.n3881 240.244
R4916 gnd.n3878 gnd.n3877 240.244
R4917 gnd.n3874 gnd.n3873 240.244
R4918 gnd.n3147 gnd.n2859 240.244
R4919 gnd.n3157 gnd.n2859 240.244
R4920 gnd.n3157 gnd.n2850 240.244
R4921 gnd.n2850 gnd.n2839 240.244
R4922 gnd.n3178 gnd.n2839 240.244
R4923 gnd.n3178 gnd.n2833 240.244
R4924 gnd.n3188 gnd.n2833 240.244
R4925 gnd.n3188 gnd.n2822 240.244
R4926 gnd.n2822 gnd.n2814 240.244
R4927 gnd.n3206 gnd.n2814 240.244
R4928 gnd.n3207 gnd.n3206 240.244
R4929 gnd.n3207 gnd.n2799 240.244
R4930 gnd.n3209 gnd.n2799 240.244
R4931 gnd.n3209 gnd.n2785 240.244
R4932 gnd.n3251 gnd.n2785 240.244
R4933 gnd.n3252 gnd.n3251 240.244
R4934 gnd.n3255 gnd.n3252 240.244
R4935 gnd.n3255 gnd.n2740 240.244
R4936 gnd.n2780 gnd.n2740 240.244
R4937 gnd.n2780 gnd.n2750 240.244
R4938 gnd.n3265 gnd.n2750 240.244
R4939 gnd.n3265 gnd.n2771 240.244
R4940 gnd.n3275 gnd.n2771 240.244
R4941 gnd.n3275 gnd.n2669 240.244
R4942 gnd.n3320 gnd.n2669 240.244
R4943 gnd.n3320 gnd.n2655 240.244
R4944 gnd.n3342 gnd.n2655 240.244
R4945 gnd.n3343 gnd.n3342 240.244
R4946 gnd.n3343 gnd.n2642 240.244
R4947 gnd.n2642 gnd.n2631 240.244
R4948 gnd.n3374 gnd.n2631 240.244
R4949 gnd.n3375 gnd.n3374 240.244
R4950 gnd.n3376 gnd.n3375 240.244
R4951 gnd.n3376 gnd.n2616 240.244
R4952 gnd.n2616 gnd.n2615 240.244
R4953 gnd.n2615 gnd.n2600 240.244
R4954 gnd.n3427 gnd.n2600 240.244
R4955 gnd.n3428 gnd.n3427 240.244
R4956 gnd.n3428 gnd.n2587 240.244
R4957 gnd.n2587 gnd.n2576 240.244
R4958 gnd.n3459 gnd.n2576 240.244
R4959 gnd.n3460 gnd.n3459 240.244
R4960 gnd.n3461 gnd.n3460 240.244
R4961 gnd.n3461 gnd.n2560 240.244
R4962 gnd.n2560 gnd.n2559 240.244
R4963 gnd.n2559 gnd.n2546 240.244
R4964 gnd.n3516 gnd.n2546 240.244
R4965 gnd.n3517 gnd.n3516 240.244
R4966 gnd.n3517 gnd.n2533 240.244
R4967 gnd.n2533 gnd.n2523 240.244
R4968 gnd.n3805 gnd.n2523 240.244
R4969 gnd.n3808 gnd.n3805 240.244
R4970 gnd.n3808 gnd.n3807 240.244
R4971 gnd.n3137 gnd.n2872 240.244
R4972 gnd.n2893 gnd.n2872 240.244
R4973 gnd.n2896 gnd.n2895 240.244
R4974 gnd.n2903 gnd.n2902 240.244
R4975 gnd.n2906 gnd.n2905 240.244
R4976 gnd.n2913 gnd.n2912 240.244
R4977 gnd.n2916 gnd.n2915 240.244
R4978 gnd.n2923 gnd.n2922 240.244
R4979 gnd.n3145 gnd.n2869 240.244
R4980 gnd.n2869 gnd.n2848 240.244
R4981 gnd.n3168 gnd.n2848 240.244
R4982 gnd.n3168 gnd.n2842 240.244
R4983 gnd.n3176 gnd.n2842 240.244
R4984 gnd.n3176 gnd.n2844 240.244
R4985 gnd.n2844 gnd.n2820 240.244
R4986 gnd.n3198 gnd.n2820 240.244
R4987 gnd.n3198 gnd.n2816 240.244
R4988 gnd.n3204 gnd.n2816 240.244
R4989 gnd.n3204 gnd.n2798 240.244
R4990 gnd.n3229 gnd.n2798 240.244
R4991 gnd.n3229 gnd.n2793 240.244
R4992 gnd.n3241 gnd.n2793 240.244
R4993 gnd.n3241 gnd.n2794 240.244
R4994 gnd.n3237 gnd.n2794 240.244
R4995 gnd.n3237 gnd.n2742 240.244
R4996 gnd.n3289 gnd.n2742 240.244
R4997 gnd.n3289 gnd.n2743 240.244
R4998 gnd.n3285 gnd.n2743 240.244
R4999 gnd.n3285 gnd.n2749 240.244
R5000 gnd.n2769 gnd.n2749 240.244
R5001 gnd.n2769 gnd.n2667 240.244
R5002 gnd.n3324 gnd.n2667 240.244
R5003 gnd.n3324 gnd.n2662 240.244
R5004 gnd.n3332 gnd.n2662 240.244
R5005 gnd.n3332 gnd.n2663 240.244
R5006 gnd.n2663 gnd.n2640 240.244
R5007 gnd.n3364 gnd.n2640 240.244
R5008 gnd.n3364 gnd.n2635 240.244
R5009 gnd.n3372 gnd.n2635 240.244
R5010 gnd.n3372 gnd.n2636 240.244
R5011 gnd.n2636 gnd.n2613 240.244
R5012 gnd.n3409 gnd.n2613 240.244
R5013 gnd.n3409 gnd.n2608 240.244
R5014 gnd.n3417 gnd.n2608 240.244
R5015 gnd.n3417 gnd.n2609 240.244
R5016 gnd.n2609 gnd.n2585 240.244
R5017 gnd.n3449 gnd.n2585 240.244
R5018 gnd.n3449 gnd.n2580 240.244
R5019 gnd.n3457 gnd.n2580 240.244
R5020 gnd.n3457 gnd.n2581 240.244
R5021 gnd.n2581 gnd.n2558 240.244
R5022 gnd.n3498 gnd.n2558 240.244
R5023 gnd.n3498 gnd.n2553 240.244
R5024 gnd.n3506 gnd.n2553 240.244
R5025 gnd.n3506 gnd.n2554 240.244
R5026 gnd.n2554 gnd.n2531 240.244
R5027 gnd.n3793 gnd.n2531 240.244
R5028 gnd.n3793 gnd.n2526 240.244
R5029 gnd.n3803 gnd.n2526 240.244
R5030 gnd.n3803 gnd.n2527 240.244
R5031 gnd.n2527 gnd.n2466 240.244
R5032 gnd.n169 gnd.n166 240.244
R5033 gnd.n276 gnd.n275 240.244
R5034 gnd.n273 gnd.n173 240.244
R5035 gnd.n269 gnd.n268 240.244
R5036 gnd.n266 gnd.n180 240.244
R5037 gnd.n262 gnd.n261 240.244
R5038 gnd.n259 gnd.n187 240.244
R5039 gnd.n255 gnd.n254 240.244
R5040 gnd.n252 gnd.n194 240.244
R5041 gnd.n5571 gnd.n1668 240.244
R5042 gnd.n5571 gnd.n1677 240.244
R5043 gnd.n5538 gnd.n1677 240.244
R5044 gnd.n5538 gnd.n1693 240.244
R5045 gnd.n5539 gnd.n1693 240.244
R5046 gnd.n5539 gnd.n1706 240.244
R5047 gnd.n5551 gnd.n1706 240.244
R5048 gnd.n5551 gnd.n1718 240.244
R5049 gnd.n1731 gnd.n1718 240.244
R5050 gnd.n5552 gnd.n1731 240.244
R5051 gnd.n5552 gnd.n548 240.244
R5052 gnd.n548 gnd.n535 240.244
R5053 gnd.n6876 gnd.n535 240.244
R5054 gnd.n6876 gnd.n531 240.244
R5055 gnd.n6882 gnd.n531 240.244
R5056 gnd.n6882 gnd.n516 240.244
R5057 gnd.n6903 gnd.n516 240.244
R5058 gnd.n6903 gnd.n511 240.244
R5059 gnd.n6909 gnd.n511 240.244
R5060 gnd.n6909 gnd.n507 240.244
R5061 gnd.n507 gnd.n506 240.244
R5062 gnd.n506 gnd.n66 240.244
R5063 gnd.n7026 gnd.n66 240.244
R5064 gnd.n7026 gnd.n68 240.244
R5065 gnd.n216 gnd.n68 240.244
R5066 gnd.n216 gnd.n87 240.244
R5067 gnd.n212 gnd.n87 240.244
R5068 gnd.n212 gnd.n98 240.244
R5069 gnd.n223 gnd.n98 240.244
R5070 gnd.n223 gnd.n107 240.244
R5071 gnd.n209 gnd.n107 240.244
R5072 gnd.n209 gnd.n116 240.244
R5073 gnd.n230 gnd.n116 240.244
R5074 gnd.n230 gnd.n126 240.244
R5075 gnd.n206 gnd.n126 240.244
R5076 gnd.n206 gnd.n135 240.244
R5077 gnd.n237 gnd.n135 240.244
R5078 gnd.n237 gnd.n146 240.244
R5079 gnd.n203 gnd.n146 240.244
R5080 gnd.n203 gnd.n155 240.244
R5081 gnd.n244 gnd.n155 240.244
R5082 gnd.n244 gnd.n164 240.244
R5083 gnd.n1512 gnd.n1511 240.244
R5084 gnd.n1587 gnd.n1519 240.244
R5085 gnd.n1590 gnd.n1520 240.244
R5086 gnd.n1528 gnd.n1527 240.244
R5087 gnd.n1592 gnd.n1535 240.244
R5088 gnd.n1595 gnd.n1536 240.244
R5089 gnd.n1544 gnd.n1543 240.244
R5090 gnd.n1597 gnd.n1553 240.244
R5091 gnd.n5757 gnd.n1556 240.244
R5092 gnd.n5633 gnd.n1671 240.244
R5093 gnd.n1679 gnd.n1671 240.244
R5094 gnd.n1695 gnd.n1679 240.244
R5095 gnd.n5619 gnd.n1695 240.244
R5096 gnd.n5619 gnd.n1696 240.244
R5097 gnd.n5615 gnd.n1696 240.244
R5098 gnd.n5615 gnd.n1703 240.244
R5099 gnd.n5607 gnd.n1703 240.244
R5100 gnd.n5607 gnd.n1720 240.244
R5101 gnd.n1720 gnd.n550 240.244
R5102 gnd.n6863 gnd.n550 240.244
R5103 gnd.n6863 gnd.n551 240.244
R5104 gnd.n551 gnd.n539 240.244
R5105 gnd.n6858 gnd.n539 240.244
R5106 gnd.n6858 gnd.n524 240.244
R5107 gnd.n6896 gnd.n524 240.244
R5108 gnd.n6896 gnd.n519 240.244
R5109 gnd.n6892 gnd.n519 240.244
R5110 gnd.n6892 gnd.n504 240.244
R5111 gnd.n6919 gnd.n504 240.244
R5112 gnd.n6919 gnd.n498 240.244
R5113 gnd.n6928 gnd.n498 240.244
R5114 gnd.n6928 gnd.n71 240.244
R5115 gnd.n6931 gnd.n71 240.244
R5116 gnd.n6931 gnd.n89 240.244
R5117 gnd.n7016 gnd.n89 240.244
R5118 gnd.n7016 gnd.n90 240.244
R5119 gnd.n7012 gnd.n90 240.244
R5120 gnd.n7012 gnd.n96 240.244
R5121 gnd.n7004 gnd.n96 240.244
R5122 gnd.n7004 gnd.n108 240.244
R5123 gnd.n7000 gnd.n108 240.244
R5124 gnd.n7000 gnd.n113 240.244
R5125 gnd.n6992 gnd.n113 240.244
R5126 gnd.n6992 gnd.n128 240.244
R5127 gnd.n6988 gnd.n128 240.244
R5128 gnd.n6988 gnd.n133 240.244
R5129 gnd.n6980 gnd.n133 240.244
R5130 gnd.n6980 gnd.n148 240.244
R5131 gnd.n6976 gnd.n148 240.244
R5132 gnd.n6976 gnd.n153 240.244
R5133 gnd.n6968 gnd.n153 240.244
R5134 gnd.n2486 gnd.n2444 240.244
R5135 gnd.n3864 gnd.n3863 240.244
R5136 gnd.n3860 gnd.n3859 240.244
R5137 gnd.n3856 gnd.n3855 240.244
R5138 gnd.n3852 gnd.n3851 240.244
R5139 gnd.n3848 gnd.n3847 240.244
R5140 gnd.n3844 gnd.n3843 240.244
R5141 gnd.n3840 gnd.n3839 240.244
R5142 gnd.n3836 gnd.n3835 240.244
R5143 gnd.n3832 gnd.n3831 240.244
R5144 gnd.n3828 gnd.n3827 240.244
R5145 gnd.n3824 gnd.n3823 240.244
R5146 gnd.n3820 gnd.n3819 240.244
R5147 gnd.n3060 gnd.n2957 240.244
R5148 gnd.n3060 gnd.n2950 240.244
R5149 gnd.n3071 gnd.n2950 240.244
R5150 gnd.n3071 gnd.n2946 240.244
R5151 gnd.n3077 gnd.n2946 240.244
R5152 gnd.n3077 gnd.n2938 240.244
R5153 gnd.n3087 gnd.n2938 240.244
R5154 gnd.n3087 gnd.n2933 240.244
R5155 gnd.n3123 gnd.n2933 240.244
R5156 gnd.n3123 gnd.n2934 240.244
R5157 gnd.n2934 gnd.n2881 240.244
R5158 gnd.n3118 gnd.n2881 240.244
R5159 gnd.n3118 gnd.n3117 240.244
R5160 gnd.n3117 gnd.n2860 240.244
R5161 gnd.n3113 gnd.n2860 240.244
R5162 gnd.n3113 gnd.n2851 240.244
R5163 gnd.n3110 gnd.n2851 240.244
R5164 gnd.n3110 gnd.n3109 240.244
R5165 gnd.n3109 gnd.n2834 240.244
R5166 gnd.n3105 gnd.n2834 240.244
R5167 gnd.n3105 gnd.n2823 240.244
R5168 gnd.n2823 gnd.n2804 240.244
R5169 gnd.n3218 gnd.n2804 240.244
R5170 gnd.n3218 gnd.n2800 240.244
R5171 gnd.n3226 gnd.n2800 240.244
R5172 gnd.n3226 gnd.n2791 240.244
R5173 gnd.n2791 gnd.n2727 240.244
R5174 gnd.n3298 gnd.n2727 240.244
R5175 gnd.n3298 gnd.n2728 240.244
R5176 gnd.n2739 gnd.n2728 240.244
R5177 gnd.n2774 gnd.n2739 240.244
R5178 gnd.n2777 gnd.n2774 240.244
R5179 gnd.n2777 gnd.n2751 240.244
R5180 gnd.n2764 gnd.n2751 240.244
R5181 gnd.n2764 gnd.n2761 240.244
R5182 gnd.n2761 gnd.n2670 240.244
R5183 gnd.n3319 gnd.n2670 240.244
R5184 gnd.n3319 gnd.n2660 240.244
R5185 gnd.n3315 gnd.n2660 240.244
R5186 gnd.n3315 gnd.n2654 240.244
R5187 gnd.n3312 gnd.n2654 240.244
R5188 gnd.n3312 gnd.n2643 240.244
R5189 gnd.n3309 gnd.n2643 240.244
R5190 gnd.n3309 gnd.n2621 240.244
R5191 gnd.n3385 gnd.n2621 240.244
R5192 gnd.n3385 gnd.n2617 240.244
R5193 gnd.n3406 gnd.n2617 240.244
R5194 gnd.n3406 gnd.n2606 240.244
R5195 gnd.n3402 gnd.n2606 240.244
R5196 gnd.n3402 gnd.n2599 240.244
R5197 gnd.n3399 gnd.n2599 240.244
R5198 gnd.n3399 gnd.n2588 240.244
R5199 gnd.n3396 gnd.n2588 240.244
R5200 gnd.n3396 gnd.n2565 240.244
R5201 gnd.n3470 gnd.n2565 240.244
R5202 gnd.n3470 gnd.n2561 240.244
R5203 gnd.n3495 gnd.n2561 240.244
R5204 gnd.n3495 gnd.n2552 240.244
R5205 gnd.n3491 gnd.n2552 240.244
R5206 gnd.n3491 gnd.n2545 240.244
R5207 gnd.n3487 gnd.n2545 240.244
R5208 gnd.n3487 gnd.n2534 240.244
R5209 gnd.n3484 gnd.n2534 240.244
R5210 gnd.n3484 gnd.n2515 240.244
R5211 gnd.n3815 gnd.n2515 240.244
R5212 gnd.n2974 gnd.n2973 240.244
R5213 gnd.n3045 gnd.n2973 240.244
R5214 gnd.n3043 gnd.n3042 240.244
R5215 gnd.n3039 gnd.n3038 240.244
R5216 gnd.n3035 gnd.n3034 240.244
R5217 gnd.n3031 gnd.n3030 240.244
R5218 gnd.n3027 gnd.n3026 240.244
R5219 gnd.n3023 gnd.n3022 240.244
R5220 gnd.n3019 gnd.n3018 240.244
R5221 gnd.n3015 gnd.n3014 240.244
R5222 gnd.n3011 gnd.n3010 240.244
R5223 gnd.n3007 gnd.n3006 240.244
R5224 gnd.n3003 gnd.n2961 240.244
R5225 gnd.n3063 gnd.n2955 240.244
R5226 gnd.n3063 gnd.n2951 240.244
R5227 gnd.n3069 gnd.n2951 240.244
R5228 gnd.n3069 gnd.n2944 240.244
R5229 gnd.n3079 gnd.n2944 240.244
R5230 gnd.n3079 gnd.n2940 240.244
R5231 gnd.n3085 gnd.n2940 240.244
R5232 gnd.n3085 gnd.n2931 240.244
R5233 gnd.n3125 gnd.n2931 240.244
R5234 gnd.n3125 gnd.n2882 240.244
R5235 gnd.n3133 gnd.n2882 240.244
R5236 gnd.n3133 gnd.n2883 240.244
R5237 gnd.n2883 gnd.n2861 240.244
R5238 gnd.n3154 gnd.n2861 240.244
R5239 gnd.n3154 gnd.n2853 240.244
R5240 gnd.n3165 gnd.n2853 240.244
R5241 gnd.n3165 gnd.n2854 240.244
R5242 gnd.n2854 gnd.n2835 240.244
R5243 gnd.n3185 gnd.n2835 240.244
R5244 gnd.n3185 gnd.n2825 240.244
R5245 gnd.n3195 gnd.n2825 240.244
R5246 gnd.n3195 gnd.n2806 240.244
R5247 gnd.n3216 gnd.n2806 240.244
R5248 gnd.n3216 gnd.n2808 240.244
R5249 gnd.n2808 gnd.n2789 240.244
R5250 gnd.n3244 gnd.n2789 240.244
R5251 gnd.n3244 gnd.n2731 240.244
R5252 gnd.n3296 gnd.n2731 240.244
R5253 gnd.n3296 gnd.n2732 240.244
R5254 gnd.n3292 gnd.n2732 240.244
R5255 gnd.n3292 gnd.n2738 240.244
R5256 gnd.n2753 gnd.n2738 240.244
R5257 gnd.n3282 gnd.n2753 240.244
R5258 gnd.n3282 gnd.n2754 240.244
R5259 gnd.n3278 gnd.n2754 240.244
R5260 gnd.n3278 gnd.n2760 240.244
R5261 gnd.n2760 gnd.n2659 240.244
R5262 gnd.n3335 gnd.n2659 240.244
R5263 gnd.n3335 gnd.n2652 240.244
R5264 gnd.n3346 gnd.n2652 240.244
R5265 gnd.n3346 gnd.n2645 240.244
R5266 gnd.n3361 gnd.n2645 240.244
R5267 gnd.n3361 gnd.n2646 240.244
R5268 gnd.n2646 gnd.n2624 240.244
R5269 gnd.n3383 gnd.n2624 240.244
R5270 gnd.n3383 gnd.n2625 240.244
R5271 gnd.n2625 gnd.n2604 240.244
R5272 gnd.n3420 gnd.n2604 240.244
R5273 gnd.n3420 gnd.n2597 240.244
R5274 gnd.n3431 gnd.n2597 240.244
R5275 gnd.n3431 gnd.n2590 240.244
R5276 gnd.n3446 gnd.n2590 240.244
R5277 gnd.n3446 gnd.n2591 240.244
R5278 gnd.n2591 gnd.n2568 240.244
R5279 gnd.n3468 gnd.n2568 240.244
R5280 gnd.n3468 gnd.n2570 240.244
R5281 gnd.n2570 gnd.n2550 240.244
R5282 gnd.n3509 gnd.n2550 240.244
R5283 gnd.n3509 gnd.n2543 240.244
R5284 gnd.n3521 gnd.n2543 240.244
R5285 gnd.n3521 gnd.n2536 240.244
R5286 gnd.n3790 gnd.n2536 240.244
R5287 gnd.n3790 gnd.n2537 240.244
R5288 gnd.n2537 gnd.n2518 240.244
R5289 gnd.n3813 gnd.n2518 240.244
R5290 gnd.n4463 gnd.n1145 240.244
R5291 gnd.n4473 gnd.n4472 240.244
R5292 gnd.n4475 gnd.n4474 240.244
R5293 gnd.n4483 gnd.n4482 240.244
R5294 gnd.n4493 gnd.n4492 240.244
R5295 gnd.n4495 gnd.n4494 240.244
R5296 gnd.n4503 gnd.n4502 240.244
R5297 gnd.n4513 gnd.n4512 240.244
R5298 gnd.n4515 gnd.n4514 240.244
R5299 gnd.n4081 gnd.n2432 240.244
R5300 gnd.n4078 gnd.n2432 240.244
R5301 gnd.n4078 gnd.n2423 240.244
R5302 gnd.n4075 gnd.n2423 240.244
R5303 gnd.n4075 gnd.n2413 240.244
R5304 gnd.n4072 gnd.n2413 240.244
R5305 gnd.n4072 gnd.n2404 240.244
R5306 gnd.n4069 gnd.n2404 240.244
R5307 gnd.n4069 gnd.n2396 240.244
R5308 gnd.n4066 gnd.n2396 240.244
R5309 gnd.n4066 gnd.n2387 240.244
R5310 gnd.n4063 gnd.n2387 240.244
R5311 gnd.n4063 gnd.n2377 240.244
R5312 gnd.n4060 gnd.n2377 240.244
R5313 gnd.n4060 gnd.n2368 240.244
R5314 gnd.n4057 gnd.n2368 240.244
R5315 gnd.n4057 gnd.n2360 240.244
R5316 gnd.n4054 gnd.n2360 240.244
R5317 gnd.n4054 gnd.n2353 240.244
R5318 gnd.n4051 gnd.n2353 240.244
R5319 gnd.n4051 gnd.n2341 240.244
R5320 gnd.n2341 gnd.n2333 240.244
R5321 gnd.n4368 gnd.n2333 240.244
R5322 gnd.n4369 gnd.n4368 240.244
R5323 gnd.n4369 gnd.n1052 240.244
R5324 gnd.n4375 gnd.n1052 240.244
R5325 gnd.n4375 gnd.n1064 240.244
R5326 gnd.n4394 gnd.n1064 240.244
R5327 gnd.n4394 gnd.n1075 240.244
R5328 gnd.n4388 gnd.n1075 240.244
R5329 gnd.n4388 gnd.n1086 240.244
R5330 gnd.n4423 gnd.n1086 240.244
R5331 gnd.n4423 gnd.n1095 240.244
R5332 gnd.n4429 gnd.n1095 240.244
R5333 gnd.n4429 gnd.n1106 240.244
R5334 gnd.n4689 gnd.n1106 240.244
R5335 gnd.n4689 gnd.n1115 240.244
R5336 gnd.n2312 gnd.n1115 240.244
R5337 gnd.n2312 gnd.n1126 240.244
R5338 gnd.n4678 gnd.n1126 240.244
R5339 gnd.n4678 gnd.n1136 240.244
R5340 gnd.n4715 gnd.n1136 240.244
R5341 gnd.n4118 gnd.n4117 240.244
R5342 gnd.n4114 gnd.n4113 240.244
R5343 gnd.n4110 gnd.n4109 240.244
R5344 gnd.n4106 gnd.n4105 240.244
R5345 gnd.n4102 gnd.n4101 240.244
R5346 gnd.n4098 gnd.n4097 240.244
R5347 gnd.n4094 gnd.n4093 240.244
R5348 gnd.n4090 gnd.n4089 240.244
R5349 gnd.n4023 gnd.n3942 240.244
R5350 gnd.n4250 gnd.n2433 240.244
R5351 gnd.n4250 gnd.n2434 240.244
R5352 gnd.n2434 gnd.n2424 240.244
R5353 gnd.n2424 gnd.n2415 240.244
R5354 gnd.n4270 gnd.n2415 240.244
R5355 gnd.n4270 gnd.n2416 240.244
R5356 gnd.n2416 gnd.n2405 240.244
R5357 gnd.n2405 gnd.n2397 240.244
R5358 gnd.n4290 gnd.n2397 240.244
R5359 gnd.n4290 gnd.n2398 240.244
R5360 gnd.n2398 gnd.n2388 240.244
R5361 gnd.n2388 gnd.n2379 240.244
R5362 gnd.n4310 gnd.n2379 240.244
R5363 gnd.n4310 gnd.n2380 240.244
R5364 gnd.n2380 gnd.n2369 240.244
R5365 gnd.n2369 gnd.n2361 240.244
R5366 gnd.n4331 gnd.n2361 240.244
R5367 gnd.n4331 gnd.n2362 240.244
R5368 gnd.n2362 gnd.n2354 240.244
R5369 gnd.n2354 gnd.n2343 240.244
R5370 gnd.n4358 gnd.n2343 240.244
R5371 gnd.n4358 gnd.n2344 240.244
R5372 gnd.n2344 gnd.n2335 240.244
R5373 gnd.n4353 gnd.n2335 240.244
R5374 gnd.n4353 gnd.n1054 240.244
R5375 gnd.n1065 gnd.n1054 240.244
R5376 gnd.n6133 gnd.n1065 240.244
R5377 gnd.n6133 gnd.n1066 240.244
R5378 gnd.n6129 gnd.n1066 240.244
R5379 gnd.n6129 gnd.n1072 240.244
R5380 gnd.n6121 gnd.n1072 240.244
R5381 gnd.n6121 gnd.n1088 240.244
R5382 gnd.n6117 gnd.n1088 240.244
R5383 gnd.n6117 gnd.n1093 240.244
R5384 gnd.n6109 gnd.n1093 240.244
R5385 gnd.n6109 gnd.n1107 240.244
R5386 gnd.n6105 gnd.n1107 240.244
R5387 gnd.n6105 gnd.n1112 240.244
R5388 gnd.n6097 gnd.n1112 240.244
R5389 gnd.n6097 gnd.n1128 240.244
R5390 gnd.n6093 gnd.n1128 240.244
R5391 gnd.n6093 gnd.n1133 240.244
R5392 gnd.n6316 gnd.n879 240.244
R5393 gnd.n6316 gnd.n877 240.244
R5394 gnd.n6320 gnd.n877 240.244
R5395 gnd.n6320 gnd.n873 240.244
R5396 gnd.n6326 gnd.n873 240.244
R5397 gnd.n6326 gnd.n871 240.244
R5398 gnd.n6330 gnd.n871 240.244
R5399 gnd.n6330 gnd.n867 240.244
R5400 gnd.n6336 gnd.n867 240.244
R5401 gnd.n6336 gnd.n865 240.244
R5402 gnd.n6340 gnd.n865 240.244
R5403 gnd.n6340 gnd.n861 240.244
R5404 gnd.n6346 gnd.n861 240.244
R5405 gnd.n6346 gnd.n859 240.244
R5406 gnd.n6350 gnd.n859 240.244
R5407 gnd.n6350 gnd.n855 240.244
R5408 gnd.n6356 gnd.n855 240.244
R5409 gnd.n6356 gnd.n853 240.244
R5410 gnd.n6360 gnd.n853 240.244
R5411 gnd.n6360 gnd.n849 240.244
R5412 gnd.n6366 gnd.n849 240.244
R5413 gnd.n6366 gnd.n847 240.244
R5414 gnd.n6370 gnd.n847 240.244
R5415 gnd.n6370 gnd.n843 240.244
R5416 gnd.n6376 gnd.n843 240.244
R5417 gnd.n6376 gnd.n841 240.244
R5418 gnd.n6380 gnd.n841 240.244
R5419 gnd.n6380 gnd.n837 240.244
R5420 gnd.n6386 gnd.n837 240.244
R5421 gnd.n6386 gnd.n835 240.244
R5422 gnd.n6390 gnd.n835 240.244
R5423 gnd.n6390 gnd.n831 240.244
R5424 gnd.n6396 gnd.n831 240.244
R5425 gnd.n6396 gnd.n829 240.244
R5426 gnd.n6400 gnd.n829 240.244
R5427 gnd.n6400 gnd.n825 240.244
R5428 gnd.n6406 gnd.n825 240.244
R5429 gnd.n6406 gnd.n823 240.244
R5430 gnd.n6410 gnd.n823 240.244
R5431 gnd.n6410 gnd.n819 240.244
R5432 gnd.n6416 gnd.n819 240.244
R5433 gnd.n6416 gnd.n817 240.244
R5434 gnd.n6420 gnd.n817 240.244
R5435 gnd.n6420 gnd.n813 240.244
R5436 gnd.n6426 gnd.n813 240.244
R5437 gnd.n6426 gnd.n811 240.244
R5438 gnd.n6430 gnd.n811 240.244
R5439 gnd.n6430 gnd.n807 240.244
R5440 gnd.n6436 gnd.n807 240.244
R5441 gnd.n6436 gnd.n805 240.244
R5442 gnd.n6440 gnd.n805 240.244
R5443 gnd.n6440 gnd.n801 240.244
R5444 gnd.n6446 gnd.n801 240.244
R5445 gnd.n6446 gnd.n799 240.244
R5446 gnd.n6450 gnd.n799 240.244
R5447 gnd.n6450 gnd.n795 240.244
R5448 gnd.n6456 gnd.n795 240.244
R5449 gnd.n6456 gnd.n793 240.244
R5450 gnd.n6460 gnd.n793 240.244
R5451 gnd.n6460 gnd.n789 240.244
R5452 gnd.n6466 gnd.n789 240.244
R5453 gnd.n6466 gnd.n787 240.244
R5454 gnd.n6470 gnd.n787 240.244
R5455 gnd.n6470 gnd.n783 240.244
R5456 gnd.n6476 gnd.n783 240.244
R5457 gnd.n6476 gnd.n781 240.244
R5458 gnd.n6480 gnd.n781 240.244
R5459 gnd.n6480 gnd.n777 240.244
R5460 gnd.n6486 gnd.n777 240.244
R5461 gnd.n6486 gnd.n775 240.244
R5462 gnd.n6490 gnd.n775 240.244
R5463 gnd.n6490 gnd.n771 240.244
R5464 gnd.n6496 gnd.n771 240.244
R5465 gnd.n6496 gnd.n769 240.244
R5466 gnd.n6500 gnd.n769 240.244
R5467 gnd.n6500 gnd.n765 240.244
R5468 gnd.n6506 gnd.n765 240.244
R5469 gnd.n6506 gnd.n763 240.244
R5470 gnd.n6510 gnd.n763 240.244
R5471 gnd.n6510 gnd.n759 240.244
R5472 gnd.n6516 gnd.n759 240.244
R5473 gnd.n6516 gnd.n757 240.244
R5474 gnd.n6520 gnd.n757 240.244
R5475 gnd.n6520 gnd.n753 240.244
R5476 gnd.n6526 gnd.n753 240.244
R5477 gnd.n6526 gnd.n751 240.244
R5478 gnd.n6530 gnd.n751 240.244
R5479 gnd.n6530 gnd.n747 240.244
R5480 gnd.n6536 gnd.n747 240.244
R5481 gnd.n6536 gnd.n745 240.244
R5482 gnd.n6540 gnd.n745 240.244
R5483 gnd.n6540 gnd.n741 240.244
R5484 gnd.n6546 gnd.n741 240.244
R5485 gnd.n6546 gnd.n739 240.244
R5486 gnd.n6550 gnd.n739 240.244
R5487 gnd.n6550 gnd.n735 240.244
R5488 gnd.n6556 gnd.n735 240.244
R5489 gnd.n6556 gnd.n733 240.244
R5490 gnd.n6560 gnd.n733 240.244
R5491 gnd.n6560 gnd.n729 240.244
R5492 gnd.n6566 gnd.n729 240.244
R5493 gnd.n6566 gnd.n727 240.244
R5494 gnd.n6570 gnd.n727 240.244
R5495 gnd.n6570 gnd.n723 240.244
R5496 gnd.n6576 gnd.n723 240.244
R5497 gnd.n6576 gnd.n721 240.244
R5498 gnd.n6580 gnd.n721 240.244
R5499 gnd.n6580 gnd.n717 240.244
R5500 gnd.n6586 gnd.n717 240.244
R5501 gnd.n6586 gnd.n715 240.244
R5502 gnd.n6590 gnd.n715 240.244
R5503 gnd.n6590 gnd.n711 240.244
R5504 gnd.n6596 gnd.n711 240.244
R5505 gnd.n6596 gnd.n709 240.244
R5506 gnd.n6600 gnd.n709 240.244
R5507 gnd.n6600 gnd.n705 240.244
R5508 gnd.n6606 gnd.n705 240.244
R5509 gnd.n6606 gnd.n703 240.244
R5510 gnd.n6610 gnd.n703 240.244
R5511 gnd.n6610 gnd.n699 240.244
R5512 gnd.n6616 gnd.n699 240.244
R5513 gnd.n6616 gnd.n697 240.244
R5514 gnd.n6620 gnd.n697 240.244
R5515 gnd.n6620 gnd.n693 240.244
R5516 gnd.n6627 gnd.n693 240.244
R5517 gnd.n6627 gnd.n691 240.244
R5518 gnd.n6631 gnd.n691 240.244
R5519 gnd.n6631 gnd.n688 240.244
R5520 gnd.n6637 gnd.n686 240.244
R5521 gnd.n6641 gnd.n686 240.244
R5522 gnd.n6641 gnd.n682 240.244
R5523 gnd.n6647 gnd.n682 240.244
R5524 gnd.n6647 gnd.n680 240.244
R5525 gnd.n6651 gnd.n680 240.244
R5526 gnd.n6651 gnd.n676 240.244
R5527 gnd.n6657 gnd.n676 240.244
R5528 gnd.n6657 gnd.n674 240.244
R5529 gnd.n6661 gnd.n674 240.244
R5530 gnd.n6661 gnd.n670 240.244
R5531 gnd.n6667 gnd.n670 240.244
R5532 gnd.n6667 gnd.n668 240.244
R5533 gnd.n6671 gnd.n668 240.244
R5534 gnd.n6671 gnd.n664 240.244
R5535 gnd.n6677 gnd.n664 240.244
R5536 gnd.n6677 gnd.n662 240.244
R5537 gnd.n6681 gnd.n662 240.244
R5538 gnd.n6681 gnd.n658 240.244
R5539 gnd.n6687 gnd.n658 240.244
R5540 gnd.n6687 gnd.n656 240.244
R5541 gnd.n6691 gnd.n656 240.244
R5542 gnd.n6691 gnd.n652 240.244
R5543 gnd.n6697 gnd.n652 240.244
R5544 gnd.n6697 gnd.n650 240.244
R5545 gnd.n6701 gnd.n650 240.244
R5546 gnd.n6701 gnd.n646 240.244
R5547 gnd.n6707 gnd.n646 240.244
R5548 gnd.n6707 gnd.n644 240.244
R5549 gnd.n6711 gnd.n644 240.244
R5550 gnd.n6711 gnd.n640 240.244
R5551 gnd.n6717 gnd.n640 240.244
R5552 gnd.n6717 gnd.n638 240.244
R5553 gnd.n6721 gnd.n638 240.244
R5554 gnd.n6721 gnd.n634 240.244
R5555 gnd.n6727 gnd.n634 240.244
R5556 gnd.n6727 gnd.n632 240.244
R5557 gnd.n6731 gnd.n632 240.244
R5558 gnd.n6731 gnd.n628 240.244
R5559 gnd.n6737 gnd.n628 240.244
R5560 gnd.n6737 gnd.n626 240.244
R5561 gnd.n6741 gnd.n626 240.244
R5562 gnd.n6741 gnd.n622 240.244
R5563 gnd.n6747 gnd.n622 240.244
R5564 gnd.n6747 gnd.n620 240.244
R5565 gnd.n6751 gnd.n620 240.244
R5566 gnd.n6751 gnd.n616 240.244
R5567 gnd.n6757 gnd.n616 240.244
R5568 gnd.n6757 gnd.n614 240.244
R5569 gnd.n6761 gnd.n614 240.244
R5570 gnd.n6761 gnd.n610 240.244
R5571 gnd.n6767 gnd.n610 240.244
R5572 gnd.n6767 gnd.n608 240.244
R5573 gnd.n6771 gnd.n608 240.244
R5574 gnd.n6771 gnd.n604 240.244
R5575 gnd.n6777 gnd.n604 240.244
R5576 gnd.n6777 gnd.n602 240.244
R5577 gnd.n6781 gnd.n602 240.244
R5578 gnd.n6781 gnd.n598 240.244
R5579 gnd.n6787 gnd.n598 240.244
R5580 gnd.n6787 gnd.n596 240.244
R5581 gnd.n6791 gnd.n596 240.244
R5582 gnd.n6791 gnd.n592 240.244
R5583 gnd.n6797 gnd.n592 240.244
R5584 gnd.n6797 gnd.n590 240.244
R5585 gnd.n6801 gnd.n590 240.244
R5586 gnd.n6801 gnd.n586 240.244
R5587 gnd.n6807 gnd.n586 240.244
R5588 gnd.n6807 gnd.n584 240.244
R5589 gnd.n6811 gnd.n584 240.244
R5590 gnd.n6811 gnd.n580 240.244
R5591 gnd.n6817 gnd.n580 240.244
R5592 gnd.n6817 gnd.n578 240.244
R5593 gnd.n6821 gnd.n578 240.244
R5594 gnd.n6821 gnd.n574 240.244
R5595 gnd.n6827 gnd.n574 240.244
R5596 gnd.n6827 gnd.n572 240.244
R5597 gnd.n6831 gnd.n572 240.244
R5598 gnd.n6831 gnd.n568 240.244
R5599 gnd.n6837 gnd.n568 240.244
R5600 gnd.n6837 gnd.n566 240.244
R5601 gnd.n6842 gnd.n566 240.244
R5602 gnd.n6842 gnd.n562 240.244
R5603 gnd.n6849 gnd.n562 240.244
R5604 gnd.n4402 gnd.n1049 240.244
R5605 gnd.n4402 gnd.n4397 240.244
R5606 gnd.n4408 gnd.n4397 240.244
R5607 gnd.n4409 gnd.n4408 240.244
R5608 gnd.n4410 gnd.n4409 240.244
R5609 gnd.n4410 gnd.n2319 240.244
R5610 gnd.n4420 gnd.n2319 240.244
R5611 gnd.n4420 gnd.n2320 240.244
R5612 gnd.n2320 gnd.n2306 240.244
R5613 gnd.n4692 gnd.n2306 240.244
R5614 gnd.n4693 gnd.n4692 240.244
R5615 gnd.n4693 gnd.n2302 240.244
R5616 gnd.n4699 gnd.n2302 240.244
R5617 gnd.n4700 gnd.n4699 240.244
R5618 gnd.n4701 gnd.n4700 240.244
R5619 gnd.n4701 gnd.n2297 240.244
R5620 gnd.n4712 gnd.n2297 240.244
R5621 gnd.n4712 gnd.n2298 240.244
R5622 gnd.n4708 gnd.n2298 240.244
R5623 gnd.n4708 gnd.n2272 240.244
R5624 gnd.n4739 gnd.n2272 240.244
R5625 gnd.n4739 gnd.n2267 240.244
R5626 gnd.n4754 gnd.n2267 240.244
R5627 gnd.n4754 gnd.n2268 240.244
R5628 gnd.n4750 gnd.n2268 240.244
R5629 gnd.n4750 gnd.n4749 240.244
R5630 gnd.n4749 gnd.n1282 240.244
R5631 gnd.n5957 gnd.n1282 240.244
R5632 gnd.n5957 gnd.n1283 240.244
R5633 gnd.n5953 gnd.n1283 240.244
R5634 gnd.n5953 gnd.n1289 240.244
R5635 gnd.n1382 gnd.n1289 240.244
R5636 gnd.n5938 gnd.n1382 240.244
R5637 gnd.n5938 gnd.n1383 240.244
R5638 gnd.n5934 gnd.n1383 240.244
R5639 gnd.n5934 gnd.n1391 240.244
R5640 gnd.n4838 gnd.n1391 240.244
R5641 gnd.n4844 gnd.n4838 240.244
R5642 gnd.n4844 gnd.n2228 240.244
R5643 gnd.n4880 gnd.n2228 240.244
R5644 gnd.n4880 gnd.n2224 240.244
R5645 gnd.n4887 gnd.n2224 240.244
R5646 gnd.n4887 gnd.n2193 240.244
R5647 gnd.n4939 gnd.n2193 240.244
R5648 gnd.n4939 gnd.n2194 240.244
R5649 gnd.n4935 gnd.n2194 240.244
R5650 gnd.n4935 gnd.n4934 240.244
R5651 gnd.n4934 gnd.n4933 240.244
R5652 gnd.n4933 gnd.n2200 240.244
R5653 gnd.n2208 gnd.n2200 240.244
R5654 gnd.n2208 gnd.n2207 240.244
R5655 gnd.n2207 gnd.n2155 240.244
R5656 gnd.n4995 gnd.n2155 240.244
R5657 gnd.n4995 gnd.n2150 240.244
R5658 gnd.n5003 gnd.n2150 240.244
R5659 gnd.n5003 gnd.n2151 240.244
R5660 gnd.n2151 gnd.n2129 240.244
R5661 gnd.n5051 gnd.n2129 240.244
R5662 gnd.n5051 gnd.n2124 240.244
R5663 gnd.n5059 gnd.n2124 240.244
R5664 gnd.n5059 gnd.n2125 240.244
R5665 gnd.n2125 gnd.n2107 240.244
R5666 gnd.n5098 gnd.n2107 240.244
R5667 gnd.n5098 gnd.n2103 240.244
R5668 gnd.n5104 gnd.n2103 240.244
R5669 gnd.n5104 gnd.n2083 240.244
R5670 gnd.n5128 gnd.n2083 240.244
R5671 gnd.n5128 gnd.n2079 240.244
R5672 gnd.n5134 gnd.n2079 240.244
R5673 gnd.n5134 gnd.n2065 240.244
R5674 gnd.n5176 gnd.n2065 240.244
R5675 gnd.n5176 gnd.n2059 240.244
R5676 gnd.n5184 gnd.n2059 240.244
R5677 gnd.n5184 gnd.n2061 240.244
R5678 gnd.n2061 gnd.n2039 240.244
R5679 gnd.n5212 gnd.n2039 240.244
R5680 gnd.n5212 gnd.n2034 240.244
R5681 gnd.n5220 gnd.n2034 240.244
R5682 gnd.n5220 gnd.n2035 240.244
R5683 gnd.n2035 gnd.n2009 240.244
R5684 gnd.n5276 gnd.n2009 240.244
R5685 gnd.n5276 gnd.n2005 240.244
R5686 gnd.n5282 gnd.n2005 240.244
R5687 gnd.n5282 gnd.n1992 240.244
R5688 gnd.n5305 gnd.n1992 240.244
R5689 gnd.n5305 gnd.n1987 240.244
R5690 gnd.n5313 gnd.n1987 240.244
R5691 gnd.n5313 gnd.n1988 240.244
R5692 gnd.n1988 gnd.n1966 240.244
R5693 gnd.n5341 gnd.n1966 240.244
R5694 gnd.n5341 gnd.n1962 240.244
R5695 gnd.n5347 gnd.n1962 240.244
R5696 gnd.n5347 gnd.n1938 240.244
R5697 gnd.n5378 gnd.n1938 240.244
R5698 gnd.n5378 gnd.n1933 240.244
R5699 gnd.n5386 gnd.n1933 240.244
R5700 gnd.n5386 gnd.n1934 240.244
R5701 gnd.n1934 gnd.n1789 240.244
R5702 gnd.n5486 gnd.n1789 240.244
R5703 gnd.n5486 gnd.n1785 240.244
R5704 gnd.n5495 gnd.n1785 240.244
R5705 gnd.n5495 gnd.n1778 240.244
R5706 gnd.n5505 gnd.n1778 240.244
R5707 gnd.n5506 gnd.n5505 240.244
R5708 gnd.n5506 gnd.n1489 240.244
R5709 gnd.n1773 gnd.n1489 240.244
R5710 gnd.n5527 gnd.n1773 240.244
R5711 gnd.n5527 gnd.n1774 240.244
R5712 gnd.n5523 gnd.n1774 240.244
R5713 gnd.n5523 gnd.n5522 240.244
R5714 gnd.n5522 gnd.n5521 240.244
R5715 gnd.n5521 gnd.n1742 240.244
R5716 gnd.n5574 gnd.n1742 240.244
R5717 gnd.n5575 gnd.n5574 240.244
R5718 gnd.n5576 gnd.n5575 240.244
R5719 gnd.n5576 gnd.n1738 240.244
R5720 gnd.n5582 gnd.n1738 240.244
R5721 gnd.n5583 gnd.n5582 240.244
R5722 gnd.n5584 gnd.n5583 240.244
R5723 gnd.n5584 gnd.n1733 240.244
R5724 gnd.n5599 gnd.n1733 240.244
R5725 gnd.n5599 gnd.n1734 240.244
R5726 gnd.n5595 gnd.n1734 240.244
R5727 gnd.n5595 gnd.n5594 240.244
R5728 gnd.n5594 gnd.n557 240.244
R5729 gnd.n6855 gnd.n557 240.244
R5730 gnd.n6855 gnd.n558 240.244
R5731 gnd.n6850 gnd.n558 240.244
R5732 gnd.n6310 gnd.n883 240.244
R5733 gnd.n6306 gnd.n883 240.244
R5734 gnd.n6306 gnd.n885 240.244
R5735 gnd.n6302 gnd.n885 240.244
R5736 gnd.n6302 gnd.n890 240.244
R5737 gnd.n6298 gnd.n890 240.244
R5738 gnd.n6298 gnd.n892 240.244
R5739 gnd.n6294 gnd.n892 240.244
R5740 gnd.n6294 gnd.n898 240.244
R5741 gnd.n6290 gnd.n898 240.244
R5742 gnd.n6290 gnd.n900 240.244
R5743 gnd.n6286 gnd.n900 240.244
R5744 gnd.n6286 gnd.n906 240.244
R5745 gnd.n6282 gnd.n906 240.244
R5746 gnd.n6282 gnd.n908 240.244
R5747 gnd.n6278 gnd.n908 240.244
R5748 gnd.n6278 gnd.n914 240.244
R5749 gnd.n6274 gnd.n914 240.244
R5750 gnd.n6274 gnd.n916 240.244
R5751 gnd.n6270 gnd.n916 240.244
R5752 gnd.n6270 gnd.n922 240.244
R5753 gnd.n6266 gnd.n922 240.244
R5754 gnd.n6266 gnd.n924 240.244
R5755 gnd.n6262 gnd.n924 240.244
R5756 gnd.n6262 gnd.n930 240.244
R5757 gnd.n6258 gnd.n930 240.244
R5758 gnd.n6258 gnd.n932 240.244
R5759 gnd.n6254 gnd.n932 240.244
R5760 gnd.n6254 gnd.n938 240.244
R5761 gnd.n6250 gnd.n938 240.244
R5762 gnd.n6250 gnd.n940 240.244
R5763 gnd.n6246 gnd.n940 240.244
R5764 gnd.n6246 gnd.n946 240.244
R5765 gnd.n6242 gnd.n946 240.244
R5766 gnd.n6242 gnd.n948 240.244
R5767 gnd.n6238 gnd.n948 240.244
R5768 gnd.n6238 gnd.n954 240.244
R5769 gnd.n6234 gnd.n954 240.244
R5770 gnd.n6234 gnd.n956 240.244
R5771 gnd.n6230 gnd.n956 240.244
R5772 gnd.n6230 gnd.n962 240.244
R5773 gnd.n6226 gnd.n962 240.244
R5774 gnd.n6226 gnd.n964 240.244
R5775 gnd.n6222 gnd.n964 240.244
R5776 gnd.n6222 gnd.n970 240.244
R5777 gnd.n6218 gnd.n970 240.244
R5778 gnd.n6218 gnd.n972 240.244
R5779 gnd.n6214 gnd.n972 240.244
R5780 gnd.n6214 gnd.n978 240.244
R5781 gnd.n6210 gnd.n978 240.244
R5782 gnd.n6210 gnd.n980 240.244
R5783 gnd.n6206 gnd.n980 240.244
R5784 gnd.n6206 gnd.n986 240.244
R5785 gnd.n6202 gnd.n986 240.244
R5786 gnd.n6202 gnd.n988 240.244
R5787 gnd.n6198 gnd.n988 240.244
R5788 gnd.n6198 gnd.n994 240.244
R5789 gnd.n6194 gnd.n994 240.244
R5790 gnd.n6194 gnd.n996 240.244
R5791 gnd.n6190 gnd.n996 240.244
R5792 gnd.n6190 gnd.n1002 240.244
R5793 gnd.n6186 gnd.n1002 240.244
R5794 gnd.n6186 gnd.n1004 240.244
R5795 gnd.n6182 gnd.n1004 240.244
R5796 gnd.n6182 gnd.n1010 240.244
R5797 gnd.n6178 gnd.n1010 240.244
R5798 gnd.n6178 gnd.n1012 240.244
R5799 gnd.n6174 gnd.n1012 240.244
R5800 gnd.n6174 gnd.n1018 240.244
R5801 gnd.n6170 gnd.n1018 240.244
R5802 gnd.n6170 gnd.n1020 240.244
R5803 gnd.n6166 gnd.n1020 240.244
R5804 gnd.n6166 gnd.n1026 240.244
R5805 gnd.n6162 gnd.n1026 240.244
R5806 gnd.n6162 gnd.n1028 240.244
R5807 gnd.n6158 gnd.n1028 240.244
R5808 gnd.n6158 gnd.n1034 240.244
R5809 gnd.n6154 gnd.n1034 240.244
R5810 gnd.n6154 gnd.n1036 240.244
R5811 gnd.n6150 gnd.n1036 240.244
R5812 gnd.n6150 gnd.n1042 240.244
R5813 gnd.n6146 gnd.n1042 240.244
R5814 gnd.n6146 gnd.n1044 240.244
R5815 gnd.n6142 gnd.n1044 240.244
R5816 gnd.n4756 gnd.n2260 240.244
R5817 gnd.n4762 gnd.n2260 240.244
R5818 gnd.n4763 gnd.n4762 240.244
R5819 gnd.n4764 gnd.n4763 240.244
R5820 gnd.n4764 gnd.n1279 240.244
R5821 gnd.n4770 gnd.n1279 240.244
R5822 gnd.n4770 gnd.n1291 240.244
R5823 gnd.n4789 gnd.n1291 240.244
R5824 gnd.n4789 gnd.n2251 240.244
R5825 gnd.n2251 gnd.n1379 240.244
R5826 gnd.n4824 gnd.n1379 240.244
R5827 gnd.n4824 gnd.n1393 240.244
R5828 gnd.n2244 gnd.n1393 240.244
R5829 gnd.n4836 gnd.n2244 240.244
R5830 gnd.n4836 gnd.n2242 240.244
R5831 gnd.n2242 gnd.n2238 240.244
R5832 gnd.n2238 gnd.n2229 240.244
R5833 gnd.n2229 gnd.n2220 240.244
R5834 gnd.n4888 gnd.n2220 240.244
R5835 gnd.n4888 gnd.n2221 240.244
R5836 gnd.n2221 gnd.n2190 240.244
R5837 gnd.n4895 gnd.n2190 240.244
R5838 gnd.n4896 gnd.n4895 240.244
R5839 gnd.n4896 gnd.n2212 240.244
R5840 gnd.n4929 gnd.n2212 240.244
R5841 gnd.n4929 gnd.n2213 240.244
R5842 gnd.n4901 gnd.n2213 240.244
R5843 gnd.n4902 gnd.n4901 240.244
R5844 gnd.n4902 gnd.n2164 240.244
R5845 gnd.n2164 gnd.n2156 240.244
R5846 gnd.n4906 gnd.n2156 240.244
R5847 gnd.n4906 gnd.n2149 240.244
R5848 gnd.n4907 gnd.n2149 240.244
R5849 gnd.n4910 gnd.n4907 240.244
R5850 gnd.n4910 gnd.n2131 240.244
R5851 gnd.n2131 gnd.n2120 240.244
R5852 gnd.n5061 gnd.n2120 240.244
R5853 gnd.n5061 gnd.n2115 240.244
R5854 gnd.n5088 gnd.n2115 240.244
R5855 gnd.n5088 gnd.n2109 240.244
R5856 gnd.n5066 gnd.n2109 240.244
R5857 gnd.n5066 gnd.n2101 240.244
R5858 gnd.n5067 gnd.n2101 240.244
R5859 gnd.n5067 gnd.n2085 240.244
R5860 gnd.n5070 gnd.n2085 240.244
R5861 gnd.n5070 gnd.n2078 240.244
R5862 gnd.n5071 gnd.n2078 240.244
R5863 gnd.n5071 gnd.n2066 240.244
R5864 gnd.n2066 gnd.n2056 240.244
R5865 gnd.n5186 gnd.n2056 240.244
R5866 gnd.n5186 gnd.n2051 240.244
R5867 gnd.n5196 gnd.n2051 240.244
R5868 gnd.n5196 gnd.n2041 240.244
R5869 gnd.n2041 gnd.n2029 240.244
R5870 gnd.n5222 gnd.n2029 240.244
R5871 gnd.n5223 gnd.n5222 240.244
R5872 gnd.n5224 gnd.n5223 240.244
R5873 gnd.n5224 gnd.n2012 240.244
R5874 gnd.n5259 gnd.n2012 240.244
R5875 gnd.n5259 gnd.n2004 240.244
R5876 gnd.n2004 gnd.n2000 240.244
R5877 gnd.n2000 gnd.n1993 240.244
R5878 gnd.n5229 gnd.n1993 240.244
R5879 gnd.n5229 gnd.n1986 240.244
R5880 gnd.n5232 gnd.n1986 240.244
R5881 gnd.n5233 gnd.n5232 240.244
R5882 gnd.n5233 gnd.n1968 240.244
R5883 gnd.n5235 gnd.n1968 240.244
R5884 gnd.n5235 gnd.n1959 240.244
R5885 gnd.n5238 gnd.n1959 240.244
R5886 gnd.n5238 gnd.n1940 240.244
R5887 gnd.n1940 gnd.n1930 240.244
R5888 gnd.n5388 gnd.n1930 240.244
R5889 gnd.n5388 gnd.n1925 240.244
R5890 gnd.n5395 gnd.n1925 240.244
R5891 gnd.n5395 gnd.n1791 240.244
R5892 gnd.n1791 gnd.n1783 240.244
R5893 gnd.n5497 gnd.n1783 240.244
R5894 gnd.n5497 gnd.n1779 240.244
R5895 gnd.n5503 gnd.n1779 240.244
R5896 gnd.n5503 gnd.n1491 240.244
R5897 gnd.n5822 gnd.n1491 240.244
R5898 gnd.n4450 gnd.n4449 240.244
R5899 gnd.n4445 gnd.n4444 240.244
R5900 gnd.n4458 gnd.n4457 240.244
R5901 gnd.n4460 gnd.n4459 240.244
R5902 gnd.n4467 gnd.n4466 240.244
R5903 gnd.n4469 gnd.n4468 240.244
R5904 gnd.n4479 gnd.n4478 240.244
R5905 gnd.n4487 gnd.n4486 240.244
R5906 gnd.n4489 gnd.n4488 240.244
R5907 gnd.n4499 gnd.n4498 240.244
R5908 gnd.n4507 gnd.n4506 240.244
R5909 gnd.n4509 gnd.n4508 240.244
R5910 gnd.n4521 gnd.n4520 240.244
R5911 gnd.n4737 gnd.n2288 240.244
R5912 gnd.n4722 gnd.n2266 240.244
R5913 gnd.n4723 gnd.n4722 240.244
R5914 gnd.n4725 gnd.n4723 240.244
R5915 gnd.n4726 gnd.n4725 240.244
R5916 gnd.n4726 gnd.n1281 240.244
R5917 gnd.n4778 gnd.n1281 240.244
R5918 gnd.n4778 gnd.n1293 240.244
R5919 gnd.n4787 gnd.n1293 240.244
R5920 gnd.n4787 gnd.n2252 240.244
R5921 gnd.n2252 gnd.n1381 240.244
R5922 gnd.n1395 gnd.n1381 240.244
R5923 gnd.n5932 gnd.n1395 240.244
R5924 gnd.n5932 gnd.n1396 240.244
R5925 gnd.n1401 gnd.n1396 240.244
R5926 gnd.n1402 gnd.n1401 240.244
R5927 gnd.n1403 gnd.n1402 240.244
R5928 gnd.n4878 gnd.n1403 240.244
R5929 gnd.n4878 gnd.n1406 240.244
R5930 gnd.n1407 gnd.n1406 240.244
R5931 gnd.n1408 gnd.n1407 240.244
R5932 gnd.n2192 gnd.n1408 240.244
R5933 gnd.n2192 gnd.n1411 240.244
R5934 gnd.n1412 gnd.n1411 240.244
R5935 gnd.n1413 gnd.n1412 240.244
R5936 gnd.n4931 gnd.n1413 240.244
R5937 gnd.n4931 gnd.n1416 240.244
R5938 gnd.n1417 gnd.n1416 240.244
R5939 gnd.n1418 gnd.n1417 240.244
R5940 gnd.n4985 gnd.n1418 240.244
R5941 gnd.n4985 gnd.n1421 240.244
R5942 gnd.n1422 gnd.n1421 240.244
R5943 gnd.n1423 gnd.n1422 240.244
R5944 gnd.n2143 gnd.n1423 240.244
R5945 gnd.n2143 gnd.n1426 240.244
R5946 gnd.n1427 gnd.n1426 240.244
R5947 gnd.n1428 gnd.n1427 240.244
R5948 gnd.n2123 gnd.n1428 240.244
R5949 gnd.n2123 gnd.n1431 240.244
R5950 gnd.n1432 gnd.n1431 240.244
R5951 gnd.n1433 gnd.n1432 240.244
R5952 gnd.n2098 gnd.n1433 240.244
R5953 gnd.n2098 gnd.n1436 240.244
R5954 gnd.n1437 gnd.n1436 240.244
R5955 gnd.n1438 gnd.n1437 240.244
R5956 gnd.n2087 gnd.n1438 240.244
R5957 gnd.n2087 gnd.n1441 240.244
R5958 gnd.n1442 gnd.n1441 240.244
R5959 gnd.n1443 gnd.n1442 240.244
R5960 gnd.n2068 gnd.n1443 240.244
R5961 gnd.n2068 gnd.n1446 240.244
R5962 gnd.n1447 gnd.n1446 240.244
R5963 gnd.n1448 gnd.n1447 240.244
R5964 gnd.n5210 gnd.n1448 240.244
R5965 gnd.n5210 gnd.n1451 240.244
R5966 gnd.n1452 gnd.n1451 240.244
R5967 gnd.n1453 gnd.n1452 240.244
R5968 gnd.n2018 gnd.n1453 240.244
R5969 gnd.n2018 gnd.n1456 240.244
R5970 gnd.n1457 gnd.n1456 240.244
R5971 gnd.n1458 gnd.n1457 240.244
R5972 gnd.n5295 gnd.n1458 240.244
R5973 gnd.n5295 gnd.n1461 240.244
R5974 gnd.n1462 gnd.n1461 240.244
R5975 gnd.n1463 gnd.n1462 240.244
R5976 gnd.n1980 gnd.n1463 240.244
R5977 gnd.n1980 gnd.n1466 240.244
R5978 gnd.n1467 gnd.n1466 240.244
R5979 gnd.n1468 gnd.n1467 240.244
R5980 gnd.n1961 gnd.n1468 240.244
R5981 gnd.n1961 gnd.n1471 240.244
R5982 gnd.n1472 gnd.n1471 240.244
R5983 gnd.n1473 gnd.n1472 240.244
R5984 gnd.n1932 gnd.n1473 240.244
R5985 gnd.n1932 gnd.n1476 240.244
R5986 gnd.n1477 gnd.n1476 240.244
R5987 gnd.n1478 gnd.n1477 240.244
R5988 gnd.n5402 gnd.n1478 240.244
R5989 gnd.n5402 gnd.n1481 240.244
R5990 gnd.n1482 gnd.n1481 240.244
R5991 gnd.n1483 gnd.n1482 240.244
R5992 gnd.n1486 gnd.n1483 240.244
R5993 gnd.n5824 gnd.n1486 240.244
R5994 gnd.n1497 gnd.n1496 240.244
R5995 gnd.n1751 gnd.n1500 240.244
R5996 gnd.n1502 gnd.n1501 240.244
R5997 gnd.n1754 gnd.n1506 240.244
R5998 gnd.n1757 gnd.n1507 240.244
R5999 gnd.n1516 gnd.n1515 240.244
R6000 gnd.n1759 gnd.n1523 240.244
R6001 gnd.n1762 gnd.n1524 240.244
R6002 gnd.n1532 gnd.n1531 240.244
R6003 gnd.n1764 gnd.n1539 240.244
R6004 gnd.n1767 gnd.n1540 240.244
R6005 gnd.n1548 gnd.n1547 240.244
R6006 gnd.n1770 gnd.n1749 240.244
R6007 gnd.n5530 gnd.n1487 240.244
R6008 gnd.n1260 gnd.n1259 240.132
R6009 gnd.n1828 gnd.n1827 240.132
R6010 gnd.n6317 gnd.n878 225.874
R6011 gnd.n6318 gnd.n6317 225.874
R6012 gnd.n6319 gnd.n6318 225.874
R6013 gnd.n6319 gnd.n872 225.874
R6014 gnd.n6327 gnd.n872 225.874
R6015 gnd.n6328 gnd.n6327 225.874
R6016 gnd.n6329 gnd.n6328 225.874
R6017 gnd.n6329 gnd.n866 225.874
R6018 gnd.n6337 gnd.n866 225.874
R6019 gnd.n6338 gnd.n6337 225.874
R6020 gnd.n6339 gnd.n6338 225.874
R6021 gnd.n6339 gnd.n860 225.874
R6022 gnd.n6347 gnd.n860 225.874
R6023 gnd.n6348 gnd.n6347 225.874
R6024 gnd.n6349 gnd.n6348 225.874
R6025 gnd.n6349 gnd.n854 225.874
R6026 gnd.n6357 gnd.n854 225.874
R6027 gnd.n6358 gnd.n6357 225.874
R6028 gnd.n6359 gnd.n6358 225.874
R6029 gnd.n6359 gnd.n848 225.874
R6030 gnd.n6367 gnd.n848 225.874
R6031 gnd.n6368 gnd.n6367 225.874
R6032 gnd.n6369 gnd.n6368 225.874
R6033 gnd.n6369 gnd.n842 225.874
R6034 gnd.n6377 gnd.n842 225.874
R6035 gnd.n6378 gnd.n6377 225.874
R6036 gnd.n6379 gnd.n6378 225.874
R6037 gnd.n6379 gnd.n836 225.874
R6038 gnd.n6387 gnd.n836 225.874
R6039 gnd.n6388 gnd.n6387 225.874
R6040 gnd.n6389 gnd.n6388 225.874
R6041 gnd.n6389 gnd.n830 225.874
R6042 gnd.n6397 gnd.n830 225.874
R6043 gnd.n6398 gnd.n6397 225.874
R6044 gnd.n6399 gnd.n6398 225.874
R6045 gnd.n6399 gnd.n824 225.874
R6046 gnd.n6407 gnd.n824 225.874
R6047 gnd.n6408 gnd.n6407 225.874
R6048 gnd.n6409 gnd.n6408 225.874
R6049 gnd.n6409 gnd.n818 225.874
R6050 gnd.n6417 gnd.n818 225.874
R6051 gnd.n6418 gnd.n6417 225.874
R6052 gnd.n6419 gnd.n6418 225.874
R6053 gnd.n6419 gnd.n812 225.874
R6054 gnd.n6427 gnd.n812 225.874
R6055 gnd.n6428 gnd.n6427 225.874
R6056 gnd.n6429 gnd.n6428 225.874
R6057 gnd.n6429 gnd.n806 225.874
R6058 gnd.n6437 gnd.n806 225.874
R6059 gnd.n6438 gnd.n6437 225.874
R6060 gnd.n6439 gnd.n6438 225.874
R6061 gnd.n6439 gnd.n800 225.874
R6062 gnd.n6447 gnd.n800 225.874
R6063 gnd.n6448 gnd.n6447 225.874
R6064 gnd.n6449 gnd.n6448 225.874
R6065 gnd.n6449 gnd.n794 225.874
R6066 gnd.n6457 gnd.n794 225.874
R6067 gnd.n6458 gnd.n6457 225.874
R6068 gnd.n6459 gnd.n6458 225.874
R6069 gnd.n6459 gnd.n788 225.874
R6070 gnd.n6467 gnd.n788 225.874
R6071 gnd.n6468 gnd.n6467 225.874
R6072 gnd.n6469 gnd.n6468 225.874
R6073 gnd.n6469 gnd.n782 225.874
R6074 gnd.n6477 gnd.n782 225.874
R6075 gnd.n6478 gnd.n6477 225.874
R6076 gnd.n6479 gnd.n6478 225.874
R6077 gnd.n6479 gnd.n776 225.874
R6078 gnd.n6487 gnd.n776 225.874
R6079 gnd.n6488 gnd.n6487 225.874
R6080 gnd.n6489 gnd.n6488 225.874
R6081 gnd.n6489 gnd.n770 225.874
R6082 gnd.n6497 gnd.n770 225.874
R6083 gnd.n6498 gnd.n6497 225.874
R6084 gnd.n6499 gnd.n6498 225.874
R6085 gnd.n6499 gnd.n764 225.874
R6086 gnd.n6507 gnd.n764 225.874
R6087 gnd.n6508 gnd.n6507 225.874
R6088 gnd.n6509 gnd.n6508 225.874
R6089 gnd.n6509 gnd.n758 225.874
R6090 gnd.n6517 gnd.n758 225.874
R6091 gnd.n6518 gnd.n6517 225.874
R6092 gnd.n6519 gnd.n6518 225.874
R6093 gnd.n6519 gnd.n752 225.874
R6094 gnd.n6527 gnd.n752 225.874
R6095 gnd.n6528 gnd.n6527 225.874
R6096 gnd.n6529 gnd.n6528 225.874
R6097 gnd.n6529 gnd.n746 225.874
R6098 gnd.n6537 gnd.n746 225.874
R6099 gnd.n6538 gnd.n6537 225.874
R6100 gnd.n6539 gnd.n6538 225.874
R6101 gnd.n6539 gnd.n740 225.874
R6102 gnd.n6547 gnd.n740 225.874
R6103 gnd.n6548 gnd.n6547 225.874
R6104 gnd.n6549 gnd.n6548 225.874
R6105 gnd.n6549 gnd.n734 225.874
R6106 gnd.n6557 gnd.n734 225.874
R6107 gnd.n6558 gnd.n6557 225.874
R6108 gnd.n6559 gnd.n6558 225.874
R6109 gnd.n6559 gnd.n728 225.874
R6110 gnd.n6567 gnd.n728 225.874
R6111 gnd.n6568 gnd.n6567 225.874
R6112 gnd.n6569 gnd.n6568 225.874
R6113 gnd.n6569 gnd.n722 225.874
R6114 gnd.n6577 gnd.n722 225.874
R6115 gnd.n6578 gnd.n6577 225.874
R6116 gnd.n6579 gnd.n6578 225.874
R6117 gnd.n6579 gnd.n716 225.874
R6118 gnd.n6587 gnd.n716 225.874
R6119 gnd.n6588 gnd.n6587 225.874
R6120 gnd.n6589 gnd.n6588 225.874
R6121 gnd.n6589 gnd.n710 225.874
R6122 gnd.n6597 gnd.n710 225.874
R6123 gnd.n6598 gnd.n6597 225.874
R6124 gnd.n6599 gnd.n6598 225.874
R6125 gnd.n6599 gnd.n704 225.874
R6126 gnd.n6607 gnd.n704 225.874
R6127 gnd.n6608 gnd.n6607 225.874
R6128 gnd.n6609 gnd.n6608 225.874
R6129 gnd.n6609 gnd.n698 225.874
R6130 gnd.n6617 gnd.n698 225.874
R6131 gnd.n6618 gnd.n6617 225.874
R6132 gnd.n6619 gnd.n6618 225.874
R6133 gnd.n6619 gnd.n692 225.874
R6134 gnd.n6628 gnd.n692 225.874
R6135 gnd.n6629 gnd.n6628 225.874
R6136 gnd.n6630 gnd.n6629 225.874
R6137 gnd.n6630 gnd.n687 225.874
R6138 gnd.n2998 gnd.t183 224.174
R6139 gnd.n2508 gnd.t172 224.174
R6140 gnd.n1632 gnd.n1569 199.319
R6141 gnd.n1632 gnd.n1570 199.319
R6142 gnd.n1212 gnd.n1172 199.319
R6143 gnd.n1212 gnd.n1171 199.319
R6144 gnd.n1261 gnd.n1258 186.49
R6145 gnd.n1829 gnd.n1826 186.49
R6146 gnd.n3774 gnd.n3773 185
R6147 gnd.n3772 gnd.n3771 185
R6148 gnd.n3751 gnd.n3750 185
R6149 gnd.n3766 gnd.n3765 185
R6150 gnd.n3764 gnd.n3763 185
R6151 gnd.n3755 gnd.n3754 185
R6152 gnd.n3758 gnd.n3757 185
R6153 gnd.n3742 gnd.n3741 185
R6154 gnd.n3740 gnd.n3739 185
R6155 gnd.n3719 gnd.n3718 185
R6156 gnd.n3734 gnd.n3733 185
R6157 gnd.n3732 gnd.n3731 185
R6158 gnd.n3723 gnd.n3722 185
R6159 gnd.n3726 gnd.n3725 185
R6160 gnd.n3710 gnd.n3709 185
R6161 gnd.n3708 gnd.n3707 185
R6162 gnd.n3687 gnd.n3686 185
R6163 gnd.n3702 gnd.n3701 185
R6164 gnd.n3700 gnd.n3699 185
R6165 gnd.n3691 gnd.n3690 185
R6166 gnd.n3694 gnd.n3693 185
R6167 gnd.n3679 gnd.n3678 185
R6168 gnd.n3677 gnd.n3676 185
R6169 gnd.n3656 gnd.n3655 185
R6170 gnd.n3671 gnd.n3670 185
R6171 gnd.n3669 gnd.n3668 185
R6172 gnd.n3660 gnd.n3659 185
R6173 gnd.n3663 gnd.n3662 185
R6174 gnd.n3647 gnd.n3646 185
R6175 gnd.n3645 gnd.n3644 185
R6176 gnd.n3624 gnd.n3623 185
R6177 gnd.n3639 gnd.n3638 185
R6178 gnd.n3637 gnd.n3636 185
R6179 gnd.n3628 gnd.n3627 185
R6180 gnd.n3631 gnd.n3630 185
R6181 gnd.n3615 gnd.n3614 185
R6182 gnd.n3613 gnd.n3612 185
R6183 gnd.n3592 gnd.n3591 185
R6184 gnd.n3607 gnd.n3606 185
R6185 gnd.n3605 gnd.n3604 185
R6186 gnd.n3596 gnd.n3595 185
R6187 gnd.n3599 gnd.n3598 185
R6188 gnd.n3583 gnd.n3582 185
R6189 gnd.n3581 gnd.n3580 185
R6190 gnd.n3560 gnd.n3559 185
R6191 gnd.n3575 gnd.n3574 185
R6192 gnd.n3573 gnd.n3572 185
R6193 gnd.n3564 gnd.n3563 185
R6194 gnd.n3567 gnd.n3566 185
R6195 gnd.n3552 gnd.n3551 185
R6196 gnd.n3550 gnd.n3549 185
R6197 gnd.n3529 gnd.n3528 185
R6198 gnd.n3544 gnd.n3543 185
R6199 gnd.n3542 gnd.n3541 185
R6200 gnd.n3533 gnd.n3532 185
R6201 gnd.n3536 gnd.n3535 185
R6202 gnd.n2999 gnd.t182 178.987
R6203 gnd.n2509 gnd.t173 178.987
R6204 gnd.n1 gnd.t320 170.774
R6205 gnd.n7 gnd.t23 170.103
R6206 gnd.n6 gnd.t322 170.103
R6207 gnd.n5 gnd.t313 170.103
R6208 gnd.n4 gnd.t35 170.103
R6209 gnd.n3 gnd.t39 170.103
R6210 gnd.n2 gnd.t325 170.103
R6211 gnd.n1 gnd.t3 170.103
R6212 gnd.n1840 gnd.n1839 163.367
R6213 gnd.n1844 gnd.n1843 163.367
R6214 gnd.n1848 gnd.n1847 163.367
R6215 gnd.n1852 gnd.n1851 163.367
R6216 gnd.n1856 gnd.n1855 163.367
R6217 gnd.n1860 gnd.n1859 163.367
R6218 gnd.n1864 gnd.n1863 163.367
R6219 gnd.n1868 gnd.n1867 163.367
R6220 gnd.n1872 gnd.n1871 163.367
R6221 gnd.n1876 gnd.n1875 163.367
R6222 gnd.n1880 gnd.n1879 163.367
R6223 gnd.n1884 gnd.n1883 163.367
R6224 gnd.n1888 gnd.n1887 163.367
R6225 gnd.n1892 gnd.n1891 163.367
R6226 gnd.n1897 gnd.n1896 163.367
R6227 gnd.n1901 gnd.n1900 163.367
R6228 gnd.n5474 gnd.n5473 163.367
R6229 gnd.n5470 gnd.n5469 163.367
R6230 gnd.n5465 gnd.n5464 163.367
R6231 gnd.n5461 gnd.n5460 163.367
R6232 gnd.n5457 gnd.n5456 163.367
R6233 gnd.n5453 gnd.n5452 163.367
R6234 gnd.n5449 gnd.n5448 163.367
R6235 gnd.n5445 gnd.n5444 163.367
R6236 gnd.n5441 gnd.n5440 163.367
R6237 gnd.n5437 gnd.n5436 163.367
R6238 gnd.n5433 gnd.n5432 163.367
R6239 gnd.n5429 gnd.n5428 163.367
R6240 gnd.n5425 gnd.n5424 163.367
R6241 gnd.n5421 gnd.n5420 163.367
R6242 gnd.n5417 gnd.n5416 163.367
R6243 gnd.n5413 gnd.n5412 163.367
R6244 gnd.n1362 gnd.n1277 163.367
R6245 gnd.n1278 gnd.n1277 163.367
R6246 gnd.n1366 gnd.n1278 163.367
R6247 gnd.n1366 gnd.n1294 163.367
R6248 gnd.n5951 gnd.n1294 163.367
R6249 gnd.n5951 gnd.n1295 163.367
R6250 gnd.n5947 gnd.n1295 163.367
R6251 gnd.n5947 gnd.n1370 163.367
R6252 gnd.n1378 gnd.n1370 163.367
R6253 gnd.n4806 gnd.n1378 163.367
R6254 gnd.n4806 gnd.n4795 163.367
R6255 gnd.n4809 gnd.n4795 163.367
R6256 gnd.n4809 gnd.n4803 163.367
R6257 gnd.n4814 gnd.n4803 163.367
R6258 gnd.n4814 gnd.n4804 163.367
R6259 gnd.n4804 gnd.n2240 163.367
R6260 gnd.n4847 gnd.n2240 163.367
R6261 gnd.n4847 gnd.n2237 163.367
R6262 gnd.n4863 gnd.n2237 163.367
R6263 gnd.n4863 gnd.n2230 163.367
R6264 gnd.n4859 gnd.n2230 163.367
R6265 gnd.n4859 gnd.n4858 163.367
R6266 gnd.n4858 gnd.n4857 163.367
R6267 gnd.n4857 gnd.n4853 163.367
R6268 gnd.n4853 gnd.n2189 163.367
R6269 gnd.n2189 gnd.n2183 163.367
R6270 gnd.n4948 gnd.n2183 163.367
R6271 gnd.n4948 gnd.n2181 163.367
R6272 gnd.n4952 gnd.n2181 163.367
R6273 gnd.n4952 gnd.n2175 163.367
R6274 gnd.n4960 gnd.n2175 163.367
R6275 gnd.n4960 gnd.n2173 163.367
R6276 gnd.n4965 gnd.n2173 163.367
R6277 gnd.n4965 gnd.n2166 163.367
R6278 gnd.n4974 gnd.n2166 163.367
R6279 gnd.n4975 gnd.n4974 163.367
R6280 gnd.n4975 gnd.n2163 163.367
R6281 gnd.n4983 gnd.n2163 163.367
R6282 gnd.n4983 gnd.n2157 163.367
R6283 gnd.n4979 gnd.n2157 163.367
R6284 gnd.n4979 gnd.n2148 163.367
R6285 gnd.n2148 gnd.n2141 163.367
R6286 gnd.n5012 gnd.n2141 163.367
R6287 gnd.n5012 gnd.n2138 163.367
R6288 gnd.n5037 gnd.n2138 163.367
R6289 gnd.n5037 gnd.n2139 163.367
R6290 gnd.n2139 gnd.n2132 163.367
R6291 gnd.n5032 gnd.n2132 163.367
R6292 gnd.n5032 gnd.n5030 163.367
R6293 gnd.n5030 gnd.n5029 163.367
R6294 gnd.n5029 gnd.n5018 163.367
R6295 gnd.n5018 gnd.n2114 163.367
R6296 gnd.n5024 gnd.n2114 163.367
R6297 gnd.n5024 gnd.n2110 163.367
R6298 gnd.n5021 gnd.n2110 163.367
R6299 gnd.n5021 gnd.n2100 163.367
R6300 gnd.n2100 gnd.n2093 163.367
R6301 gnd.n5113 gnd.n2093 163.367
R6302 gnd.n5114 gnd.n5113 163.367
R6303 gnd.n5114 gnd.n2086 163.367
R6304 gnd.n5118 gnd.n2086 163.367
R6305 gnd.n5118 gnd.n2077 163.367
R6306 gnd.n5137 gnd.n2077 163.367
R6307 gnd.n5137 gnd.n2075 163.367
R6308 gnd.n5161 gnd.n2075 163.367
R6309 gnd.n5161 gnd.n2067 163.367
R6310 gnd.n5157 gnd.n2067 163.367
R6311 gnd.n5157 gnd.n5155 163.367
R6312 gnd.n5155 gnd.n5154 163.367
R6313 gnd.n5154 gnd.n5141 163.367
R6314 gnd.n5141 gnd.n2050 163.367
R6315 gnd.n5149 gnd.n2050 163.367
R6316 gnd.n5149 gnd.n2042 163.367
R6317 gnd.n5146 gnd.n2042 163.367
R6318 gnd.n5146 gnd.n5145 163.367
R6319 gnd.n5145 gnd.n5144 163.367
R6320 gnd.n5144 gnd.n2016 163.367
R6321 gnd.n5269 gnd.n2016 163.367
R6322 gnd.n5269 gnd.n2013 163.367
R6323 gnd.n5274 gnd.n2013 163.367
R6324 gnd.n5274 gnd.n2014 163.367
R6325 gnd.n2014 gnd.n2002 163.367
R6326 gnd.n5285 gnd.n2002 163.367
R6327 gnd.n5285 gnd.n1999 163.367
R6328 gnd.n5293 gnd.n1999 163.367
R6329 gnd.n5293 gnd.n1994 163.367
R6330 gnd.n5289 gnd.n1994 163.367
R6331 gnd.n5289 gnd.n1985 163.367
R6332 gnd.n1985 gnd.n1977 163.367
R6333 gnd.n5322 gnd.n1977 163.367
R6334 gnd.n5322 gnd.n1974 163.367
R6335 gnd.n5332 gnd.n1974 163.367
R6336 gnd.n5332 gnd.n1975 163.367
R6337 gnd.n1975 gnd.n1969 163.367
R6338 gnd.n5327 gnd.n1969 163.367
R6339 gnd.n5327 gnd.n1958 163.367
R6340 gnd.n1958 gnd.n1952 163.367
R6341 gnd.n5356 gnd.n1952 163.367
R6342 gnd.n5357 gnd.n5356 163.367
R6343 gnd.n5357 gnd.n1941 163.367
R6344 gnd.n5361 gnd.n1941 163.367
R6345 gnd.n5361 gnd.n1950 163.367
R6346 gnd.n5366 gnd.n1950 163.367
R6347 gnd.n5366 gnd.n1923 163.367
R6348 gnd.n5397 gnd.n1923 163.367
R6349 gnd.n5398 gnd.n5397 163.367
R6350 gnd.n5398 gnd.n1792 163.367
R6351 gnd.n5405 gnd.n1792 163.367
R6352 gnd.n5406 gnd.n5405 163.367
R6353 gnd.n5406 gnd.n1798 163.367
R6354 gnd.n1252 gnd.n1251 163.367
R6355 gnd.n6023 gnd.n1251 163.367
R6356 gnd.n6021 gnd.n6020 163.367
R6357 gnd.n6017 gnd.n6016 163.367
R6358 gnd.n6013 gnd.n6012 163.367
R6359 gnd.n6009 gnd.n6008 163.367
R6360 gnd.n6005 gnd.n6004 163.367
R6361 gnd.n6001 gnd.n6000 163.367
R6362 gnd.n5997 gnd.n5996 163.367
R6363 gnd.n5993 gnd.n5992 163.367
R6364 gnd.n5989 gnd.n5988 163.367
R6365 gnd.n5985 gnd.n5984 163.367
R6366 gnd.n5981 gnd.n5980 163.367
R6367 gnd.n5977 gnd.n5976 163.367
R6368 gnd.n5973 gnd.n5972 163.367
R6369 gnd.n5969 gnd.n5968 163.367
R6370 gnd.n6032 gnd.n1217 163.367
R6371 gnd.n1300 gnd.n1299 163.367
R6372 gnd.n1305 gnd.n1304 163.367
R6373 gnd.n1309 gnd.n1308 163.367
R6374 gnd.n1313 gnd.n1312 163.367
R6375 gnd.n1317 gnd.n1316 163.367
R6376 gnd.n1321 gnd.n1320 163.367
R6377 gnd.n1325 gnd.n1324 163.367
R6378 gnd.n1329 gnd.n1328 163.367
R6379 gnd.n1333 gnd.n1332 163.367
R6380 gnd.n1337 gnd.n1336 163.367
R6381 gnd.n1341 gnd.n1340 163.367
R6382 gnd.n1345 gnd.n1344 163.367
R6383 gnd.n1349 gnd.n1348 163.367
R6384 gnd.n1353 gnd.n1352 163.367
R6385 gnd.n1357 gnd.n1356 163.367
R6386 gnd.n5961 gnd.n1253 163.367
R6387 gnd.n5961 gnd.n1275 163.367
R6388 gnd.n4771 gnd.n1275 163.367
R6389 gnd.n4775 gnd.n4771 163.367
R6390 gnd.n4775 gnd.n1290 163.367
R6391 gnd.n1372 gnd.n1290 163.367
R6392 gnd.n5945 gnd.n1372 163.367
R6393 gnd.n5945 gnd.n1373 163.367
R6394 gnd.n5941 gnd.n1373 163.367
R6395 gnd.n5941 gnd.n1376 163.367
R6396 gnd.n4821 gnd.n1376 163.367
R6397 gnd.n4821 gnd.n4796 163.367
R6398 gnd.n4817 gnd.n4796 163.367
R6399 gnd.n4817 gnd.n4816 163.367
R6400 gnd.n4816 gnd.n4801 163.367
R6401 gnd.n4801 gnd.n4798 163.367
R6402 gnd.n4798 gnd.n2236 163.367
R6403 gnd.n4867 gnd.n2236 163.367
R6404 gnd.n4867 gnd.n2233 163.367
R6405 gnd.n4876 gnd.n2233 163.367
R6406 gnd.n4876 gnd.n2234 163.367
R6407 gnd.n4872 gnd.n2234 163.367
R6408 gnd.n4872 gnd.n4871 163.367
R6409 gnd.n4871 gnd.n2188 163.367
R6410 gnd.n4942 gnd.n2188 163.367
R6411 gnd.n4942 gnd.n2186 163.367
R6412 gnd.n4946 gnd.n2186 163.367
R6413 gnd.n4946 gnd.n2179 163.367
R6414 gnd.n4954 gnd.n2179 163.367
R6415 gnd.n4954 gnd.n2177 163.367
R6416 gnd.n4958 gnd.n2177 163.367
R6417 gnd.n4958 gnd.n2171 163.367
R6418 gnd.n4968 gnd.n2171 163.367
R6419 gnd.n4968 gnd.n2169 163.367
R6420 gnd.n4972 gnd.n2169 163.367
R6421 gnd.n4972 gnd.n2161 163.367
R6422 gnd.n4988 gnd.n2161 163.367
R6423 gnd.n4988 gnd.n2159 163.367
R6424 gnd.n4992 gnd.n2159 163.367
R6425 gnd.n4992 gnd.n2147 163.367
R6426 gnd.n5006 gnd.n2147 163.367
R6427 gnd.n5006 gnd.n2145 163.367
R6428 gnd.n5010 gnd.n2145 163.367
R6429 gnd.n5010 gnd.n2137 163.367
R6430 gnd.n5039 gnd.n2137 163.367
R6431 gnd.n5039 gnd.n2134 163.367
R6432 gnd.n5048 gnd.n2134 163.367
R6433 gnd.n5048 gnd.n2135 163.367
R6434 gnd.n5044 gnd.n2135 163.367
R6435 gnd.n5044 gnd.n5043 163.367
R6436 gnd.n5043 gnd.n2113 163.367
R6437 gnd.n5091 gnd.n2113 163.367
R6438 gnd.n5091 gnd.n2111 163.367
R6439 gnd.n5095 gnd.n2111 163.367
R6440 gnd.n5095 gnd.n2097 163.367
R6441 gnd.n5107 gnd.n2097 163.367
R6442 gnd.n5107 gnd.n2095 163.367
R6443 gnd.n5111 gnd.n2095 163.367
R6444 gnd.n5111 gnd.n2089 163.367
R6445 gnd.n5125 gnd.n2089 163.367
R6446 gnd.n5125 gnd.n2090 163.367
R6447 gnd.n5121 gnd.n2090 163.367
R6448 gnd.n5121 gnd.n2073 163.367
R6449 gnd.n5164 gnd.n2073 163.367
R6450 gnd.n5164 gnd.n2070 163.367
R6451 gnd.n5173 gnd.n2070 163.367
R6452 gnd.n5173 gnd.n2071 163.367
R6453 gnd.n5169 gnd.n2071 163.367
R6454 gnd.n5169 gnd.n5168 163.367
R6455 gnd.n5168 gnd.n2048 163.367
R6456 gnd.n5199 gnd.n2048 163.367
R6457 gnd.n5199 gnd.n2045 163.367
R6458 gnd.n5208 gnd.n2045 163.367
R6459 gnd.n5208 gnd.n2046 163.367
R6460 gnd.n5204 gnd.n2046 163.367
R6461 gnd.n5204 gnd.n5203 163.367
R6462 gnd.n5203 gnd.n2020 163.367
R6463 gnd.n5267 gnd.n2020 163.367
R6464 gnd.n5267 gnd.n2021 163.367
R6465 gnd.n2021 gnd.n2011 163.367
R6466 gnd.n5262 gnd.n2011 163.367
R6467 gnd.n5262 gnd.n2024 163.367
R6468 gnd.n2024 gnd.n1998 163.367
R6469 gnd.n5298 gnd.n1998 163.367
R6470 gnd.n5298 gnd.n1996 163.367
R6471 gnd.n5302 gnd.n1996 163.367
R6472 gnd.n5302 gnd.n1984 163.367
R6473 gnd.n5316 gnd.n1984 163.367
R6474 gnd.n5316 gnd.n1982 163.367
R6475 gnd.n5320 gnd.n1982 163.367
R6476 gnd.n5320 gnd.n1972 163.367
R6477 gnd.n5334 gnd.n1972 163.367
R6478 gnd.n5334 gnd.n1970 163.367
R6479 gnd.n5338 gnd.n1970 163.367
R6480 gnd.n5338 gnd.n1956 163.367
R6481 gnd.n5350 gnd.n1956 163.367
R6482 gnd.n5350 gnd.n1954 163.367
R6483 gnd.n5354 gnd.n1954 163.367
R6484 gnd.n5354 gnd.n1943 163.367
R6485 gnd.n5375 gnd.n1943 163.367
R6486 gnd.n5375 gnd.n1944 163.367
R6487 gnd.n5371 gnd.n1944 163.367
R6488 gnd.n5371 gnd.n5370 163.367
R6489 gnd.n5370 gnd.n1949 163.367
R6490 gnd.n1949 gnd.n1924 163.367
R6491 gnd.n1924 gnd.n1793 163.367
R6492 gnd.n5483 gnd.n1793 163.367
R6493 gnd.n5483 gnd.n1794 163.367
R6494 gnd.n5479 gnd.n1794 163.367
R6495 gnd.n5479 gnd.n5478 163.367
R6496 gnd.n1835 gnd.n1834 156.462
R6497 gnd.n3714 gnd.n3682 153.042
R6498 gnd.n3778 gnd.n3777 152.079
R6499 gnd.n3746 gnd.n3745 152.079
R6500 gnd.n3714 gnd.n3713 152.079
R6501 gnd.n1266 gnd.n1265 152
R6502 gnd.n1267 gnd.n1256 152
R6503 gnd.n1269 gnd.n1268 152
R6504 gnd.n1271 gnd.n1254 152
R6505 gnd.n1273 gnd.n1272 152
R6506 gnd.n1833 gnd.n1817 152
R6507 gnd.n1825 gnd.n1818 152
R6508 gnd.n1824 gnd.n1823 152
R6509 gnd.n1822 gnd.n1819 152
R6510 gnd.n1820 gnd.t148 150.546
R6511 gnd.t26 gnd.n3756 147.661
R6512 gnd.t47 gnd.n3724 147.661
R6513 gnd.t49 gnd.n3692 147.661
R6514 gnd.t318 gnd.n3661 147.661
R6515 gnd.t63 gnd.n3629 147.661
R6516 gnd.t37 gnd.n3597 147.661
R6517 gnd.t41 gnd.n3565 147.661
R6518 gnd.t311 gnd.n3534 147.661
R6519 gnd.n1919 gnd.n1902 143.351
R6520 gnd.n1233 gnd.n1216 143.351
R6521 gnd.n6031 gnd.n1216 143.351
R6522 gnd.n1263 gnd.t70 130.484
R6523 gnd.n1272 gnd.t136 126.766
R6524 gnd.n1270 gnd.t67 126.766
R6525 gnd.n1256 gnd.t95 126.766
R6526 gnd.n1264 gnd.t177 126.766
R6527 gnd.n1821 gnd.t119 126.766
R6528 gnd.n1823 gnd.t64 126.766
R6529 gnd.n1832 gnd.t109 126.766
R6530 gnd.n1834 gnd.t85 126.766
R6531 gnd.n6639 gnd.n6638 106.719
R6532 gnd.n6640 gnd.n6639 106.719
R6533 gnd.n6640 gnd.n681 106.719
R6534 gnd.n6648 gnd.n681 106.719
R6535 gnd.n6649 gnd.n6648 106.719
R6536 gnd.n6650 gnd.n6649 106.719
R6537 gnd.n6650 gnd.n675 106.719
R6538 gnd.n6658 gnd.n675 106.719
R6539 gnd.n6659 gnd.n6658 106.719
R6540 gnd.n6660 gnd.n6659 106.719
R6541 gnd.n6660 gnd.n669 106.719
R6542 gnd.n6668 gnd.n669 106.719
R6543 gnd.n6669 gnd.n6668 106.719
R6544 gnd.n6670 gnd.n6669 106.719
R6545 gnd.n6670 gnd.n663 106.719
R6546 gnd.n6678 gnd.n663 106.719
R6547 gnd.n6679 gnd.n6678 106.719
R6548 gnd.n6680 gnd.n6679 106.719
R6549 gnd.n6680 gnd.n657 106.719
R6550 gnd.n6688 gnd.n657 106.719
R6551 gnd.n6689 gnd.n6688 106.719
R6552 gnd.n6690 gnd.n6689 106.719
R6553 gnd.n6690 gnd.n651 106.719
R6554 gnd.n6698 gnd.n651 106.719
R6555 gnd.n6699 gnd.n6698 106.719
R6556 gnd.n6700 gnd.n6699 106.719
R6557 gnd.n6700 gnd.n645 106.719
R6558 gnd.n6708 gnd.n645 106.719
R6559 gnd.n6709 gnd.n6708 106.719
R6560 gnd.n6710 gnd.n6709 106.719
R6561 gnd.n6710 gnd.n639 106.719
R6562 gnd.n6718 gnd.n639 106.719
R6563 gnd.n6719 gnd.n6718 106.719
R6564 gnd.n6720 gnd.n6719 106.719
R6565 gnd.n6720 gnd.n633 106.719
R6566 gnd.n6728 gnd.n633 106.719
R6567 gnd.n6729 gnd.n6728 106.719
R6568 gnd.n6730 gnd.n6729 106.719
R6569 gnd.n6730 gnd.n627 106.719
R6570 gnd.n6738 gnd.n627 106.719
R6571 gnd.n6739 gnd.n6738 106.719
R6572 gnd.n6740 gnd.n6739 106.719
R6573 gnd.n6740 gnd.n621 106.719
R6574 gnd.n6748 gnd.n621 106.719
R6575 gnd.n6749 gnd.n6748 106.719
R6576 gnd.n6750 gnd.n6749 106.719
R6577 gnd.n6750 gnd.n615 106.719
R6578 gnd.n6758 gnd.n615 106.719
R6579 gnd.n6759 gnd.n6758 106.719
R6580 gnd.n6760 gnd.n6759 106.719
R6581 gnd.n6760 gnd.n609 106.719
R6582 gnd.n6768 gnd.n609 106.719
R6583 gnd.n6769 gnd.n6768 106.719
R6584 gnd.n6770 gnd.n6769 106.719
R6585 gnd.n6770 gnd.n603 106.719
R6586 gnd.n6778 gnd.n603 106.719
R6587 gnd.n6779 gnd.n6778 106.719
R6588 gnd.n6780 gnd.n6779 106.719
R6589 gnd.n6780 gnd.n597 106.719
R6590 gnd.n6788 gnd.n597 106.719
R6591 gnd.n6789 gnd.n6788 106.719
R6592 gnd.n6790 gnd.n6789 106.719
R6593 gnd.n6790 gnd.n591 106.719
R6594 gnd.n6798 gnd.n591 106.719
R6595 gnd.n6799 gnd.n6798 106.719
R6596 gnd.n6800 gnd.n6799 106.719
R6597 gnd.n6800 gnd.n585 106.719
R6598 gnd.n6808 gnd.n585 106.719
R6599 gnd.n6809 gnd.n6808 106.719
R6600 gnd.n6810 gnd.n6809 106.719
R6601 gnd.n6810 gnd.n579 106.719
R6602 gnd.n6818 gnd.n579 106.719
R6603 gnd.n6819 gnd.n6818 106.719
R6604 gnd.n6820 gnd.n6819 106.719
R6605 gnd.n6820 gnd.n573 106.719
R6606 gnd.n6828 gnd.n573 106.719
R6607 gnd.n6829 gnd.n6828 106.719
R6608 gnd.n6830 gnd.n6829 106.719
R6609 gnd.n6830 gnd.n567 106.719
R6610 gnd.n6838 gnd.n567 106.719
R6611 gnd.n6839 gnd.n6838 106.719
R6612 gnd.n6841 gnd.n6839 106.719
R6613 gnd.n6841 gnd.n6840 106.719
R6614 gnd.n3773 gnd.n3772 104.615
R6615 gnd.n3772 gnd.n3750 104.615
R6616 gnd.n3765 gnd.n3750 104.615
R6617 gnd.n3765 gnd.n3764 104.615
R6618 gnd.n3764 gnd.n3754 104.615
R6619 gnd.n3757 gnd.n3754 104.615
R6620 gnd.n3741 gnd.n3740 104.615
R6621 gnd.n3740 gnd.n3718 104.615
R6622 gnd.n3733 gnd.n3718 104.615
R6623 gnd.n3733 gnd.n3732 104.615
R6624 gnd.n3732 gnd.n3722 104.615
R6625 gnd.n3725 gnd.n3722 104.615
R6626 gnd.n3709 gnd.n3708 104.615
R6627 gnd.n3708 gnd.n3686 104.615
R6628 gnd.n3701 gnd.n3686 104.615
R6629 gnd.n3701 gnd.n3700 104.615
R6630 gnd.n3700 gnd.n3690 104.615
R6631 gnd.n3693 gnd.n3690 104.615
R6632 gnd.n3678 gnd.n3677 104.615
R6633 gnd.n3677 gnd.n3655 104.615
R6634 gnd.n3670 gnd.n3655 104.615
R6635 gnd.n3670 gnd.n3669 104.615
R6636 gnd.n3669 gnd.n3659 104.615
R6637 gnd.n3662 gnd.n3659 104.615
R6638 gnd.n3646 gnd.n3645 104.615
R6639 gnd.n3645 gnd.n3623 104.615
R6640 gnd.n3638 gnd.n3623 104.615
R6641 gnd.n3638 gnd.n3637 104.615
R6642 gnd.n3637 gnd.n3627 104.615
R6643 gnd.n3630 gnd.n3627 104.615
R6644 gnd.n3614 gnd.n3613 104.615
R6645 gnd.n3613 gnd.n3591 104.615
R6646 gnd.n3606 gnd.n3591 104.615
R6647 gnd.n3606 gnd.n3605 104.615
R6648 gnd.n3605 gnd.n3595 104.615
R6649 gnd.n3598 gnd.n3595 104.615
R6650 gnd.n3582 gnd.n3581 104.615
R6651 gnd.n3581 gnd.n3559 104.615
R6652 gnd.n3574 gnd.n3559 104.615
R6653 gnd.n3574 gnd.n3573 104.615
R6654 gnd.n3573 gnd.n3563 104.615
R6655 gnd.n3566 gnd.n3563 104.615
R6656 gnd.n3551 gnd.n3550 104.615
R6657 gnd.n3550 gnd.n3528 104.615
R6658 gnd.n3543 gnd.n3528 104.615
R6659 gnd.n3543 gnd.n3542 104.615
R6660 gnd.n3542 gnd.n3532 104.615
R6661 gnd.n3535 gnd.n3532 104.615
R6662 gnd.n2924 gnd.t128 100.632
R6663 gnd.n2482 gnd.t159 100.632
R6664 gnd.n350 gnd.n348 99.6594
R6665 gnd.n356 gnd.n341 99.6594
R6666 gnd.n360 gnd.n358 99.6594
R6667 gnd.n366 gnd.n337 99.6594
R6668 gnd.n370 gnd.n368 99.6594
R6669 gnd.n376 gnd.n333 99.6594
R6670 gnd.n381 gnd.n378 99.6594
R6671 gnd.n379 gnd.n329 99.6594
R6672 gnd.n391 gnd.n389 99.6594
R6673 gnd.n397 gnd.n323 99.6594
R6674 gnd.n401 gnd.n399 99.6594
R6675 gnd.n407 gnd.n319 99.6594
R6676 gnd.n411 gnd.n409 99.6594
R6677 gnd.n417 gnd.n315 99.6594
R6678 gnd.n421 gnd.n419 99.6594
R6679 gnd.n427 gnd.n311 99.6594
R6680 gnd.n431 gnd.n429 99.6594
R6681 gnd.n437 gnd.n307 99.6594
R6682 gnd.n441 gnd.n439 99.6594
R6683 gnd.n447 gnd.n301 99.6594
R6684 gnd.n451 gnd.n449 99.6594
R6685 gnd.n457 gnd.n297 99.6594
R6686 gnd.n461 gnd.n459 99.6594
R6687 gnd.n467 gnd.n293 99.6594
R6688 gnd.n471 gnd.n469 99.6594
R6689 gnd.n477 gnd.n289 99.6594
R6690 gnd.n481 gnd.n479 99.6594
R6691 gnd.n487 gnd.n285 99.6594
R6692 gnd.n490 gnd.n489 99.6594
R6693 gnd.n5754 gnd.n5753 99.6594
R6694 gnd.n5748 gnd.n1558 99.6594
R6695 gnd.n5745 gnd.n1559 99.6594
R6696 gnd.n5741 gnd.n1560 99.6594
R6697 gnd.n5737 gnd.n1561 99.6594
R6698 gnd.n5733 gnd.n1562 99.6594
R6699 gnd.n5729 gnd.n1563 99.6594
R6700 gnd.n5725 gnd.n1564 99.6594
R6701 gnd.n5721 gnd.n1565 99.6594
R6702 gnd.n5716 gnd.n1566 99.6594
R6703 gnd.n5712 gnd.n1567 99.6594
R6704 gnd.n5708 gnd.n1568 99.6594
R6705 gnd.n5704 gnd.n1569 99.6594
R6706 gnd.n5699 gnd.n1571 99.6594
R6707 gnd.n5695 gnd.n1572 99.6594
R6708 gnd.n5691 gnd.n1573 99.6594
R6709 gnd.n5687 gnd.n1574 99.6594
R6710 gnd.n5683 gnd.n1575 99.6594
R6711 gnd.n5679 gnd.n1576 99.6594
R6712 gnd.n5675 gnd.n1577 99.6594
R6713 gnd.n5671 gnd.n1578 99.6594
R6714 gnd.n5667 gnd.n1579 99.6594
R6715 gnd.n5663 gnd.n1580 99.6594
R6716 gnd.n5659 gnd.n1581 99.6594
R6717 gnd.n5655 gnd.n1582 99.6594
R6718 gnd.n5651 gnd.n1583 99.6594
R6719 gnd.n5647 gnd.n1584 99.6594
R6720 gnd.n5643 gnd.n1585 99.6594
R6721 gnd.n6083 gnd.n6082 99.6594
R6722 gnd.n6078 gnd.n1183 99.6594
R6723 gnd.n6074 gnd.n1182 99.6594
R6724 gnd.n6070 gnd.n1181 99.6594
R6725 gnd.n6066 gnd.n1180 99.6594
R6726 gnd.n6062 gnd.n1179 99.6594
R6727 gnd.n6058 gnd.n1178 99.6594
R6728 gnd.n6054 gnd.n1177 99.6594
R6729 gnd.n6049 gnd.n1176 99.6594
R6730 gnd.n6045 gnd.n1175 99.6594
R6731 gnd.n6041 gnd.n1174 99.6594
R6732 gnd.n6037 gnd.n1173 99.6594
R6733 gnd.n4597 gnd.n1171 99.6594
R6734 gnd.n4601 gnd.n1170 99.6594
R6735 gnd.n4607 gnd.n1169 99.6594
R6736 gnd.n4611 gnd.n1168 99.6594
R6737 gnd.n4616 gnd.n1167 99.6594
R6738 gnd.n4620 gnd.n1166 99.6594
R6739 gnd.n4626 gnd.n1165 99.6594
R6740 gnd.n4630 gnd.n1164 99.6594
R6741 gnd.n4636 gnd.n1163 99.6594
R6742 gnd.n4640 gnd.n1162 99.6594
R6743 gnd.n4646 gnd.n1161 99.6594
R6744 gnd.n4650 gnd.n1160 99.6594
R6745 gnd.n4656 gnd.n1159 99.6594
R6746 gnd.n4660 gnd.n1158 99.6594
R6747 gnd.n4665 gnd.n1157 99.6594
R6748 gnd.n4668 gnd.n1156 99.6594
R6749 gnd.n4240 gnd.n4239 99.6594
R6750 gnd.n4234 gnd.n3906 99.6594
R6751 gnd.n4231 gnd.n3907 99.6594
R6752 gnd.n4227 gnd.n3908 99.6594
R6753 gnd.n4223 gnd.n3909 99.6594
R6754 gnd.n4219 gnd.n3910 99.6594
R6755 gnd.n4215 gnd.n3911 99.6594
R6756 gnd.n4211 gnd.n3912 99.6594
R6757 gnd.n4207 gnd.n3913 99.6594
R6758 gnd.n4202 gnd.n3914 99.6594
R6759 gnd.n4198 gnd.n3915 99.6594
R6760 gnd.n4194 gnd.n3916 99.6594
R6761 gnd.n4190 gnd.n3917 99.6594
R6762 gnd.n4186 gnd.n3918 99.6594
R6763 gnd.n4182 gnd.n3919 99.6594
R6764 gnd.n4178 gnd.n3920 99.6594
R6765 gnd.n4174 gnd.n3921 99.6594
R6766 gnd.n4170 gnd.n3922 99.6594
R6767 gnd.n4166 gnd.n3923 99.6594
R6768 gnd.n4162 gnd.n3924 99.6594
R6769 gnd.n4158 gnd.n3925 99.6594
R6770 gnd.n4154 gnd.n3926 99.6594
R6771 gnd.n4150 gnd.n3927 99.6594
R6772 gnd.n4146 gnd.n3928 99.6594
R6773 gnd.n4142 gnd.n3929 99.6594
R6774 gnd.n4138 gnd.n3930 99.6594
R6775 gnd.n4134 gnd.n3931 99.6594
R6776 gnd.n4130 gnd.n3932 99.6594
R6777 gnd.n4242 gnd.n2442 99.6594
R6778 gnd.n3896 gnd.n2465 99.6594
R6779 gnd.n3894 gnd.n2464 99.6594
R6780 gnd.n3890 gnd.n2463 99.6594
R6781 gnd.n3886 gnd.n2462 99.6594
R6782 gnd.n3882 gnd.n2461 99.6594
R6783 gnd.n3878 gnd.n2460 99.6594
R6784 gnd.n3874 gnd.n2459 99.6594
R6785 gnd.n3806 gnd.n2458 99.6594
R6786 gnd.n3136 gnd.n2867 99.6594
R6787 gnd.n2893 gnd.n2874 99.6594
R6788 gnd.n2895 gnd.n2875 99.6594
R6789 gnd.n2903 gnd.n2876 99.6594
R6790 gnd.n2905 gnd.n2877 99.6594
R6791 gnd.n2913 gnd.n2878 99.6594
R6792 gnd.n2915 gnd.n2879 99.6594
R6793 gnd.n2923 gnd.n2880 99.6594
R6794 gnd.n276 gnd.n172 99.6594
R6795 gnd.n274 gnd.n273 99.6594
R6796 gnd.n269 gnd.n179 99.6594
R6797 gnd.n267 gnd.n266 99.6594
R6798 gnd.n262 gnd.n186 99.6594
R6799 gnd.n260 gnd.n259 99.6594
R6800 gnd.n255 gnd.n193 99.6594
R6801 gnd.n253 gnd.n252 99.6594
R6802 gnd.n198 gnd.n197 99.6594
R6803 gnd.n1670 gnd.n1586 99.6594
R6804 gnd.n1588 gnd.n1512 99.6594
R6805 gnd.n1589 gnd.n1519 99.6594
R6806 gnd.n1591 gnd.n1590 99.6594
R6807 gnd.n1593 gnd.n1528 99.6594
R6808 gnd.n1594 gnd.n1535 99.6594
R6809 gnd.n1596 gnd.n1595 99.6594
R6810 gnd.n1598 gnd.n1544 99.6594
R6811 gnd.n5756 gnd.n1553 99.6594
R6812 gnd.n3864 gnd.n2445 99.6594
R6813 gnd.n3860 gnd.n2446 99.6594
R6814 gnd.n3856 gnd.n2447 99.6594
R6815 gnd.n3852 gnd.n2448 99.6594
R6816 gnd.n3848 gnd.n2449 99.6594
R6817 gnd.n3844 gnd.n2450 99.6594
R6818 gnd.n3840 gnd.n2451 99.6594
R6819 gnd.n3836 gnd.n2452 99.6594
R6820 gnd.n3832 gnd.n2453 99.6594
R6821 gnd.n3828 gnd.n2454 99.6594
R6822 gnd.n3824 gnd.n2455 99.6594
R6823 gnd.n3820 gnd.n2456 99.6594
R6824 gnd.n3816 gnd.n2457 99.6594
R6825 gnd.n3051 gnd.n3050 99.6594
R6826 gnd.n3045 gnd.n2962 99.6594
R6827 gnd.n3042 gnd.n2963 99.6594
R6828 gnd.n3038 gnd.n2964 99.6594
R6829 gnd.n3034 gnd.n2965 99.6594
R6830 gnd.n3030 gnd.n2966 99.6594
R6831 gnd.n3026 gnd.n2967 99.6594
R6832 gnd.n3022 gnd.n2968 99.6594
R6833 gnd.n3018 gnd.n2969 99.6594
R6834 gnd.n3014 gnd.n2970 99.6594
R6835 gnd.n3010 gnd.n2971 99.6594
R6836 gnd.n3006 gnd.n2972 99.6594
R6837 gnd.n3053 gnd.n2961 99.6594
R6838 gnd.n4472 gnd.n1146 99.6594
R6839 gnd.n4474 gnd.n1147 99.6594
R6840 gnd.n4482 gnd.n1148 99.6594
R6841 gnd.n4492 gnd.n1149 99.6594
R6842 gnd.n4494 gnd.n1150 99.6594
R6843 gnd.n4502 gnd.n1151 99.6594
R6844 gnd.n4512 gnd.n1152 99.6594
R6845 gnd.n4515 gnd.n1153 99.6594
R6846 gnd.n4716 gnd.n1154 99.6594
R6847 gnd.n4120 gnd.n3933 99.6594
R6848 gnd.n4117 gnd.n3934 99.6594
R6849 gnd.n4113 gnd.n3935 99.6594
R6850 gnd.n4109 gnd.n3936 99.6594
R6851 gnd.n4105 gnd.n3937 99.6594
R6852 gnd.n4101 gnd.n3938 99.6594
R6853 gnd.n4097 gnd.n3939 99.6594
R6854 gnd.n4093 gnd.n3940 99.6594
R6855 gnd.n4089 gnd.n3941 99.6594
R6856 gnd.n4118 gnd.n3933 99.6594
R6857 gnd.n4114 gnd.n3934 99.6594
R6858 gnd.n4110 gnd.n3935 99.6594
R6859 gnd.n4106 gnd.n3936 99.6594
R6860 gnd.n4102 gnd.n3937 99.6594
R6861 gnd.n4098 gnd.n3938 99.6594
R6862 gnd.n4094 gnd.n3939 99.6594
R6863 gnd.n4090 gnd.n3940 99.6594
R6864 gnd.n4023 gnd.n3941 99.6594
R6865 gnd.n4514 gnd.n1154 99.6594
R6866 gnd.n4513 gnd.n1153 99.6594
R6867 gnd.n4503 gnd.n1152 99.6594
R6868 gnd.n4495 gnd.n1151 99.6594
R6869 gnd.n4493 gnd.n1150 99.6594
R6870 gnd.n4483 gnd.n1149 99.6594
R6871 gnd.n4475 gnd.n1148 99.6594
R6872 gnd.n4473 gnd.n1147 99.6594
R6873 gnd.n4463 gnd.n1146 99.6594
R6874 gnd.n3051 gnd.n2974 99.6594
R6875 gnd.n3043 gnd.n2962 99.6594
R6876 gnd.n3039 gnd.n2963 99.6594
R6877 gnd.n3035 gnd.n2964 99.6594
R6878 gnd.n3031 gnd.n2965 99.6594
R6879 gnd.n3027 gnd.n2966 99.6594
R6880 gnd.n3023 gnd.n2967 99.6594
R6881 gnd.n3019 gnd.n2968 99.6594
R6882 gnd.n3015 gnd.n2969 99.6594
R6883 gnd.n3011 gnd.n2970 99.6594
R6884 gnd.n3007 gnd.n2971 99.6594
R6885 gnd.n3003 gnd.n2972 99.6594
R6886 gnd.n3054 gnd.n3053 99.6594
R6887 gnd.n3819 gnd.n2457 99.6594
R6888 gnd.n3823 gnd.n2456 99.6594
R6889 gnd.n3827 gnd.n2455 99.6594
R6890 gnd.n3831 gnd.n2454 99.6594
R6891 gnd.n3835 gnd.n2453 99.6594
R6892 gnd.n3839 gnd.n2452 99.6594
R6893 gnd.n3843 gnd.n2451 99.6594
R6894 gnd.n3847 gnd.n2450 99.6594
R6895 gnd.n3851 gnd.n2449 99.6594
R6896 gnd.n3855 gnd.n2448 99.6594
R6897 gnd.n3859 gnd.n2447 99.6594
R6898 gnd.n3863 gnd.n2446 99.6594
R6899 gnd.n2486 gnd.n2445 99.6594
R6900 gnd.n1586 gnd.n1511 99.6594
R6901 gnd.n1588 gnd.n1587 99.6594
R6902 gnd.n1589 gnd.n1520 99.6594
R6903 gnd.n1591 gnd.n1527 99.6594
R6904 gnd.n1593 gnd.n1592 99.6594
R6905 gnd.n1594 gnd.n1536 99.6594
R6906 gnd.n1596 gnd.n1543 99.6594
R6907 gnd.n1598 gnd.n1597 99.6594
R6908 gnd.n5757 gnd.n5756 99.6594
R6909 gnd.n197 gnd.n194 99.6594
R6910 gnd.n254 gnd.n253 99.6594
R6911 gnd.n193 gnd.n187 99.6594
R6912 gnd.n261 gnd.n260 99.6594
R6913 gnd.n186 gnd.n180 99.6594
R6914 gnd.n268 gnd.n267 99.6594
R6915 gnd.n179 gnd.n173 99.6594
R6916 gnd.n275 gnd.n274 99.6594
R6917 gnd.n172 gnd.n169 99.6594
R6918 gnd.n3137 gnd.n3136 99.6594
R6919 gnd.n2896 gnd.n2874 99.6594
R6920 gnd.n2902 gnd.n2875 99.6594
R6921 gnd.n2906 gnd.n2876 99.6594
R6922 gnd.n2912 gnd.n2877 99.6594
R6923 gnd.n2916 gnd.n2878 99.6594
R6924 gnd.n2922 gnd.n2879 99.6594
R6925 gnd.n2880 gnd.n2864 99.6594
R6926 gnd.n3873 gnd.n2458 99.6594
R6927 gnd.n3877 gnd.n2459 99.6594
R6928 gnd.n3881 gnd.n2460 99.6594
R6929 gnd.n3885 gnd.n2461 99.6594
R6930 gnd.n3889 gnd.n2462 99.6594
R6931 gnd.n3893 gnd.n2463 99.6594
R6932 gnd.n3897 gnd.n2464 99.6594
R6933 gnd.n2467 gnd.n2465 99.6594
R6934 gnd.n4240 gnd.n3944 99.6594
R6935 gnd.n4232 gnd.n3906 99.6594
R6936 gnd.n4228 gnd.n3907 99.6594
R6937 gnd.n4224 gnd.n3908 99.6594
R6938 gnd.n4220 gnd.n3909 99.6594
R6939 gnd.n4216 gnd.n3910 99.6594
R6940 gnd.n4212 gnd.n3911 99.6594
R6941 gnd.n4208 gnd.n3912 99.6594
R6942 gnd.n4203 gnd.n3913 99.6594
R6943 gnd.n4199 gnd.n3914 99.6594
R6944 gnd.n4195 gnd.n3915 99.6594
R6945 gnd.n4191 gnd.n3916 99.6594
R6946 gnd.n4187 gnd.n3917 99.6594
R6947 gnd.n4183 gnd.n3918 99.6594
R6948 gnd.n4179 gnd.n3919 99.6594
R6949 gnd.n4175 gnd.n3920 99.6594
R6950 gnd.n4171 gnd.n3921 99.6594
R6951 gnd.n4167 gnd.n3922 99.6594
R6952 gnd.n4163 gnd.n3923 99.6594
R6953 gnd.n4159 gnd.n3924 99.6594
R6954 gnd.n4155 gnd.n3925 99.6594
R6955 gnd.n4151 gnd.n3926 99.6594
R6956 gnd.n4147 gnd.n3927 99.6594
R6957 gnd.n4143 gnd.n3928 99.6594
R6958 gnd.n4139 gnd.n3929 99.6594
R6959 gnd.n4135 gnd.n3930 99.6594
R6960 gnd.n4131 gnd.n3931 99.6594
R6961 gnd.n4127 gnd.n3932 99.6594
R6962 gnd.n4243 gnd.n4242 99.6594
R6963 gnd.n4578 gnd.n1156 99.6594
R6964 gnd.n4659 gnd.n1157 99.6594
R6965 gnd.n4657 gnd.n1158 99.6594
R6966 gnd.n4649 gnd.n1159 99.6594
R6967 gnd.n4647 gnd.n1160 99.6594
R6968 gnd.n4639 gnd.n1161 99.6594
R6969 gnd.n4637 gnd.n1162 99.6594
R6970 gnd.n4629 gnd.n1163 99.6594
R6971 gnd.n4627 gnd.n1164 99.6594
R6972 gnd.n4619 gnd.n1165 99.6594
R6973 gnd.n4591 gnd.n1166 99.6594
R6974 gnd.n4610 gnd.n1167 99.6594
R6975 gnd.n4608 gnd.n1168 99.6594
R6976 gnd.n4600 gnd.n1169 99.6594
R6977 gnd.n4598 gnd.n1170 99.6594
R6978 gnd.n6036 gnd.n1172 99.6594
R6979 gnd.n6040 gnd.n1173 99.6594
R6980 gnd.n6044 gnd.n1174 99.6594
R6981 gnd.n6048 gnd.n1175 99.6594
R6982 gnd.n6053 gnd.n1176 99.6594
R6983 gnd.n6057 gnd.n1177 99.6594
R6984 gnd.n6061 gnd.n1178 99.6594
R6985 gnd.n6065 gnd.n1179 99.6594
R6986 gnd.n6069 gnd.n1180 99.6594
R6987 gnd.n6073 gnd.n1181 99.6594
R6988 gnd.n6077 gnd.n1182 99.6594
R6989 gnd.n1184 gnd.n1183 99.6594
R6990 gnd.n6083 gnd.n1143 99.6594
R6991 gnd.n5754 gnd.n1601 99.6594
R6992 gnd.n5746 gnd.n1558 99.6594
R6993 gnd.n5742 gnd.n1559 99.6594
R6994 gnd.n5738 gnd.n1560 99.6594
R6995 gnd.n5734 gnd.n1561 99.6594
R6996 gnd.n5730 gnd.n1562 99.6594
R6997 gnd.n5726 gnd.n1563 99.6594
R6998 gnd.n5722 gnd.n1564 99.6594
R6999 gnd.n5717 gnd.n1565 99.6594
R7000 gnd.n5713 gnd.n1566 99.6594
R7001 gnd.n5709 gnd.n1567 99.6594
R7002 gnd.n5705 gnd.n1568 99.6594
R7003 gnd.n5700 gnd.n1570 99.6594
R7004 gnd.n5696 gnd.n1571 99.6594
R7005 gnd.n5692 gnd.n1572 99.6594
R7006 gnd.n5688 gnd.n1573 99.6594
R7007 gnd.n5684 gnd.n1574 99.6594
R7008 gnd.n5680 gnd.n1575 99.6594
R7009 gnd.n5676 gnd.n1576 99.6594
R7010 gnd.n5672 gnd.n1577 99.6594
R7011 gnd.n5668 gnd.n1578 99.6594
R7012 gnd.n5664 gnd.n1579 99.6594
R7013 gnd.n5660 gnd.n1580 99.6594
R7014 gnd.n5656 gnd.n1581 99.6594
R7015 gnd.n5652 gnd.n1582 99.6594
R7016 gnd.n5648 gnd.n1583 99.6594
R7017 gnd.n5644 gnd.n1584 99.6594
R7018 gnd.n5636 gnd.n1585 99.6594
R7019 gnd.n489 gnd.n488 99.6594
R7020 gnd.n480 gnd.n285 99.6594
R7021 gnd.n479 gnd.n478 99.6594
R7022 gnd.n470 gnd.n289 99.6594
R7023 gnd.n469 gnd.n468 99.6594
R7024 gnd.n460 gnd.n293 99.6594
R7025 gnd.n459 gnd.n458 99.6594
R7026 gnd.n450 gnd.n297 99.6594
R7027 gnd.n449 gnd.n448 99.6594
R7028 gnd.n440 gnd.n301 99.6594
R7029 gnd.n439 gnd.n438 99.6594
R7030 gnd.n430 gnd.n307 99.6594
R7031 gnd.n429 gnd.n428 99.6594
R7032 gnd.n420 gnd.n311 99.6594
R7033 gnd.n419 gnd.n418 99.6594
R7034 gnd.n410 gnd.n315 99.6594
R7035 gnd.n409 gnd.n408 99.6594
R7036 gnd.n400 gnd.n319 99.6594
R7037 gnd.n399 gnd.n398 99.6594
R7038 gnd.n390 gnd.n323 99.6594
R7039 gnd.n389 gnd.n388 99.6594
R7040 gnd.n380 gnd.n379 99.6594
R7041 gnd.n378 gnd.n377 99.6594
R7042 gnd.n369 gnd.n333 99.6594
R7043 gnd.n368 gnd.n367 99.6594
R7044 gnd.n359 gnd.n337 99.6594
R7045 gnd.n358 gnd.n357 99.6594
R7046 gnd.n349 gnd.n341 99.6594
R7047 gnd.n348 gnd.n347 99.6594
R7048 gnd.n2274 gnd.n2263 99.6594
R7049 gnd.n4450 gnd.n2275 99.6594
R7050 gnd.n4445 gnd.n2276 99.6594
R7051 gnd.n4458 gnd.n2277 99.6594
R7052 gnd.n4460 gnd.n2278 99.6594
R7053 gnd.n4467 gnd.n2279 99.6594
R7054 gnd.n4469 gnd.n2280 99.6594
R7055 gnd.n4479 gnd.n2281 99.6594
R7056 gnd.n4487 gnd.n2282 99.6594
R7057 gnd.n4489 gnd.n2283 99.6594
R7058 gnd.n4499 gnd.n2284 99.6594
R7059 gnd.n4507 gnd.n2285 99.6594
R7060 gnd.n4509 gnd.n2286 99.6594
R7061 gnd.n4521 gnd.n2287 99.6594
R7062 gnd.n4449 gnd.n2274 99.6594
R7063 gnd.n4444 gnd.n2275 99.6594
R7064 gnd.n4457 gnd.n2276 99.6594
R7065 gnd.n4459 gnd.n2277 99.6594
R7066 gnd.n4466 gnd.n2278 99.6594
R7067 gnd.n4468 gnd.n2279 99.6594
R7068 gnd.n4478 gnd.n2280 99.6594
R7069 gnd.n4486 gnd.n2281 99.6594
R7070 gnd.n4488 gnd.n2282 99.6594
R7071 gnd.n4498 gnd.n2283 99.6594
R7072 gnd.n4506 gnd.n2284 99.6594
R7073 gnd.n4508 gnd.n2285 99.6594
R7074 gnd.n4520 gnd.n2286 99.6594
R7075 gnd.n2288 gnd.n2287 99.6594
R7076 gnd.n1750 gnd.n1492 99.6594
R7077 gnd.n1752 gnd.n1497 99.6594
R7078 gnd.n1753 gnd.n1500 99.6594
R7079 gnd.n1755 gnd.n1502 99.6594
R7080 gnd.n1756 gnd.n1506 99.6594
R7081 gnd.n1758 gnd.n1757 99.6594
R7082 gnd.n1760 gnd.n1516 99.6594
R7083 gnd.n1761 gnd.n1523 99.6594
R7084 gnd.n1763 gnd.n1762 99.6594
R7085 gnd.n1765 gnd.n1532 99.6594
R7086 gnd.n1766 gnd.n1539 99.6594
R7087 gnd.n1768 gnd.n1767 99.6594
R7088 gnd.n1771 gnd.n1548 99.6594
R7089 gnd.n5529 gnd.n1749 99.6594
R7090 gnd.n1768 gnd.n1547 99.6594
R7091 gnd.n1766 gnd.n1540 99.6594
R7092 gnd.n1765 gnd.n1764 99.6594
R7093 gnd.n1763 gnd.n1531 99.6594
R7094 gnd.n1761 gnd.n1524 99.6594
R7095 gnd.n1760 gnd.n1759 99.6594
R7096 gnd.n1758 gnd.n1515 99.6594
R7097 gnd.n1756 gnd.n1507 99.6594
R7098 gnd.n1755 gnd.n1754 99.6594
R7099 gnd.n1753 gnd.n1501 99.6594
R7100 gnd.n1752 gnd.n1751 99.6594
R7101 gnd.n1750 gnd.n1496 99.6594
R7102 gnd.n5530 gnd.n5529 99.6594
R7103 gnd.n1771 gnd.n1770 99.6594
R7104 gnd.n4517 gnd.t135 98.63
R7105 gnd.n5758 gnd.t156 98.63
R7106 gnd.n2292 gnd.t175 98.63
R7107 gnd.n1621 gnd.t153 98.63
R7108 gnd.n1644 gnd.t141 98.63
R7109 gnd.n5638 gnd.t84 98.63
R7110 gnd.n282 gnd.t89 98.63
R7111 gnd.n304 gnd.t79 98.63
R7112 gnd.n326 gnd.t146 98.63
R7113 gnd.n200 gnd.t162 98.63
R7114 gnd.n3963 gnd.t118 98.63
R7115 gnd.n3985 gnd.t100 98.63
R7116 gnd.n4006 gnd.t124 98.63
R7117 gnd.n4024 gnd.t76 98.63
R7118 gnd.n1201 gnd.t165 98.63
R7119 gnd.n4576 gnd.t107 98.63
R7120 gnd.n4589 gnd.t130 98.63
R7121 gnd.n1549 gnd.t114 98.63
R7122 gnd.n1296 gnd.t169 96.6984
R7123 gnd.n1920 gnd.t93 96.6984
R7124 gnd.n5965 gnd.t104 96.6906
R7125 gnd.n1815 gnd.t143 96.6906
R7126 gnd.n1263 gnd.n1262 81.8399
R7127 gnd.n2925 gnd.t127 74.8376
R7128 gnd.n2483 gnd.t160 74.8376
R7129 gnd.n1297 gnd.t168 72.8438
R7130 gnd.n1921 gnd.t94 72.8438
R7131 gnd.n1264 gnd.n1257 72.8411
R7132 gnd.n1270 gnd.n1255 72.8411
R7133 gnd.n1832 gnd.n1831 72.8411
R7134 gnd.n4518 gnd.t134 72.836
R7135 gnd.n5966 gnd.t103 72.836
R7136 gnd.n1816 gnd.t144 72.836
R7137 gnd.n5759 gnd.t155 72.836
R7138 gnd.n2293 gnd.t176 72.836
R7139 gnd.n1622 gnd.t152 72.836
R7140 gnd.n1645 gnd.t140 72.836
R7141 gnd.n5639 gnd.t83 72.836
R7142 gnd.n283 gnd.t90 72.836
R7143 gnd.n305 gnd.t80 72.836
R7144 gnd.n327 gnd.t147 72.836
R7145 gnd.n201 gnd.t163 72.836
R7146 gnd.n3964 gnd.t117 72.836
R7147 gnd.n3986 gnd.t99 72.836
R7148 gnd.n4007 gnd.t123 72.836
R7149 gnd.n4025 gnd.t75 72.836
R7150 gnd.n1202 gnd.t166 72.836
R7151 gnd.n4577 gnd.t108 72.836
R7152 gnd.n4590 gnd.t131 72.836
R7153 gnd.n1550 gnd.t115 72.836
R7154 gnd.n1839 gnd.n1799 71.676
R7155 gnd.n1843 gnd.n1800 71.676
R7156 gnd.n1847 gnd.n1801 71.676
R7157 gnd.n1851 gnd.n1802 71.676
R7158 gnd.n1855 gnd.n1803 71.676
R7159 gnd.n1859 gnd.n1804 71.676
R7160 gnd.n1863 gnd.n1805 71.676
R7161 gnd.n1867 gnd.n1806 71.676
R7162 gnd.n1871 gnd.n1807 71.676
R7163 gnd.n1875 gnd.n1808 71.676
R7164 gnd.n1879 gnd.n1809 71.676
R7165 gnd.n1883 gnd.n1810 71.676
R7166 gnd.n1887 gnd.n1811 71.676
R7167 gnd.n1891 gnd.n1812 71.676
R7168 gnd.n1896 gnd.n1813 71.676
R7169 gnd.n1900 gnd.n1814 71.676
R7170 gnd.n5474 gnd.n1919 71.676
R7171 gnd.n5470 gnd.n1918 71.676
R7172 gnd.n5465 gnd.n1917 71.676
R7173 gnd.n5461 gnd.n1916 71.676
R7174 gnd.n5457 gnd.n1915 71.676
R7175 gnd.n5453 gnd.n1914 71.676
R7176 gnd.n5449 gnd.n1913 71.676
R7177 gnd.n5445 gnd.n1912 71.676
R7178 gnd.n5441 gnd.n1911 71.676
R7179 gnd.n5437 gnd.n1910 71.676
R7180 gnd.n5433 gnd.n1909 71.676
R7181 gnd.n5429 gnd.n1908 71.676
R7182 gnd.n5425 gnd.n1907 71.676
R7183 gnd.n5421 gnd.n1906 71.676
R7184 gnd.n5417 gnd.n1905 71.676
R7185 gnd.n5413 gnd.n1904 71.676
R7186 gnd.n5409 gnd.n1903 71.676
R7187 gnd.n6029 gnd.n6028 71.676
R7188 gnd.n6023 gnd.n1219 71.676
R7189 gnd.n6020 gnd.n1220 71.676
R7190 gnd.n6016 gnd.n1221 71.676
R7191 gnd.n6012 gnd.n1222 71.676
R7192 gnd.n6008 gnd.n1223 71.676
R7193 gnd.n6004 gnd.n1224 71.676
R7194 gnd.n6000 gnd.n1225 71.676
R7195 gnd.n5996 gnd.n1226 71.676
R7196 gnd.n5992 gnd.n1227 71.676
R7197 gnd.n5988 gnd.n1228 71.676
R7198 gnd.n5984 gnd.n1229 71.676
R7199 gnd.n5980 gnd.n1230 71.676
R7200 gnd.n5976 gnd.n1231 71.676
R7201 gnd.n5972 gnd.n1232 71.676
R7202 gnd.n5968 gnd.n1233 71.676
R7203 gnd.n1234 gnd.n1217 71.676
R7204 gnd.n1300 gnd.n1235 71.676
R7205 gnd.n1305 gnd.n1236 71.676
R7206 gnd.n1309 gnd.n1237 71.676
R7207 gnd.n1313 gnd.n1238 71.676
R7208 gnd.n1317 gnd.n1239 71.676
R7209 gnd.n1321 gnd.n1240 71.676
R7210 gnd.n1325 gnd.n1241 71.676
R7211 gnd.n1329 gnd.n1242 71.676
R7212 gnd.n1333 gnd.n1243 71.676
R7213 gnd.n1337 gnd.n1244 71.676
R7214 gnd.n1341 gnd.n1245 71.676
R7215 gnd.n1345 gnd.n1246 71.676
R7216 gnd.n1349 gnd.n1247 71.676
R7217 gnd.n1353 gnd.n1248 71.676
R7218 gnd.n1357 gnd.n1249 71.676
R7219 gnd.n6029 gnd.n1252 71.676
R7220 gnd.n6021 gnd.n1219 71.676
R7221 gnd.n6017 gnd.n1220 71.676
R7222 gnd.n6013 gnd.n1221 71.676
R7223 gnd.n6009 gnd.n1222 71.676
R7224 gnd.n6005 gnd.n1223 71.676
R7225 gnd.n6001 gnd.n1224 71.676
R7226 gnd.n5997 gnd.n1225 71.676
R7227 gnd.n5993 gnd.n1226 71.676
R7228 gnd.n5989 gnd.n1227 71.676
R7229 gnd.n5985 gnd.n1228 71.676
R7230 gnd.n5981 gnd.n1229 71.676
R7231 gnd.n5977 gnd.n1230 71.676
R7232 gnd.n5973 gnd.n1231 71.676
R7233 gnd.n5969 gnd.n1232 71.676
R7234 gnd.n6032 gnd.n6031 71.676
R7235 gnd.n1299 gnd.n1234 71.676
R7236 gnd.n1304 gnd.n1235 71.676
R7237 gnd.n1308 gnd.n1236 71.676
R7238 gnd.n1312 gnd.n1237 71.676
R7239 gnd.n1316 gnd.n1238 71.676
R7240 gnd.n1320 gnd.n1239 71.676
R7241 gnd.n1324 gnd.n1240 71.676
R7242 gnd.n1328 gnd.n1241 71.676
R7243 gnd.n1332 gnd.n1242 71.676
R7244 gnd.n1336 gnd.n1243 71.676
R7245 gnd.n1340 gnd.n1244 71.676
R7246 gnd.n1344 gnd.n1245 71.676
R7247 gnd.n1348 gnd.n1246 71.676
R7248 gnd.n1352 gnd.n1247 71.676
R7249 gnd.n1356 gnd.n1248 71.676
R7250 gnd.n1360 gnd.n1249 71.676
R7251 gnd.n5412 gnd.n1903 71.676
R7252 gnd.n5416 gnd.n1904 71.676
R7253 gnd.n5420 gnd.n1905 71.676
R7254 gnd.n5424 gnd.n1906 71.676
R7255 gnd.n5428 gnd.n1907 71.676
R7256 gnd.n5432 gnd.n1908 71.676
R7257 gnd.n5436 gnd.n1909 71.676
R7258 gnd.n5440 gnd.n1910 71.676
R7259 gnd.n5444 gnd.n1911 71.676
R7260 gnd.n5448 gnd.n1912 71.676
R7261 gnd.n5452 gnd.n1913 71.676
R7262 gnd.n5456 gnd.n1914 71.676
R7263 gnd.n5460 gnd.n1915 71.676
R7264 gnd.n5464 gnd.n1916 71.676
R7265 gnd.n5469 gnd.n1917 71.676
R7266 gnd.n5473 gnd.n1918 71.676
R7267 gnd.n1902 gnd.n1901 71.676
R7268 gnd.n1897 gnd.n1814 71.676
R7269 gnd.n1892 gnd.n1813 71.676
R7270 gnd.n1888 gnd.n1812 71.676
R7271 gnd.n1884 gnd.n1811 71.676
R7272 gnd.n1880 gnd.n1810 71.676
R7273 gnd.n1876 gnd.n1809 71.676
R7274 gnd.n1872 gnd.n1808 71.676
R7275 gnd.n1868 gnd.n1807 71.676
R7276 gnd.n1864 gnd.n1806 71.676
R7277 gnd.n1860 gnd.n1805 71.676
R7278 gnd.n1856 gnd.n1804 71.676
R7279 gnd.n1852 gnd.n1803 71.676
R7280 gnd.n1848 gnd.n1802 71.676
R7281 gnd.n1844 gnd.n1801 71.676
R7282 gnd.n1840 gnd.n1800 71.676
R7283 gnd.n1799 gnd.n1797 71.676
R7284 gnd.n8 gnd.t307 69.1507
R7285 gnd.n14 gnd.t43 68.4792
R7286 gnd.n13 gnd.t5 68.4792
R7287 gnd.n12 gnd.t56 68.4792
R7288 gnd.n11 gnd.t327 68.4792
R7289 gnd.n10 gnd.t309 68.4792
R7290 gnd.n9 gnd.t54 68.4792
R7291 gnd.n8 gnd.t14 68.4792
R7292 gnd.n3052 gnd.n2956 64.369
R7293 gnd.n6840 gnd.n136 64.0315
R7294 gnd.n4241 gnd.n2430 63.0944
R7295 gnd.n6969 gnd.n165 63.0944
R7296 gnd.n1302 gnd.n1297 59.5399
R7297 gnd.n5467 gnd.n1921 59.5399
R7298 gnd.n5967 gnd.n5966 59.5399
R7299 gnd.n1894 gnd.n1816 59.5399
R7300 gnd.n5964 gnd.n1273 59.1804
R7301 gnd.n3905 gnd.n2443 57.3586
R7302 gnd.n2711 gnd.t242 56.407
R7303 gnd.n2676 gnd.t291 56.407
R7304 gnd.n2687 gnd.t201 56.407
R7305 gnd.n2699 gnd.t282 56.407
R7306 gnd.n52 gnd.t222 56.407
R7307 gnd.n17 gnd.t208 56.407
R7308 gnd.n28 gnd.t300 56.407
R7309 gnd.n40 gnd.t257 56.407
R7310 gnd.n2720 gnd.t268 55.8337
R7311 gnd.n2685 gnd.t197 55.8337
R7312 gnd.n2696 gnd.t298 55.8337
R7313 gnd.n2708 gnd.t204 55.8337
R7314 gnd.n61 gnd.t240 55.8337
R7315 gnd.n26 gnd.t232 55.8337
R7316 gnd.n37 gnd.t283 55.8337
R7317 gnd.n49 gnd.t279 55.8337
R7318 gnd.n1261 gnd.n1260 54.358
R7319 gnd.n1829 gnd.n1828 54.358
R7320 gnd.n2711 gnd.n2710 53.0052
R7321 gnd.n2713 gnd.n2712 53.0052
R7322 gnd.n2715 gnd.n2714 53.0052
R7323 gnd.n2717 gnd.n2716 53.0052
R7324 gnd.n2719 gnd.n2718 53.0052
R7325 gnd.n2676 gnd.n2675 53.0052
R7326 gnd.n2678 gnd.n2677 53.0052
R7327 gnd.n2680 gnd.n2679 53.0052
R7328 gnd.n2682 gnd.n2681 53.0052
R7329 gnd.n2684 gnd.n2683 53.0052
R7330 gnd.n2687 gnd.n2686 53.0052
R7331 gnd.n2689 gnd.n2688 53.0052
R7332 gnd.n2691 gnd.n2690 53.0052
R7333 gnd.n2693 gnd.n2692 53.0052
R7334 gnd.n2695 gnd.n2694 53.0052
R7335 gnd.n2699 gnd.n2698 53.0052
R7336 gnd.n2701 gnd.n2700 53.0052
R7337 gnd.n2703 gnd.n2702 53.0052
R7338 gnd.n2705 gnd.n2704 53.0052
R7339 gnd.n2707 gnd.n2706 53.0052
R7340 gnd.n60 gnd.n59 53.0052
R7341 gnd.n58 gnd.n57 53.0052
R7342 gnd.n56 gnd.n55 53.0052
R7343 gnd.n54 gnd.n53 53.0052
R7344 gnd.n52 gnd.n51 53.0052
R7345 gnd.n25 gnd.n24 53.0052
R7346 gnd.n23 gnd.n22 53.0052
R7347 gnd.n21 gnd.n20 53.0052
R7348 gnd.n19 gnd.n18 53.0052
R7349 gnd.n17 gnd.n16 53.0052
R7350 gnd.n36 gnd.n35 53.0052
R7351 gnd.n34 gnd.n33 53.0052
R7352 gnd.n32 gnd.n31 53.0052
R7353 gnd.n30 gnd.n29 53.0052
R7354 gnd.n28 gnd.n27 53.0052
R7355 gnd.n48 gnd.n47 53.0052
R7356 gnd.n46 gnd.n45 53.0052
R7357 gnd.n44 gnd.n43 53.0052
R7358 gnd.n42 gnd.n41 53.0052
R7359 gnd.n40 gnd.n39 53.0052
R7360 gnd.n1820 gnd.n1819 52.4801
R7361 gnd.n3757 gnd.t26 52.3082
R7362 gnd.n3725 gnd.t47 52.3082
R7363 gnd.n3693 gnd.t49 52.3082
R7364 gnd.n3662 gnd.t318 52.3082
R7365 gnd.n3630 gnd.t63 52.3082
R7366 gnd.n3598 gnd.t37 52.3082
R7367 gnd.n3566 gnd.t41 52.3082
R7368 gnd.n3535 gnd.t311 52.3082
R7369 gnd.n3587 gnd.n3555 51.4173
R7370 gnd.n3651 gnd.n3650 50.455
R7371 gnd.n3619 gnd.n3618 50.455
R7372 gnd.n3587 gnd.n3586 50.455
R7373 gnd.n5702 gnd.n1631 45.6325
R7374 gnd.n6034 gnd.n6033 45.6325
R7375 gnd.n2999 gnd.n2998 45.1884
R7376 gnd.n2509 gnd.n2508 45.1884
R7377 gnd.n1836 gnd.n1835 44.3322
R7378 gnd.n1264 gnd.n1263 44.3189
R7379 gnd.n4519 gnd.n4518 42.2793
R7380 gnd.n5760 gnd.n5759 42.2793
R7381 gnd.n3000 gnd.n2999 42.2793
R7382 gnd.n2510 gnd.n2509 42.2793
R7383 gnd.n2926 gnd.n2925 42.2793
R7384 gnd.n3872 gnd.n2483 42.2793
R7385 gnd.n2294 gnd.n2293 42.2793
R7386 gnd.n5719 gnd.n1622 42.2793
R7387 gnd.n5682 gnd.n1645 42.2793
R7388 gnd.n5642 gnd.n5639 42.2793
R7389 gnd.n284 gnd.n283 42.2793
R7390 gnd.n306 gnd.n305 42.2793
R7391 gnd.n328 gnd.n327 42.2793
R7392 gnd.n250 gnd.n201 42.2793
R7393 gnd.n4205 gnd.n3964 42.2793
R7394 gnd.n4165 gnd.n3986 42.2793
R7395 gnd.n4126 gnd.n4007 42.2793
R7396 gnd.n4026 gnd.n4025 42.2793
R7397 gnd.n6051 gnd.n1202 42.2793
R7398 gnd.n4667 gnd.n4577 42.2793
R7399 gnd.n4618 gnd.n4590 42.2793
R7400 gnd.n1551 gnd.n1550 42.2793
R7401 gnd.n1262 gnd.n1261 41.6274
R7402 gnd.n1830 gnd.n1829 41.6274
R7403 gnd.n1271 gnd.n1270 40.8975
R7404 gnd.n1833 gnd.n1832 40.8975
R7405 gnd.n1270 gnd.n1269 35.055
R7406 gnd.n1265 gnd.n1264 35.055
R7407 gnd.n1822 gnd.n1821 35.055
R7408 gnd.n1832 gnd.n1818 35.055
R7409 gnd.n6309 gnd.n6308 34.6735
R7410 gnd.n6308 gnd.n6307 34.6735
R7411 gnd.n6307 gnd.n884 34.6735
R7412 gnd.n6301 gnd.n884 34.6735
R7413 gnd.n6301 gnd.n6300 34.6735
R7414 gnd.n6300 gnd.n6299 34.6735
R7415 gnd.n6299 gnd.n891 34.6735
R7416 gnd.n6293 gnd.n891 34.6735
R7417 gnd.n6293 gnd.n6292 34.6735
R7418 gnd.n6292 gnd.n6291 34.6735
R7419 gnd.n6291 gnd.n899 34.6735
R7420 gnd.n6285 gnd.n899 34.6735
R7421 gnd.n6285 gnd.n6284 34.6735
R7422 gnd.n6284 gnd.n6283 34.6735
R7423 gnd.n6283 gnd.n907 34.6735
R7424 gnd.n6277 gnd.n907 34.6735
R7425 gnd.n6277 gnd.n6276 34.6735
R7426 gnd.n6276 gnd.n6275 34.6735
R7427 gnd.n6275 gnd.n915 34.6735
R7428 gnd.n6269 gnd.n915 34.6735
R7429 gnd.n6269 gnd.n6268 34.6735
R7430 gnd.n6268 gnd.n6267 34.6735
R7431 gnd.n6267 gnd.n923 34.6735
R7432 gnd.n6261 gnd.n923 34.6735
R7433 gnd.n6261 gnd.n6260 34.6735
R7434 gnd.n6260 gnd.n6259 34.6735
R7435 gnd.n6259 gnd.n931 34.6735
R7436 gnd.n6253 gnd.n931 34.6735
R7437 gnd.n6253 gnd.n6252 34.6735
R7438 gnd.n6252 gnd.n6251 34.6735
R7439 gnd.n6251 gnd.n939 34.6735
R7440 gnd.n6245 gnd.n939 34.6735
R7441 gnd.n6245 gnd.n6244 34.6735
R7442 gnd.n6244 gnd.n6243 34.6735
R7443 gnd.n6243 gnd.n947 34.6735
R7444 gnd.n6237 gnd.n947 34.6735
R7445 gnd.n6237 gnd.n6236 34.6735
R7446 gnd.n6236 gnd.n6235 34.6735
R7447 gnd.n6235 gnd.n955 34.6735
R7448 gnd.n6229 gnd.n955 34.6735
R7449 gnd.n6229 gnd.n6228 34.6735
R7450 gnd.n6228 gnd.n6227 34.6735
R7451 gnd.n6227 gnd.n963 34.6735
R7452 gnd.n6221 gnd.n963 34.6735
R7453 gnd.n6221 gnd.n6220 34.6735
R7454 gnd.n6220 gnd.n6219 34.6735
R7455 gnd.n6219 gnd.n971 34.6735
R7456 gnd.n6213 gnd.n971 34.6735
R7457 gnd.n6213 gnd.n6212 34.6735
R7458 gnd.n6212 gnd.n6211 34.6735
R7459 gnd.n6211 gnd.n979 34.6735
R7460 gnd.n6205 gnd.n979 34.6735
R7461 gnd.n6205 gnd.n6204 34.6735
R7462 gnd.n6204 gnd.n6203 34.6735
R7463 gnd.n6203 gnd.n987 34.6735
R7464 gnd.n6197 gnd.n987 34.6735
R7465 gnd.n6197 gnd.n6196 34.6735
R7466 gnd.n6196 gnd.n6195 34.6735
R7467 gnd.n6195 gnd.n995 34.6735
R7468 gnd.n6189 gnd.n995 34.6735
R7469 gnd.n6189 gnd.n6188 34.6735
R7470 gnd.n6188 gnd.n6187 34.6735
R7471 gnd.n6187 gnd.n1003 34.6735
R7472 gnd.n6181 gnd.n1003 34.6735
R7473 gnd.n6181 gnd.n6180 34.6735
R7474 gnd.n6180 gnd.n6179 34.6735
R7475 gnd.n6179 gnd.n1011 34.6735
R7476 gnd.n6173 gnd.n1011 34.6735
R7477 gnd.n6173 gnd.n6172 34.6735
R7478 gnd.n6172 gnd.n6171 34.6735
R7479 gnd.n6171 gnd.n1019 34.6735
R7480 gnd.n6165 gnd.n1019 34.6735
R7481 gnd.n6165 gnd.n6164 34.6735
R7482 gnd.n6164 gnd.n6163 34.6735
R7483 gnd.n6163 gnd.n1027 34.6735
R7484 gnd.n6157 gnd.n1027 34.6735
R7485 gnd.n6157 gnd.n6156 34.6735
R7486 gnd.n6156 gnd.n6155 34.6735
R7487 gnd.n6155 gnd.n1035 34.6735
R7488 gnd.n6149 gnd.n1035 34.6735
R7489 gnd.n6149 gnd.n6148 34.6735
R7490 gnd.n6148 gnd.n6147 34.6735
R7491 gnd.n6147 gnd.n1043 34.6735
R7492 gnd.n5410 gnd.n5408 32.9371
R7493 gnd.n1363 gnd.n1359 32.9371
R7494 gnd.n3062 gnd.n2956 31.8661
R7495 gnd.n3062 gnd.n3061 31.8661
R7496 gnd.n3070 gnd.n2945 31.8661
R7497 gnd.n3078 gnd.n2945 31.8661
R7498 gnd.n3078 gnd.n2939 31.8661
R7499 gnd.n3086 gnd.n2939 31.8661
R7500 gnd.n3086 gnd.n2932 31.8661
R7501 gnd.n3124 gnd.n2932 31.8661
R7502 gnd.n3134 gnd.n2865 31.8661
R7503 gnd.n4251 gnd.n2430 31.8661
R7504 gnd.n4259 gnd.n2422 31.8661
R7505 gnd.n4259 gnd.n2411 31.8661
R7506 gnd.n4271 gnd.n2411 31.8661
R7507 gnd.n4271 gnd.n2414 31.8661
R7508 gnd.n4279 gnd.n2394 31.8661
R7509 gnd.n4291 gnd.n2394 31.8661
R7510 gnd.n4299 gnd.n2386 31.8661
R7511 gnd.n4311 gnd.n2375 31.8661
R7512 gnd.n4311 gnd.n2378 31.8661
R7513 gnd.n4320 gnd.n2358 31.8661
R7514 gnd.n4332 gnd.n2358 31.8661
R7515 gnd.n4340 gnd.n2352 31.8661
R7516 gnd.n4359 gnd.n2339 31.8661
R7517 gnd.n4359 gnd.n2342 31.8661
R7518 gnd.n4367 gnd.n1050 31.8661
R7519 gnd.n4713 gnd.n1144 31.8661
R7520 gnd.n2273 gnd.n1155 31.8661
R7521 gnd.n4738 gnd.n2273 31.8661
R7522 gnd.n4738 gnd.n2264 31.8661
R7523 gnd.n4755 gnd.n2264 31.8661
R7524 gnd.n4755 gnd.n2265 31.8661
R7525 gnd.n5823 gnd.n1488 31.8661
R7526 gnd.n5823 gnd.n1490 31.8661
R7527 gnd.n5528 gnd.n1490 31.8661
R7528 gnd.n5528 gnd.n1772 31.8661
R7529 gnd.n1772 gnd.n1557 31.8661
R7530 gnd.n1667 gnd.n1599 31.8661
R7531 gnd.n6910 gnd.n509 31.8661
R7532 gnd.n6918 gnd.n499 31.8661
R7533 gnd.n6927 gnd.n499 31.8661
R7534 gnd.n7025 gnd.n70 31.8661
R7535 gnd.n7017 gnd.n85 31.8661
R7536 gnd.n7017 gnd.n88 31.8661
R7537 gnd.n7011 gnd.n99 31.8661
R7538 gnd.n7005 gnd.n99 31.8661
R7539 gnd.n6999 gnd.n114 31.8661
R7540 gnd.n6993 gnd.n124 31.8661
R7541 gnd.n6993 gnd.n127 31.8661
R7542 gnd.n6981 gnd.n144 31.8661
R7543 gnd.n6981 gnd.n147 31.8661
R7544 gnd.n6975 gnd.n147 31.8661
R7545 gnd.n6969 gnd.n162 31.8661
R7546 gnd.t218 gnd.n2352 31.5474
R7547 gnd.t189 gnd.n70 31.5474
R7548 gnd.t233 gnd.n2386 30.9101
R7549 gnd.n6999 gnd.t191 30.9101
R7550 gnd.n6987 gnd.n136 28.6795
R7551 gnd.n6084 gnd.n1155 27.4049
R7552 gnd.n5755 gnd.n1557 27.4049
R7553 gnd.n6140 gnd.n1053 26.7676
R7554 gnd.n4376 gnd.n1062 26.7676
R7555 gnd.n4395 gnd.n1073 26.7676
R7556 gnd.n6128 gnd.n1076 26.7676
R7557 gnd.n6122 gnd.n1087 26.7676
R7558 gnd.n4422 gnd.n4421 26.7676
R7559 gnd.n6116 gnd.n1096 26.7676
R7560 gnd.n4430 gnd.n1104 26.7676
R7561 gnd.n4690 gnd.n1113 26.7676
R7562 gnd.n6104 gnd.n1116 26.7676
R7563 gnd.n4437 gnd.n1124 26.7676
R7564 gnd.n6098 gnd.n1127 26.7676
R7565 gnd.n6092 gnd.n1137 26.7676
R7566 gnd.n4714 gnd.n4713 26.7676
R7567 gnd.n5634 gnd.n1667 26.7676
R7568 gnd.n5572 gnd.n1669 26.7676
R7569 gnd.n5537 gnd.n1678 26.7676
R7570 gnd.n5620 gnd.n1691 26.7676
R7571 gnd.n5543 gnd.n1694 26.7676
R7572 gnd.n5614 gnd.n1704 26.7676
R7573 gnd.n5608 gnd.n1716 26.7676
R7574 gnd.n5601 gnd.n1719 26.7676
R7575 gnd.n5600 gnd.n1732 26.7676
R7576 gnd.n6864 gnd.n546 26.7676
R7577 gnd.n6875 gnd.n536 26.7676
R7578 gnd.n6857 gnd.n538 26.7676
R7579 gnd.n6897 gnd.n522 26.7676
R7580 gnd.n6902 gnd.n517 26.7676
R7581 gnd.n4518 gnd.n4517 25.7944
R7582 gnd.n5759 gnd.n5758 25.7944
R7583 gnd.n2925 gnd.n2924 25.7944
R7584 gnd.n2483 gnd.n2482 25.7944
R7585 gnd.n2293 gnd.n2292 25.7944
R7586 gnd.n1622 gnd.n1621 25.7944
R7587 gnd.n1645 gnd.n1644 25.7944
R7588 gnd.n5639 gnd.n5638 25.7944
R7589 gnd.n283 gnd.n282 25.7944
R7590 gnd.n305 gnd.n304 25.7944
R7591 gnd.n327 gnd.n326 25.7944
R7592 gnd.n201 gnd.n200 25.7944
R7593 gnd.n3964 gnd.n3963 25.7944
R7594 gnd.n3986 gnd.n3985 25.7944
R7595 gnd.n4007 gnd.n4006 25.7944
R7596 gnd.n4025 gnd.n4024 25.7944
R7597 gnd.n1202 gnd.n1201 25.7944
R7598 gnd.n4577 gnd.n4576 25.7944
R7599 gnd.n4590 gnd.n4589 25.7944
R7600 gnd.n1550 gnd.n1549 25.7944
R7601 gnd.n3146 gnd.n2866 24.8557
R7602 gnd.n3156 gnd.n2849 24.8557
R7603 gnd.n2852 gnd.n2840 24.8557
R7604 gnd.n3177 gnd.n2841 24.8557
R7605 gnd.n3187 gnd.n2821 24.8557
R7606 gnd.n3197 gnd.n3196 24.8557
R7607 gnd.n2807 gnd.n2805 24.8557
R7608 gnd.n3228 gnd.n3227 24.8557
R7609 gnd.n3243 gnd.n2790 24.8557
R7610 gnd.n3297 gnd.n2729 24.8557
R7611 gnd.n3253 gnd.n2730 24.8557
R7612 gnd.n3290 gnd.n2741 24.8557
R7613 gnd.n2779 gnd.n2778 24.8557
R7614 gnd.n3284 gnd.n3283 24.8557
R7615 gnd.n2765 gnd.n2752 24.8557
R7616 gnd.n3323 gnd.n3322 24.8557
R7617 gnd.n3333 gnd.n2661 24.8557
R7618 gnd.n3345 gnd.n2653 24.8557
R7619 gnd.n3344 gnd.n2641 24.8557
R7620 gnd.n3363 gnd.n3362 24.8557
R7621 gnd.n3373 gnd.n2634 24.8557
R7622 gnd.n3384 gnd.n2622 24.8557
R7623 gnd.n3408 gnd.n3407 24.8557
R7624 gnd.n3419 gnd.n2605 24.8557
R7625 gnd.n3418 gnd.n2607 24.8557
R7626 gnd.n3430 gnd.n2598 24.8557
R7627 gnd.n3448 gnd.n3447 24.8557
R7628 gnd.n2589 gnd.n2578 24.8557
R7629 gnd.n3469 gnd.n2566 24.8557
R7630 gnd.n3497 gnd.n3496 24.8557
R7631 gnd.n3508 gnd.n2551 24.8557
R7632 gnd.n3520 gnd.n2544 24.8557
R7633 gnd.n3792 gnd.n3791 24.8557
R7634 gnd.n3814 gnd.n2517 24.8557
R7635 gnd.n1297 gnd.n1296 23.855
R7636 gnd.n1921 gnd.n1920 23.855
R7637 gnd.n5966 gnd.n5965 23.855
R7638 gnd.n1816 gnd.n1815 23.855
R7639 gnd.n3167 gnd.t310 23.2624
R7640 gnd.n6030 gnd.n1250 23.2624
R7641 gnd.n5476 gnd.n5475 23.2624
R7642 gnd.n2868 gnd.t126 22.6251
R7643 gnd.n4299 gnd.t224 21.9878
R7644 gnd.n114 gnd.t253 21.9878
R7645 gnd.n6141 gnd.t205 21.6691
R7646 gnd.n5952 gnd.n1292 21.6691
R7647 gnd.n5940 gnd.n1377 21.6691
R7648 gnd.n4815 gnd.n2243 21.6691
R7649 gnd.n4877 gnd.n2232 21.6691
R7650 gnd.n4852 gnd.n2223 21.6691
R7651 gnd.n4959 gnd.n2176 21.6691
R7652 gnd.n4987 gnd.n2162 21.6691
R7653 gnd.n4993 gnd.n2158 21.6691
R7654 gnd.n5011 gnd.n2142 21.6691
R7655 gnd.n5038 gnd.n2130 21.6691
R7656 gnd.n5031 gnd.n2121 21.6691
R7657 gnd.n5096 gnd.n2099 21.6691
R7658 gnd.n5106 gnd.n2099 21.6691
R7659 gnd.n5120 gnd.n5119 21.6691
R7660 gnd.n5163 gnd.n5162 21.6691
R7661 gnd.n5156 gnd.n2057 21.6691
R7662 gnd.n5198 gnd.n2049 21.6691
R7663 gnd.n5209 gnd.n2044 21.6691
R7664 gnd.n5275 gnd.n2010 21.6691
R7665 gnd.n5303 gnd.n1995 21.6691
R7666 gnd.n5321 gnd.n1978 21.6691
R7667 gnd.n5349 gnd.n1957 21.6691
R7668 gnd.n5360 gnd.n1931 21.6691
R7669 gnd.n5404 gnd.n1784 21.6691
R7670 gnd.n6848 gnd.t187 21.6691
R7671 gnd.t317 gnd.n2873 21.3504
R7672 gnd.n4340 gnd.t258 21.3504
R7673 gnd.n4367 gnd.t246 21.3504
R7674 gnd.n6910 gnd.t216 21.3504
R7675 gnd.n7025 gnd.t237 21.3504
R7676 gnd.n3518 gnd.n1043 20.8043
R7677 gnd.n5964 gnd.n5963 20.7615
R7678 gnd.n1836 gnd.n1796 20.7615
R7679 gnd.t59 gnd.n2579 20.7131
R7680 gnd.n4320 gnd.t244 20.7131
R7681 gnd.n6134 gnd.t194 20.7131
R7682 gnd.n6883 gnd.t220 20.7131
R7683 gnd.t213 gnd.n88 20.7131
R7684 gnd.n5960 gnd.t68 20.3945
R7685 gnd.n5958 gnd.n1280 20.3945
R7686 gnd.n5946 gnd.n1371 20.3945
R7687 gnd.n2185 gnd.n2184 20.3945
R7688 gnd.n4930 gnd.n2172 20.3945
R7689 gnd.n5089 gnd.n2108 20.3945
R7690 gnd.n2102 gnd.n2094 20.3945
R7691 gnd.n5268 gnd.n2017 20.3945
R7692 gnd.n5283 gnd.n2003 20.3945
R7693 gnd.t57 gnd.n2614 20.0758
R7694 gnd.n4279 gnd.t196 20.0758
R7695 gnd.n6110 gnd.t200 20.0758
R7696 gnd.t92 gnd.t42 20.0758
R7697 gnd.n5550 gnd.t207 20.0758
R7698 gnd.t231 gnd.n127 20.0758
R7699 gnd.n1259 gnd.t69 19.8005
R7700 gnd.n1259 gnd.t97 19.8005
R7701 gnd.n1258 gnd.t179 19.8005
R7702 gnd.n1258 gnd.t72 19.8005
R7703 gnd.n1827 gnd.t121 19.8005
R7704 gnd.n1827 gnd.t66 19.8005
R7705 gnd.n1826 gnd.t111 19.8005
R7706 gnd.n1826 gnd.t87 19.8005
R7707 gnd.n1255 gnd.n1254 19.5087
R7708 gnd.n1268 gnd.n1255 19.5087
R7709 gnd.n1266 gnd.n1257 19.5087
R7710 gnd.n1831 gnd.n1825 19.5087
R7711 gnd.n3334 gnd.t61 19.4385
R7712 gnd.n4733 gnd.n4732 19.3944
R7713 gnd.n4732 gnd.n4731 19.3944
R7714 gnd.n4731 gnd.n4724 19.3944
R7715 gnd.n4727 gnd.n4724 19.3944
R7716 gnd.n4727 gnd.n2256 19.3944
R7717 gnd.n4779 gnd.n2256 19.3944
R7718 gnd.n4779 gnd.n2253 19.3944
R7719 gnd.n4786 gnd.n2253 19.3944
R7720 gnd.n4786 gnd.n2254 19.3944
R7721 gnd.n4782 gnd.n2254 19.3944
R7722 gnd.n4782 gnd.n1397 19.3944
R7723 gnd.n5931 gnd.n1397 19.3944
R7724 gnd.n5931 gnd.n1398 19.3944
R7725 gnd.n5927 gnd.n1398 19.3944
R7726 gnd.n5927 gnd.n5926 19.3944
R7727 gnd.n5926 gnd.n5925 19.3944
R7728 gnd.n5925 gnd.n1404 19.3944
R7729 gnd.n5921 gnd.n1404 19.3944
R7730 gnd.n5921 gnd.n5920 19.3944
R7731 gnd.n5920 gnd.n5919 19.3944
R7732 gnd.n5919 gnd.n1409 19.3944
R7733 gnd.n5915 gnd.n1409 19.3944
R7734 gnd.n5915 gnd.n5914 19.3944
R7735 gnd.n5914 gnd.n5913 19.3944
R7736 gnd.n5913 gnd.n1414 19.3944
R7737 gnd.n5909 gnd.n1414 19.3944
R7738 gnd.n5909 gnd.n5908 19.3944
R7739 gnd.n5908 gnd.n5907 19.3944
R7740 gnd.n5907 gnd.n1419 19.3944
R7741 gnd.n5903 gnd.n1419 19.3944
R7742 gnd.n5903 gnd.n5902 19.3944
R7743 gnd.n5902 gnd.n5901 19.3944
R7744 gnd.n5901 gnd.n1424 19.3944
R7745 gnd.n5897 gnd.n1424 19.3944
R7746 gnd.n5897 gnd.n5896 19.3944
R7747 gnd.n5896 gnd.n5895 19.3944
R7748 gnd.n5895 gnd.n1429 19.3944
R7749 gnd.n5891 gnd.n1429 19.3944
R7750 gnd.n5891 gnd.n5890 19.3944
R7751 gnd.n5890 gnd.n5889 19.3944
R7752 gnd.n5889 gnd.n1434 19.3944
R7753 gnd.n5885 gnd.n1434 19.3944
R7754 gnd.n5885 gnd.n5884 19.3944
R7755 gnd.n5884 gnd.n5883 19.3944
R7756 gnd.n5883 gnd.n1439 19.3944
R7757 gnd.n5879 gnd.n1439 19.3944
R7758 gnd.n5879 gnd.n5878 19.3944
R7759 gnd.n5878 gnd.n5877 19.3944
R7760 gnd.n5877 gnd.n1444 19.3944
R7761 gnd.n5873 gnd.n1444 19.3944
R7762 gnd.n5873 gnd.n5872 19.3944
R7763 gnd.n5872 gnd.n5871 19.3944
R7764 gnd.n5871 gnd.n1449 19.3944
R7765 gnd.n5867 gnd.n1449 19.3944
R7766 gnd.n5867 gnd.n5866 19.3944
R7767 gnd.n5866 gnd.n5865 19.3944
R7768 gnd.n5865 gnd.n1454 19.3944
R7769 gnd.n5861 gnd.n1454 19.3944
R7770 gnd.n5861 gnd.n5860 19.3944
R7771 gnd.n5860 gnd.n5859 19.3944
R7772 gnd.n5859 gnd.n1459 19.3944
R7773 gnd.n5855 gnd.n1459 19.3944
R7774 gnd.n5855 gnd.n5854 19.3944
R7775 gnd.n5854 gnd.n5853 19.3944
R7776 gnd.n5853 gnd.n1464 19.3944
R7777 gnd.n5849 gnd.n1464 19.3944
R7778 gnd.n5849 gnd.n5848 19.3944
R7779 gnd.n5848 gnd.n5847 19.3944
R7780 gnd.n5847 gnd.n1469 19.3944
R7781 gnd.n5843 gnd.n1469 19.3944
R7782 gnd.n5843 gnd.n5842 19.3944
R7783 gnd.n5842 gnd.n5841 19.3944
R7784 gnd.n5841 gnd.n1474 19.3944
R7785 gnd.n5837 gnd.n1474 19.3944
R7786 gnd.n5837 gnd.n5836 19.3944
R7787 gnd.n5836 gnd.n5835 19.3944
R7788 gnd.n5835 gnd.n1479 19.3944
R7789 gnd.n5831 gnd.n1479 19.3944
R7790 gnd.n5831 gnd.n5830 19.3944
R7791 gnd.n5830 gnd.n5829 19.3944
R7792 gnd.n5829 gnd.n1484 19.3944
R7793 gnd.n5825 gnd.n1484 19.3944
R7794 gnd.n4523 gnd.n4522 19.3944
R7795 gnd.n4522 gnd.n2289 19.3944
R7796 gnd.n4736 gnd.n2289 19.3944
R7797 gnd.n4448 gnd.n4447 19.3944
R7798 gnd.n4451 gnd.n4448 19.3944
R7799 gnd.n4451 gnd.n4443 19.3944
R7800 gnd.n4455 gnd.n4443 19.3944
R7801 gnd.n4456 gnd.n4455 19.3944
R7802 gnd.n4572 gnd.n4456 19.3944
R7803 gnd.n4572 gnd.n4571 19.3944
R7804 gnd.n4571 gnd.n4570 19.3944
R7805 gnd.n4570 gnd.n4461 19.3944
R7806 gnd.n4563 gnd.n4461 19.3944
R7807 gnd.n4563 gnd.n4562 19.3944
R7808 gnd.n4562 gnd.n4470 19.3944
R7809 gnd.n4555 gnd.n4470 19.3944
R7810 gnd.n4555 gnd.n4554 19.3944
R7811 gnd.n4554 gnd.n4480 19.3944
R7812 gnd.n4547 gnd.n4480 19.3944
R7813 gnd.n4547 gnd.n4546 19.3944
R7814 gnd.n4546 gnd.n4490 19.3944
R7815 gnd.n4539 gnd.n4490 19.3944
R7816 gnd.n4539 gnd.n4538 19.3944
R7817 gnd.n4538 gnd.n4500 19.3944
R7818 gnd.n4531 gnd.n4500 19.3944
R7819 gnd.n4531 gnd.n4530 19.3944
R7820 gnd.n4530 gnd.n4510 19.3944
R7821 gnd.n5801 gnd.n1510 19.3944
R7822 gnd.n5801 gnd.n5800 19.3944
R7823 gnd.n5800 gnd.n1513 19.3944
R7824 gnd.n5793 gnd.n1513 19.3944
R7825 gnd.n5793 gnd.n5792 19.3944
R7826 gnd.n5792 gnd.n1521 19.3944
R7827 gnd.n5785 gnd.n1521 19.3944
R7828 gnd.n5785 gnd.n5784 19.3944
R7829 gnd.n5784 gnd.n1529 19.3944
R7830 gnd.n5777 gnd.n1529 19.3944
R7831 gnd.n5777 gnd.n5776 19.3944
R7832 gnd.n5776 gnd.n1537 19.3944
R7833 gnd.n5769 gnd.n1537 19.3944
R7834 gnd.n5769 gnd.n5768 19.3944
R7835 gnd.n5768 gnd.n1545 19.3944
R7836 gnd.n5761 gnd.n1545 19.3944
R7837 gnd.n3049 gnd.n3048 19.3944
R7838 gnd.n3048 gnd.n3047 19.3944
R7839 gnd.n3047 gnd.n3046 19.3944
R7840 gnd.n3046 gnd.n3044 19.3944
R7841 gnd.n3044 gnd.n3041 19.3944
R7842 gnd.n3041 gnd.n3040 19.3944
R7843 gnd.n3040 gnd.n3037 19.3944
R7844 gnd.n3037 gnd.n3036 19.3944
R7845 gnd.n3036 gnd.n3033 19.3944
R7846 gnd.n3033 gnd.n3032 19.3944
R7847 gnd.n3032 gnd.n3029 19.3944
R7848 gnd.n3029 gnd.n3028 19.3944
R7849 gnd.n3028 gnd.n3025 19.3944
R7850 gnd.n3025 gnd.n3024 19.3944
R7851 gnd.n3024 gnd.n3021 19.3944
R7852 gnd.n3021 gnd.n3020 19.3944
R7853 gnd.n3020 gnd.n3017 19.3944
R7854 gnd.n3017 gnd.n3016 19.3944
R7855 gnd.n3016 gnd.n3013 19.3944
R7856 gnd.n3013 gnd.n3012 19.3944
R7857 gnd.n3012 gnd.n3009 19.3944
R7858 gnd.n3009 gnd.n3008 19.3944
R7859 gnd.n3005 gnd.n3004 19.3944
R7860 gnd.n3004 gnd.n2960 19.3944
R7861 gnd.n3055 gnd.n2960 19.3944
R7862 gnd.n3822 gnd.n3821 19.3944
R7863 gnd.n3821 gnd.n3818 19.3944
R7864 gnd.n3818 gnd.n3817 19.3944
R7865 gnd.n3867 gnd.n3866 19.3944
R7866 gnd.n3866 gnd.n3865 19.3944
R7867 gnd.n3865 gnd.n3862 19.3944
R7868 gnd.n3862 gnd.n3861 19.3944
R7869 gnd.n3861 gnd.n3858 19.3944
R7870 gnd.n3858 gnd.n3857 19.3944
R7871 gnd.n3857 gnd.n3854 19.3944
R7872 gnd.n3854 gnd.n3853 19.3944
R7873 gnd.n3853 gnd.n3850 19.3944
R7874 gnd.n3850 gnd.n3849 19.3944
R7875 gnd.n3849 gnd.n3846 19.3944
R7876 gnd.n3846 gnd.n3845 19.3944
R7877 gnd.n3845 gnd.n3842 19.3944
R7878 gnd.n3842 gnd.n3841 19.3944
R7879 gnd.n3841 gnd.n3838 19.3944
R7880 gnd.n3838 gnd.n3837 19.3944
R7881 gnd.n3837 gnd.n3834 19.3944
R7882 gnd.n3834 gnd.n3833 19.3944
R7883 gnd.n3833 gnd.n3830 19.3944
R7884 gnd.n3830 gnd.n3829 19.3944
R7885 gnd.n3829 gnd.n3826 19.3944
R7886 gnd.n3826 gnd.n3825 19.3944
R7887 gnd.n3148 gnd.n2857 19.3944
R7888 gnd.n3158 gnd.n2857 19.3944
R7889 gnd.n3159 gnd.n3158 19.3944
R7890 gnd.n3159 gnd.n2838 19.3944
R7891 gnd.n3179 gnd.n2838 19.3944
R7892 gnd.n3179 gnd.n2830 19.3944
R7893 gnd.n3189 gnd.n2830 19.3944
R7894 gnd.n3190 gnd.n3189 19.3944
R7895 gnd.n3191 gnd.n3190 19.3944
R7896 gnd.n3191 gnd.n2813 19.3944
R7897 gnd.n3208 gnd.n2813 19.3944
R7898 gnd.n3211 gnd.n3208 19.3944
R7899 gnd.n3211 gnd.n3210 19.3944
R7900 gnd.n3210 gnd.n2786 19.3944
R7901 gnd.n3250 gnd.n2786 19.3944
R7902 gnd.n3250 gnd.n2783 19.3944
R7903 gnd.n3256 gnd.n2783 19.3944
R7904 gnd.n3257 gnd.n3256 19.3944
R7905 gnd.n3257 gnd.n2781 19.3944
R7906 gnd.n3263 gnd.n2781 19.3944
R7907 gnd.n3266 gnd.n3263 19.3944
R7908 gnd.n3268 gnd.n3266 19.3944
R7909 gnd.n3274 gnd.n3268 19.3944
R7910 gnd.n3274 gnd.n3273 19.3944
R7911 gnd.n3273 gnd.n2656 19.3944
R7912 gnd.n3340 gnd.n2656 19.3944
R7913 gnd.n3341 gnd.n3340 19.3944
R7914 gnd.n3341 gnd.n2649 19.3944
R7915 gnd.n3352 gnd.n2649 19.3944
R7916 gnd.n3353 gnd.n3352 19.3944
R7917 gnd.n3353 gnd.n2632 19.3944
R7918 gnd.n2632 gnd.n2630 19.3944
R7919 gnd.n3377 gnd.n2630 19.3944
R7920 gnd.n3378 gnd.n3377 19.3944
R7921 gnd.n3378 gnd.n2601 19.3944
R7922 gnd.n3425 gnd.n2601 19.3944
R7923 gnd.n3426 gnd.n3425 19.3944
R7924 gnd.n3426 gnd.n2594 19.3944
R7925 gnd.n3437 gnd.n2594 19.3944
R7926 gnd.n3438 gnd.n3437 19.3944
R7927 gnd.n3438 gnd.n2577 19.3944
R7928 gnd.n2577 gnd.n2575 19.3944
R7929 gnd.n3462 gnd.n2575 19.3944
R7930 gnd.n3463 gnd.n3462 19.3944
R7931 gnd.n3463 gnd.n2547 19.3944
R7932 gnd.n3514 gnd.n2547 19.3944
R7933 gnd.n3515 gnd.n3514 19.3944
R7934 gnd.n3515 gnd.n2540 19.3944
R7935 gnd.n3783 gnd.n2540 19.3944
R7936 gnd.n3784 gnd.n3783 19.3944
R7937 gnd.n3784 gnd.n2521 19.3944
R7938 gnd.n3809 gnd.n2521 19.3944
R7939 gnd.n3809 gnd.n2522 19.3944
R7940 gnd.n3139 gnd.n3138 19.3944
R7941 gnd.n3138 gnd.n2871 19.3944
R7942 gnd.n2894 gnd.n2871 19.3944
R7943 gnd.n2897 gnd.n2894 19.3944
R7944 gnd.n2897 gnd.n2890 19.3944
R7945 gnd.n2901 gnd.n2890 19.3944
R7946 gnd.n2904 gnd.n2901 19.3944
R7947 gnd.n2907 gnd.n2904 19.3944
R7948 gnd.n2907 gnd.n2888 19.3944
R7949 gnd.n2911 gnd.n2888 19.3944
R7950 gnd.n2914 gnd.n2911 19.3944
R7951 gnd.n2917 gnd.n2914 19.3944
R7952 gnd.n2917 gnd.n2886 19.3944
R7953 gnd.n2921 gnd.n2886 19.3944
R7954 gnd.n3144 gnd.n3143 19.3944
R7955 gnd.n3143 gnd.n2847 19.3944
R7956 gnd.n3169 gnd.n2847 19.3944
R7957 gnd.n3169 gnd.n2845 19.3944
R7958 gnd.n3175 gnd.n2845 19.3944
R7959 gnd.n3175 gnd.n3174 19.3944
R7960 gnd.n3174 gnd.n2819 19.3944
R7961 gnd.n3199 gnd.n2819 19.3944
R7962 gnd.n3199 gnd.n2817 19.3944
R7963 gnd.n3203 gnd.n2817 19.3944
R7964 gnd.n3203 gnd.n2797 19.3944
R7965 gnd.n3230 gnd.n2797 19.3944
R7966 gnd.n3230 gnd.n2795 19.3944
R7967 gnd.n3240 gnd.n2795 19.3944
R7968 gnd.n3240 gnd.n3239 19.3944
R7969 gnd.n3239 gnd.n3238 19.3944
R7970 gnd.n3238 gnd.n2744 19.3944
R7971 gnd.n3288 gnd.n2744 19.3944
R7972 gnd.n3288 gnd.n3287 19.3944
R7973 gnd.n3287 gnd.n3286 19.3944
R7974 gnd.n3286 gnd.n2748 19.3944
R7975 gnd.n2768 gnd.n2748 19.3944
R7976 gnd.n2768 gnd.n2666 19.3944
R7977 gnd.n3325 gnd.n2666 19.3944
R7978 gnd.n3325 gnd.n2664 19.3944
R7979 gnd.n3331 gnd.n2664 19.3944
R7980 gnd.n3331 gnd.n3330 19.3944
R7981 gnd.n3330 gnd.n2639 19.3944
R7982 gnd.n3365 gnd.n2639 19.3944
R7983 gnd.n3365 gnd.n2637 19.3944
R7984 gnd.n3371 gnd.n2637 19.3944
R7985 gnd.n3371 gnd.n3370 19.3944
R7986 gnd.n3370 gnd.n2612 19.3944
R7987 gnd.n3410 gnd.n2612 19.3944
R7988 gnd.n3410 gnd.n2610 19.3944
R7989 gnd.n3416 gnd.n2610 19.3944
R7990 gnd.n3416 gnd.n3415 19.3944
R7991 gnd.n3415 gnd.n2584 19.3944
R7992 gnd.n3450 gnd.n2584 19.3944
R7993 gnd.n3450 gnd.n2582 19.3944
R7994 gnd.n3456 gnd.n2582 19.3944
R7995 gnd.n3456 gnd.n3455 19.3944
R7996 gnd.n3455 gnd.n2557 19.3944
R7997 gnd.n3499 gnd.n2557 19.3944
R7998 gnd.n3499 gnd.n2555 19.3944
R7999 gnd.n3505 gnd.n2555 19.3944
R8000 gnd.n3505 gnd.n3504 19.3944
R8001 gnd.n3504 gnd.n2530 19.3944
R8002 gnd.n3794 gnd.n2530 19.3944
R8003 gnd.n3794 gnd.n2528 19.3944
R8004 gnd.n3802 gnd.n2528 19.3944
R8005 gnd.n3802 gnd.n3801 19.3944
R8006 gnd.n3801 gnd.n3800 19.3944
R8007 gnd.n3903 gnd.n3902 19.3944
R8008 gnd.n3902 gnd.n2469 19.3944
R8009 gnd.n3898 gnd.n2469 19.3944
R8010 gnd.n3898 gnd.n3895 19.3944
R8011 gnd.n3895 gnd.n3892 19.3944
R8012 gnd.n3892 gnd.n3891 19.3944
R8013 gnd.n3891 gnd.n3888 19.3944
R8014 gnd.n3888 gnd.n3887 19.3944
R8015 gnd.n3887 gnd.n3884 19.3944
R8016 gnd.n3884 gnd.n3883 19.3944
R8017 gnd.n3883 gnd.n3880 19.3944
R8018 gnd.n3880 gnd.n3879 19.3944
R8019 gnd.n3879 gnd.n3876 19.3944
R8020 gnd.n3876 gnd.n3875 19.3944
R8021 gnd.n3059 gnd.n2958 19.3944
R8022 gnd.n3059 gnd.n2949 19.3944
R8023 gnd.n3072 gnd.n2949 19.3944
R8024 gnd.n3072 gnd.n2947 19.3944
R8025 gnd.n3076 gnd.n2947 19.3944
R8026 gnd.n3076 gnd.n2937 19.3944
R8027 gnd.n3088 gnd.n2937 19.3944
R8028 gnd.n3088 gnd.n2935 19.3944
R8029 gnd.n3122 gnd.n2935 19.3944
R8030 gnd.n3122 gnd.n3121 19.3944
R8031 gnd.n3121 gnd.n3120 19.3944
R8032 gnd.n3120 gnd.n3119 19.3944
R8033 gnd.n3119 gnd.n3116 19.3944
R8034 gnd.n3116 gnd.n3115 19.3944
R8035 gnd.n3115 gnd.n3114 19.3944
R8036 gnd.n3114 gnd.n3112 19.3944
R8037 gnd.n3112 gnd.n3111 19.3944
R8038 gnd.n3111 gnd.n3108 19.3944
R8039 gnd.n3108 gnd.n3107 19.3944
R8040 gnd.n3107 gnd.n3106 19.3944
R8041 gnd.n3106 gnd.n3104 19.3944
R8042 gnd.n3104 gnd.n2803 19.3944
R8043 gnd.n3219 gnd.n2803 19.3944
R8044 gnd.n3219 gnd.n2801 19.3944
R8045 gnd.n3225 gnd.n2801 19.3944
R8046 gnd.n3225 gnd.n3224 19.3944
R8047 gnd.n3224 gnd.n2725 19.3944
R8048 gnd.n3299 gnd.n2725 19.3944
R8049 gnd.n3299 gnd.n2726 19.3944
R8050 gnd.n2773 gnd.n2772 19.3944
R8051 gnd.n2776 gnd.n2775 19.3944
R8052 gnd.n2763 gnd.n2762 19.3944
R8053 gnd.n3318 gnd.n2671 19.3944
R8054 gnd.n3318 gnd.n3317 19.3944
R8055 gnd.n3317 gnd.n3316 19.3944
R8056 gnd.n3316 gnd.n3314 19.3944
R8057 gnd.n3314 gnd.n3313 19.3944
R8058 gnd.n3313 gnd.n3311 19.3944
R8059 gnd.n3311 gnd.n3310 19.3944
R8060 gnd.n3310 gnd.n2620 19.3944
R8061 gnd.n3386 gnd.n2620 19.3944
R8062 gnd.n3386 gnd.n2618 19.3944
R8063 gnd.n3405 gnd.n2618 19.3944
R8064 gnd.n3405 gnd.n3404 19.3944
R8065 gnd.n3404 gnd.n3403 19.3944
R8066 gnd.n3403 gnd.n3401 19.3944
R8067 gnd.n3401 gnd.n3400 19.3944
R8068 gnd.n3400 gnd.n3398 19.3944
R8069 gnd.n3398 gnd.n3397 19.3944
R8070 gnd.n3397 gnd.n2564 19.3944
R8071 gnd.n3471 gnd.n2564 19.3944
R8072 gnd.n3471 gnd.n2562 19.3944
R8073 gnd.n3494 gnd.n2562 19.3944
R8074 gnd.n3494 gnd.n3493 19.3944
R8075 gnd.n3493 gnd.n3492 19.3944
R8076 gnd.n3492 gnd.n3489 19.3944
R8077 gnd.n3489 gnd.n3488 19.3944
R8078 gnd.n3488 gnd.n3486 19.3944
R8079 gnd.n3486 gnd.n3485 19.3944
R8080 gnd.n3485 gnd.n3483 19.3944
R8081 gnd.n3483 gnd.n2516 19.3944
R8082 gnd.n3064 gnd.n2954 19.3944
R8083 gnd.n3064 gnd.n2952 19.3944
R8084 gnd.n3068 gnd.n2952 19.3944
R8085 gnd.n3068 gnd.n2943 19.3944
R8086 gnd.n3080 gnd.n2943 19.3944
R8087 gnd.n3080 gnd.n2941 19.3944
R8088 gnd.n3084 gnd.n2941 19.3944
R8089 gnd.n3084 gnd.n2930 19.3944
R8090 gnd.n3126 gnd.n2930 19.3944
R8091 gnd.n3126 gnd.n2884 19.3944
R8092 gnd.n3132 gnd.n2884 19.3944
R8093 gnd.n3132 gnd.n3131 19.3944
R8094 gnd.n3131 gnd.n2862 19.3944
R8095 gnd.n3153 gnd.n2862 19.3944
R8096 gnd.n3153 gnd.n2855 19.3944
R8097 gnd.n3164 gnd.n2855 19.3944
R8098 gnd.n3164 gnd.n3163 19.3944
R8099 gnd.n3163 gnd.n2836 19.3944
R8100 gnd.n3184 gnd.n2836 19.3944
R8101 gnd.n3184 gnd.n2826 19.3944
R8102 gnd.n3194 gnd.n2826 19.3944
R8103 gnd.n3194 gnd.n2809 19.3944
R8104 gnd.n3215 gnd.n2809 19.3944
R8105 gnd.n3215 gnd.n3214 19.3944
R8106 gnd.n3214 gnd.n2788 19.3944
R8107 gnd.n3245 gnd.n2788 19.3944
R8108 gnd.n3245 gnd.n2733 19.3944
R8109 gnd.n3295 gnd.n2733 19.3944
R8110 gnd.n3295 gnd.n3294 19.3944
R8111 gnd.n3294 gnd.n3293 19.3944
R8112 gnd.n3293 gnd.n2737 19.3944
R8113 gnd.n2755 gnd.n2737 19.3944
R8114 gnd.n3281 gnd.n2755 19.3944
R8115 gnd.n3281 gnd.n3280 19.3944
R8116 gnd.n3280 gnd.n3279 19.3944
R8117 gnd.n3279 gnd.n2759 19.3944
R8118 gnd.n2759 gnd.n2658 19.3944
R8119 gnd.n3336 gnd.n2658 19.3944
R8120 gnd.n3336 gnd.n2651 19.3944
R8121 gnd.n3347 gnd.n2651 19.3944
R8122 gnd.n3347 gnd.n2647 19.3944
R8123 gnd.n3360 gnd.n2647 19.3944
R8124 gnd.n3360 gnd.n3359 19.3944
R8125 gnd.n3359 gnd.n2626 19.3944
R8126 gnd.n3382 gnd.n2626 19.3944
R8127 gnd.n3382 gnd.n3381 19.3944
R8128 gnd.n3381 gnd.n2603 19.3944
R8129 gnd.n3421 gnd.n2603 19.3944
R8130 gnd.n3421 gnd.n2596 19.3944
R8131 gnd.n3432 gnd.n2596 19.3944
R8132 gnd.n3432 gnd.n2592 19.3944
R8133 gnd.n3445 gnd.n2592 19.3944
R8134 gnd.n3445 gnd.n3444 19.3944
R8135 gnd.n3444 gnd.n2571 19.3944
R8136 gnd.n3467 gnd.n2571 19.3944
R8137 gnd.n3467 gnd.n3466 19.3944
R8138 gnd.n3466 gnd.n2549 19.3944
R8139 gnd.n3510 gnd.n2549 19.3944
R8140 gnd.n3510 gnd.n2542 19.3944
R8141 gnd.n3522 gnd.n2542 19.3944
R8142 gnd.n3522 gnd.n2538 19.3944
R8143 gnd.n3789 gnd.n2538 19.3944
R8144 gnd.n3789 gnd.n3788 19.3944
R8145 gnd.n3788 gnd.n2519 19.3944
R8146 gnd.n3812 gnd.n2519 19.3944
R8147 gnd.n4567 gnd.n4566 19.3944
R8148 gnd.n4566 gnd.n4464 19.3944
R8149 gnd.n4559 gnd.n4464 19.3944
R8150 gnd.n4559 gnd.n4558 19.3944
R8151 gnd.n4558 gnd.n4476 19.3944
R8152 gnd.n4551 gnd.n4476 19.3944
R8153 gnd.n4551 gnd.n4550 19.3944
R8154 gnd.n4550 gnd.n4484 19.3944
R8155 gnd.n4543 gnd.n4484 19.3944
R8156 gnd.n4543 gnd.n4542 19.3944
R8157 gnd.n4542 gnd.n4496 19.3944
R8158 gnd.n4535 gnd.n4496 19.3944
R8159 gnd.n4535 gnd.n4534 19.3944
R8160 gnd.n4534 gnd.n4504 19.3944
R8161 gnd.n4527 gnd.n4504 19.3944
R8162 gnd.n4527 gnd.n4526 19.3944
R8163 gnd.n4403 gnd.n4401 19.3944
R8164 gnd.n4403 gnd.n4398 19.3944
R8165 gnd.n4407 gnd.n4398 19.3944
R8166 gnd.n4407 gnd.n2323 19.3944
R8167 gnd.n4411 gnd.n2323 19.3944
R8168 gnd.n4411 gnd.n2321 19.3944
R8169 gnd.n4419 gnd.n2321 19.3944
R8170 gnd.n4419 gnd.n4418 19.3944
R8171 gnd.n4418 gnd.n4417 19.3944
R8172 gnd.n4417 gnd.n2305 19.3944
R8173 gnd.n4694 gnd.n2305 19.3944
R8174 gnd.n4694 gnd.n2303 19.3944
R8175 gnd.n4698 gnd.n2303 19.3944
R8176 gnd.n4698 gnd.n2301 19.3944
R8177 gnd.n4702 gnd.n2301 19.3944
R8178 gnd.n4702 gnd.n2299 19.3944
R8179 gnd.n4711 gnd.n2299 19.3944
R8180 gnd.n4711 gnd.n4710 19.3944
R8181 gnd.n4710 gnd.n4709 19.3944
R8182 gnd.n4709 gnd.n2271 19.3944
R8183 gnd.n4740 gnd.n2271 19.3944
R8184 gnd.n4740 gnd.n2269 19.3944
R8185 gnd.n4753 gnd.n2269 19.3944
R8186 gnd.n4753 gnd.n4752 19.3944
R8187 gnd.n4752 gnd.n4751 19.3944
R8188 gnd.n4751 gnd.n4748 19.3944
R8189 gnd.n4748 gnd.n1284 19.3944
R8190 gnd.n5956 gnd.n1284 19.3944
R8191 gnd.n5956 gnd.n5955 19.3944
R8192 gnd.n5955 gnd.n5954 19.3944
R8193 gnd.n5954 gnd.n1288 19.3944
R8194 gnd.n1384 gnd.n1288 19.3944
R8195 gnd.n5937 gnd.n1384 19.3944
R8196 gnd.n5937 gnd.n5936 19.3944
R8197 gnd.n5936 gnd.n5935 19.3944
R8198 gnd.n5935 gnd.n1390 19.3944
R8199 gnd.n4839 gnd.n1390 19.3944
R8200 gnd.n4843 gnd.n4839 19.3944
R8201 gnd.n4843 gnd.n2227 19.3944
R8202 gnd.n4881 gnd.n2227 19.3944
R8203 gnd.n4881 gnd.n2225 19.3944
R8204 gnd.n4886 gnd.n2225 19.3944
R8205 gnd.n4886 gnd.n2195 19.3944
R8206 gnd.n4938 gnd.n2195 19.3944
R8207 gnd.n4938 gnd.n4937 19.3944
R8208 gnd.n4937 gnd.n4936 19.3944
R8209 gnd.n4936 gnd.n2199 19.3944
R8210 gnd.n2211 gnd.n2199 19.3944
R8211 gnd.n2211 gnd.n2210 19.3944
R8212 gnd.n2210 gnd.n2209 19.3944
R8213 gnd.n2209 gnd.n2206 19.3944
R8214 gnd.n2206 gnd.n2154 19.3944
R8215 gnd.n4996 gnd.n2154 19.3944
R8216 gnd.n4996 gnd.n2152 19.3944
R8217 gnd.n5002 gnd.n2152 19.3944
R8218 gnd.n5002 gnd.n5001 19.3944
R8219 gnd.n5001 gnd.n2128 19.3944
R8220 gnd.n5052 gnd.n2128 19.3944
R8221 gnd.n5052 gnd.n2126 19.3944
R8222 gnd.n5058 gnd.n2126 19.3944
R8223 gnd.n5058 gnd.n5057 19.3944
R8224 gnd.n5057 gnd.n2106 19.3944
R8225 gnd.n5099 gnd.n2106 19.3944
R8226 gnd.n5099 gnd.n2104 19.3944
R8227 gnd.n5103 gnd.n2104 19.3944
R8228 gnd.n5103 gnd.n2082 19.3944
R8229 gnd.n5129 gnd.n2082 19.3944
R8230 gnd.n5129 gnd.n2080 19.3944
R8231 gnd.n5133 gnd.n2080 19.3944
R8232 gnd.n5133 gnd.n2064 19.3944
R8233 gnd.n5177 gnd.n2064 19.3944
R8234 gnd.n5177 gnd.n2062 19.3944
R8235 gnd.n5183 gnd.n2062 19.3944
R8236 gnd.n5183 gnd.n5182 19.3944
R8237 gnd.n5182 gnd.n2038 19.3944
R8238 gnd.n5213 gnd.n2038 19.3944
R8239 gnd.n5213 gnd.n2036 19.3944
R8240 gnd.n5219 gnd.n2036 19.3944
R8241 gnd.n5219 gnd.n5218 19.3944
R8242 gnd.n5218 gnd.n2008 19.3944
R8243 gnd.n5277 gnd.n2008 19.3944
R8244 gnd.n5277 gnd.n2006 19.3944
R8245 gnd.n5281 gnd.n2006 19.3944
R8246 gnd.n5281 gnd.n1991 19.3944
R8247 gnd.n5306 gnd.n1991 19.3944
R8248 gnd.n5306 gnd.n1989 19.3944
R8249 gnd.n5312 gnd.n1989 19.3944
R8250 gnd.n5312 gnd.n5311 19.3944
R8251 gnd.n5311 gnd.n1965 19.3944
R8252 gnd.n5342 gnd.n1965 19.3944
R8253 gnd.n5342 gnd.n1963 19.3944
R8254 gnd.n5346 gnd.n1963 19.3944
R8255 gnd.n5346 gnd.n1937 19.3944
R8256 gnd.n5379 gnd.n1937 19.3944
R8257 gnd.n5379 gnd.n1935 19.3944
R8258 gnd.n5385 gnd.n1935 19.3944
R8259 gnd.n5385 gnd.n5384 19.3944
R8260 gnd.n5384 gnd.n1788 19.3944
R8261 gnd.n5487 gnd.n1788 19.3944
R8262 gnd.n5487 gnd.n1786 19.3944
R8263 gnd.n5494 gnd.n1786 19.3944
R8264 gnd.n5494 gnd.n5493 19.3944
R8265 gnd.n5493 gnd.n1777 19.3944
R8266 gnd.n5507 gnd.n1777 19.3944
R8267 gnd.n5508 gnd.n5507 19.3944
R8268 gnd.n5508 gnd.n1775 19.3944
R8269 gnd.n5526 gnd.n1775 19.3944
R8270 gnd.n5526 gnd.n5525 19.3944
R8271 gnd.n5525 gnd.n5524 19.3944
R8272 gnd.n5524 gnd.n5514 19.3944
R8273 gnd.n5520 gnd.n5514 19.3944
R8274 gnd.n5520 gnd.n5519 19.3944
R8275 gnd.n5519 gnd.n1743 19.3944
R8276 gnd.n1743 gnd.n1741 19.3944
R8277 gnd.n5577 gnd.n1741 19.3944
R8278 gnd.n5577 gnd.n1739 19.3944
R8279 gnd.n5581 gnd.n1739 19.3944
R8280 gnd.n5581 gnd.n1737 19.3944
R8281 gnd.n5585 gnd.n1737 19.3944
R8282 gnd.n5585 gnd.n1735 19.3944
R8283 gnd.n5598 gnd.n1735 19.3944
R8284 gnd.n5598 gnd.n5597 19.3944
R8285 gnd.n5597 gnd.n5596 19.3944
R8286 gnd.n5596 gnd.n5593 19.3944
R8287 gnd.n5593 gnd.n559 19.3944
R8288 gnd.n6854 gnd.n559 19.3944
R8289 gnd.n6854 gnd.n6853 19.3944
R8290 gnd.n6853 gnd.n6852 19.3944
R8291 gnd.n6636 gnd.n685 19.3944
R8292 gnd.n6642 gnd.n685 19.3944
R8293 gnd.n6642 gnd.n683 19.3944
R8294 gnd.n6646 gnd.n683 19.3944
R8295 gnd.n6646 gnd.n679 19.3944
R8296 gnd.n6652 gnd.n679 19.3944
R8297 gnd.n6652 gnd.n677 19.3944
R8298 gnd.n6656 gnd.n677 19.3944
R8299 gnd.n6656 gnd.n673 19.3944
R8300 gnd.n6662 gnd.n673 19.3944
R8301 gnd.n6662 gnd.n671 19.3944
R8302 gnd.n6666 gnd.n671 19.3944
R8303 gnd.n6666 gnd.n667 19.3944
R8304 gnd.n6672 gnd.n667 19.3944
R8305 gnd.n6672 gnd.n665 19.3944
R8306 gnd.n6676 gnd.n665 19.3944
R8307 gnd.n6676 gnd.n661 19.3944
R8308 gnd.n6682 gnd.n661 19.3944
R8309 gnd.n6682 gnd.n659 19.3944
R8310 gnd.n6686 gnd.n659 19.3944
R8311 gnd.n6686 gnd.n655 19.3944
R8312 gnd.n6692 gnd.n655 19.3944
R8313 gnd.n6692 gnd.n653 19.3944
R8314 gnd.n6696 gnd.n653 19.3944
R8315 gnd.n6696 gnd.n649 19.3944
R8316 gnd.n6702 gnd.n649 19.3944
R8317 gnd.n6702 gnd.n647 19.3944
R8318 gnd.n6706 gnd.n647 19.3944
R8319 gnd.n6706 gnd.n643 19.3944
R8320 gnd.n6712 gnd.n643 19.3944
R8321 gnd.n6712 gnd.n641 19.3944
R8322 gnd.n6716 gnd.n641 19.3944
R8323 gnd.n6716 gnd.n637 19.3944
R8324 gnd.n6722 gnd.n637 19.3944
R8325 gnd.n6722 gnd.n635 19.3944
R8326 gnd.n6726 gnd.n635 19.3944
R8327 gnd.n6726 gnd.n631 19.3944
R8328 gnd.n6732 gnd.n631 19.3944
R8329 gnd.n6732 gnd.n629 19.3944
R8330 gnd.n6736 gnd.n629 19.3944
R8331 gnd.n6736 gnd.n625 19.3944
R8332 gnd.n6742 gnd.n625 19.3944
R8333 gnd.n6742 gnd.n623 19.3944
R8334 gnd.n6746 gnd.n623 19.3944
R8335 gnd.n6746 gnd.n619 19.3944
R8336 gnd.n6752 gnd.n619 19.3944
R8337 gnd.n6752 gnd.n617 19.3944
R8338 gnd.n6756 gnd.n617 19.3944
R8339 gnd.n6756 gnd.n613 19.3944
R8340 gnd.n6762 gnd.n613 19.3944
R8341 gnd.n6762 gnd.n611 19.3944
R8342 gnd.n6766 gnd.n611 19.3944
R8343 gnd.n6766 gnd.n607 19.3944
R8344 gnd.n6772 gnd.n607 19.3944
R8345 gnd.n6772 gnd.n605 19.3944
R8346 gnd.n6776 gnd.n605 19.3944
R8347 gnd.n6776 gnd.n601 19.3944
R8348 gnd.n6782 gnd.n601 19.3944
R8349 gnd.n6782 gnd.n599 19.3944
R8350 gnd.n6786 gnd.n599 19.3944
R8351 gnd.n6786 gnd.n595 19.3944
R8352 gnd.n6792 gnd.n595 19.3944
R8353 gnd.n6792 gnd.n593 19.3944
R8354 gnd.n6796 gnd.n593 19.3944
R8355 gnd.n6796 gnd.n589 19.3944
R8356 gnd.n6802 gnd.n589 19.3944
R8357 gnd.n6802 gnd.n587 19.3944
R8358 gnd.n6806 gnd.n587 19.3944
R8359 gnd.n6806 gnd.n583 19.3944
R8360 gnd.n6812 gnd.n583 19.3944
R8361 gnd.n6812 gnd.n581 19.3944
R8362 gnd.n6816 gnd.n581 19.3944
R8363 gnd.n6816 gnd.n577 19.3944
R8364 gnd.n6822 gnd.n577 19.3944
R8365 gnd.n6822 gnd.n575 19.3944
R8366 gnd.n6826 gnd.n575 19.3944
R8367 gnd.n6826 gnd.n571 19.3944
R8368 gnd.n6832 gnd.n571 19.3944
R8369 gnd.n6832 gnd.n569 19.3944
R8370 gnd.n6836 gnd.n569 19.3944
R8371 gnd.n6836 gnd.n565 19.3944
R8372 gnd.n6843 gnd.n565 19.3944
R8373 gnd.n6843 gnd.n563 19.3944
R8374 gnd.n6847 gnd.n563 19.3944
R8375 gnd.n6315 gnd.n880 19.3944
R8376 gnd.n6315 gnd.n876 19.3944
R8377 gnd.n6321 gnd.n876 19.3944
R8378 gnd.n6321 gnd.n874 19.3944
R8379 gnd.n6325 gnd.n874 19.3944
R8380 gnd.n6325 gnd.n870 19.3944
R8381 gnd.n6331 gnd.n870 19.3944
R8382 gnd.n6331 gnd.n868 19.3944
R8383 gnd.n6335 gnd.n868 19.3944
R8384 gnd.n6335 gnd.n864 19.3944
R8385 gnd.n6341 gnd.n864 19.3944
R8386 gnd.n6341 gnd.n862 19.3944
R8387 gnd.n6345 gnd.n862 19.3944
R8388 gnd.n6345 gnd.n858 19.3944
R8389 gnd.n6351 gnd.n858 19.3944
R8390 gnd.n6351 gnd.n856 19.3944
R8391 gnd.n6355 gnd.n856 19.3944
R8392 gnd.n6355 gnd.n852 19.3944
R8393 gnd.n6361 gnd.n852 19.3944
R8394 gnd.n6361 gnd.n850 19.3944
R8395 gnd.n6365 gnd.n850 19.3944
R8396 gnd.n6365 gnd.n846 19.3944
R8397 gnd.n6371 gnd.n846 19.3944
R8398 gnd.n6371 gnd.n844 19.3944
R8399 gnd.n6375 gnd.n844 19.3944
R8400 gnd.n6375 gnd.n840 19.3944
R8401 gnd.n6381 gnd.n840 19.3944
R8402 gnd.n6381 gnd.n838 19.3944
R8403 gnd.n6385 gnd.n838 19.3944
R8404 gnd.n6385 gnd.n834 19.3944
R8405 gnd.n6391 gnd.n834 19.3944
R8406 gnd.n6391 gnd.n832 19.3944
R8407 gnd.n6395 gnd.n832 19.3944
R8408 gnd.n6395 gnd.n828 19.3944
R8409 gnd.n6401 gnd.n828 19.3944
R8410 gnd.n6401 gnd.n826 19.3944
R8411 gnd.n6405 gnd.n826 19.3944
R8412 gnd.n6405 gnd.n822 19.3944
R8413 gnd.n6411 gnd.n822 19.3944
R8414 gnd.n6411 gnd.n820 19.3944
R8415 gnd.n6415 gnd.n820 19.3944
R8416 gnd.n6415 gnd.n816 19.3944
R8417 gnd.n6421 gnd.n816 19.3944
R8418 gnd.n6421 gnd.n814 19.3944
R8419 gnd.n6425 gnd.n814 19.3944
R8420 gnd.n6425 gnd.n810 19.3944
R8421 gnd.n6431 gnd.n810 19.3944
R8422 gnd.n6431 gnd.n808 19.3944
R8423 gnd.n6435 gnd.n808 19.3944
R8424 gnd.n6435 gnd.n804 19.3944
R8425 gnd.n6441 gnd.n804 19.3944
R8426 gnd.n6441 gnd.n802 19.3944
R8427 gnd.n6445 gnd.n802 19.3944
R8428 gnd.n6445 gnd.n798 19.3944
R8429 gnd.n6451 gnd.n798 19.3944
R8430 gnd.n6451 gnd.n796 19.3944
R8431 gnd.n6455 gnd.n796 19.3944
R8432 gnd.n6455 gnd.n792 19.3944
R8433 gnd.n6461 gnd.n792 19.3944
R8434 gnd.n6461 gnd.n790 19.3944
R8435 gnd.n6465 gnd.n790 19.3944
R8436 gnd.n6465 gnd.n786 19.3944
R8437 gnd.n6471 gnd.n786 19.3944
R8438 gnd.n6471 gnd.n784 19.3944
R8439 gnd.n6475 gnd.n784 19.3944
R8440 gnd.n6475 gnd.n780 19.3944
R8441 gnd.n6481 gnd.n780 19.3944
R8442 gnd.n6481 gnd.n778 19.3944
R8443 gnd.n6485 gnd.n778 19.3944
R8444 gnd.n6485 gnd.n774 19.3944
R8445 gnd.n6491 gnd.n774 19.3944
R8446 gnd.n6491 gnd.n772 19.3944
R8447 gnd.n6495 gnd.n772 19.3944
R8448 gnd.n6495 gnd.n768 19.3944
R8449 gnd.n6501 gnd.n768 19.3944
R8450 gnd.n6501 gnd.n766 19.3944
R8451 gnd.n6505 gnd.n766 19.3944
R8452 gnd.n6505 gnd.n762 19.3944
R8453 gnd.n6511 gnd.n762 19.3944
R8454 gnd.n6511 gnd.n760 19.3944
R8455 gnd.n6515 gnd.n760 19.3944
R8456 gnd.n6515 gnd.n756 19.3944
R8457 gnd.n6521 gnd.n756 19.3944
R8458 gnd.n6521 gnd.n754 19.3944
R8459 gnd.n6525 gnd.n754 19.3944
R8460 gnd.n6525 gnd.n750 19.3944
R8461 gnd.n6531 gnd.n750 19.3944
R8462 gnd.n6531 gnd.n748 19.3944
R8463 gnd.n6535 gnd.n748 19.3944
R8464 gnd.n6535 gnd.n744 19.3944
R8465 gnd.n6541 gnd.n744 19.3944
R8466 gnd.n6541 gnd.n742 19.3944
R8467 gnd.n6545 gnd.n742 19.3944
R8468 gnd.n6545 gnd.n738 19.3944
R8469 gnd.n6551 gnd.n738 19.3944
R8470 gnd.n6551 gnd.n736 19.3944
R8471 gnd.n6555 gnd.n736 19.3944
R8472 gnd.n6555 gnd.n732 19.3944
R8473 gnd.n6561 gnd.n732 19.3944
R8474 gnd.n6561 gnd.n730 19.3944
R8475 gnd.n6565 gnd.n730 19.3944
R8476 gnd.n6565 gnd.n726 19.3944
R8477 gnd.n6571 gnd.n726 19.3944
R8478 gnd.n6571 gnd.n724 19.3944
R8479 gnd.n6575 gnd.n724 19.3944
R8480 gnd.n6575 gnd.n720 19.3944
R8481 gnd.n6581 gnd.n720 19.3944
R8482 gnd.n6581 gnd.n718 19.3944
R8483 gnd.n6585 gnd.n718 19.3944
R8484 gnd.n6585 gnd.n714 19.3944
R8485 gnd.n6591 gnd.n714 19.3944
R8486 gnd.n6591 gnd.n712 19.3944
R8487 gnd.n6595 gnd.n712 19.3944
R8488 gnd.n6595 gnd.n708 19.3944
R8489 gnd.n6601 gnd.n708 19.3944
R8490 gnd.n6601 gnd.n706 19.3944
R8491 gnd.n6605 gnd.n706 19.3944
R8492 gnd.n6605 gnd.n702 19.3944
R8493 gnd.n6611 gnd.n702 19.3944
R8494 gnd.n6611 gnd.n700 19.3944
R8495 gnd.n6615 gnd.n700 19.3944
R8496 gnd.n6615 gnd.n696 19.3944
R8497 gnd.n6621 gnd.n696 19.3944
R8498 gnd.n6621 gnd.n694 19.3944
R8499 gnd.n6626 gnd.n694 19.3944
R8500 gnd.n6626 gnd.n690 19.3944
R8501 gnd.n6632 gnd.n690 19.3944
R8502 gnd.n6633 gnd.n6632 19.3944
R8503 gnd.n5752 gnd.n5751 19.3944
R8504 gnd.n5751 gnd.n5750 19.3944
R8505 gnd.n5750 gnd.n5749 19.3944
R8506 gnd.n5749 gnd.n5747 19.3944
R8507 gnd.n5747 gnd.n5744 19.3944
R8508 gnd.n5744 gnd.n5743 19.3944
R8509 gnd.n5743 gnd.n5740 19.3944
R8510 gnd.n5740 gnd.n5739 19.3944
R8511 gnd.n5739 gnd.n5736 19.3944
R8512 gnd.n5736 gnd.n5735 19.3944
R8513 gnd.n5735 gnd.n5732 19.3944
R8514 gnd.n5732 gnd.n5731 19.3944
R8515 gnd.n5731 gnd.n5728 19.3944
R8516 gnd.n5728 gnd.n5727 19.3944
R8517 gnd.n5727 gnd.n5724 19.3944
R8518 gnd.n5724 gnd.n5723 19.3944
R8519 gnd.n5723 gnd.n5720 19.3944
R8520 gnd.n5718 gnd.n5715 19.3944
R8521 gnd.n5715 gnd.n5714 19.3944
R8522 gnd.n5714 gnd.n5711 19.3944
R8523 gnd.n5711 gnd.n5710 19.3944
R8524 gnd.n5710 gnd.n5707 19.3944
R8525 gnd.n5707 gnd.n5706 19.3944
R8526 gnd.n5706 gnd.n5703 19.3944
R8527 gnd.n5701 gnd.n5698 19.3944
R8528 gnd.n5698 gnd.n5697 19.3944
R8529 gnd.n5697 gnd.n5694 19.3944
R8530 gnd.n5694 gnd.n5693 19.3944
R8531 gnd.n5693 gnd.n5690 19.3944
R8532 gnd.n5690 gnd.n5689 19.3944
R8533 gnd.n5689 gnd.n5686 19.3944
R8534 gnd.n5686 gnd.n5685 19.3944
R8535 gnd.n5681 gnd.n5678 19.3944
R8536 gnd.n5678 gnd.n5677 19.3944
R8537 gnd.n5677 gnd.n5674 19.3944
R8538 gnd.n5674 gnd.n5673 19.3944
R8539 gnd.n5673 gnd.n5670 19.3944
R8540 gnd.n5670 gnd.n5669 19.3944
R8541 gnd.n5669 gnd.n5666 19.3944
R8542 gnd.n5666 gnd.n5665 19.3944
R8543 gnd.n5665 gnd.n5662 19.3944
R8544 gnd.n5662 gnd.n5661 19.3944
R8545 gnd.n5661 gnd.n5658 19.3944
R8546 gnd.n5658 gnd.n5657 19.3944
R8547 gnd.n5657 gnd.n5654 19.3944
R8548 gnd.n5654 gnd.n5653 19.3944
R8549 gnd.n5653 gnd.n5650 19.3944
R8550 gnd.n5650 gnd.n5649 19.3944
R8551 gnd.n5649 gnd.n5646 19.3944
R8552 gnd.n5646 gnd.n5645 19.3944
R8553 gnd.n5629 gnd.n1666 19.3944
R8554 gnd.n5629 gnd.n5628 19.3944
R8555 gnd.n5628 gnd.n1675 19.3944
R8556 gnd.n5542 gnd.n1675 19.3944
R8557 gnd.n5545 gnd.n5542 19.3944
R8558 gnd.n5546 gnd.n5545 19.3944
R8559 gnd.n5548 gnd.n5546 19.3944
R8560 gnd.n5548 gnd.n1723 19.3944
R8561 gnd.n5603 gnd.n1723 19.3944
R8562 gnd.n5603 gnd.n1729 19.3944
R8563 gnd.n1729 gnd.n1728 19.3944
R8564 gnd.n1728 gnd.n1727 19.3944
R8565 gnd.n1727 gnd.n1724 19.3944
R8566 gnd.n1724 gnd.n528 19.3944
R8567 gnd.n6885 gnd.n528 19.3944
R8568 gnd.n6886 gnd.n6885 19.3944
R8569 gnd.n6887 gnd.n6886 19.3944
R8570 gnd.n6890 gnd.n6887 19.3944
R8571 gnd.n6890 gnd.n6888 19.3944
R8572 gnd.n6888 gnd.n501 19.3944
R8573 gnd.n6923 gnd.n501 19.3944
R8574 gnd.n6925 gnd.n6923 19.3944
R8575 gnd.n6925 gnd.n6924 19.3944
R8576 gnd.n6924 gnd.n494 19.3944
R8577 gnd.n6937 gnd.n494 19.3944
R8578 gnd.n6938 gnd.n6937 19.3944
R8579 gnd.n6940 gnd.n6938 19.3944
R8580 gnd.n6941 gnd.n6940 19.3944
R8581 gnd.n6944 gnd.n6941 19.3944
R8582 gnd.n6945 gnd.n6944 19.3944
R8583 gnd.n6947 gnd.n6945 19.3944
R8584 gnd.n6948 gnd.n6947 19.3944
R8585 gnd.n6951 gnd.n6948 19.3944
R8586 gnd.n6952 gnd.n6951 19.3944
R8587 gnd.n6954 gnd.n6952 19.3944
R8588 gnd.n6955 gnd.n6954 19.3944
R8589 gnd.n6958 gnd.n6955 19.3944
R8590 gnd.n6959 gnd.n6958 19.3944
R8591 gnd.n6961 gnd.n6959 19.3944
R8592 gnd.n6962 gnd.n6961 19.3944
R8593 gnd.n6964 gnd.n6962 19.3944
R8594 gnd.n6965 gnd.n6964 19.3944
R8595 gnd.n5632 gnd.n5631 19.3944
R8596 gnd.n5631 gnd.n1673 19.3944
R8597 gnd.n1697 gnd.n1673 19.3944
R8598 gnd.n5618 gnd.n1697 19.3944
R8599 gnd.n5618 gnd.n5617 19.3944
R8600 gnd.n5617 gnd.n5616 19.3944
R8601 gnd.n5616 gnd.n1702 19.3944
R8602 gnd.n5606 gnd.n1702 19.3944
R8603 gnd.n5606 gnd.n5605 19.3944
R8604 gnd.n5605 gnd.n552 19.3944
R8605 gnd.n6862 gnd.n552 19.3944
R8606 gnd.n6862 gnd.n6861 19.3944
R8607 gnd.n6861 gnd.n6860 19.3944
R8608 gnd.n6860 gnd.n6859 19.3944
R8609 gnd.n6859 gnd.n525 19.3944
R8610 gnd.n6895 gnd.n525 19.3944
R8611 gnd.n6895 gnd.n6894 19.3944
R8612 gnd.n6894 gnd.n6893 19.3944
R8613 gnd.n6893 gnd.n503 19.3944
R8614 gnd.n6920 gnd.n503 19.3944
R8615 gnd.n6920 gnd.n496 19.3944
R8616 gnd.n6929 gnd.n496 19.3944
R8617 gnd.n6930 gnd.n6929 19.3944
R8618 gnd.n6932 gnd.n6930 19.3944
R8619 gnd.n6932 gnd.n91 19.3944
R8620 gnd.n7015 gnd.n91 19.3944
R8621 gnd.n7015 gnd.n7014 19.3944
R8622 gnd.n7014 gnd.n7013 19.3944
R8623 gnd.n7013 gnd.n95 19.3944
R8624 gnd.n7003 gnd.n95 19.3944
R8625 gnd.n7003 gnd.n7002 19.3944
R8626 gnd.n7002 gnd.n7001 19.3944
R8627 gnd.n7001 gnd.n112 19.3944
R8628 gnd.n6991 gnd.n112 19.3944
R8629 gnd.n6991 gnd.n6990 19.3944
R8630 gnd.n6990 gnd.n6989 19.3944
R8631 gnd.n6989 gnd.n132 19.3944
R8632 gnd.n6979 gnd.n132 19.3944
R8633 gnd.n6979 gnd.n6978 19.3944
R8634 gnd.n6978 gnd.n6977 19.3944
R8635 gnd.n6977 gnd.n152 19.3944
R8636 gnd.n6967 gnd.n152 19.3944
R8637 gnd.n442 gnd.n302 19.3944
R8638 gnd.n446 gnd.n302 19.3944
R8639 gnd.n446 gnd.n300 19.3944
R8640 gnd.n452 gnd.n300 19.3944
R8641 gnd.n452 gnd.n298 19.3944
R8642 gnd.n456 gnd.n298 19.3944
R8643 gnd.n456 gnd.n296 19.3944
R8644 gnd.n462 gnd.n296 19.3944
R8645 gnd.n462 gnd.n294 19.3944
R8646 gnd.n466 gnd.n294 19.3944
R8647 gnd.n466 gnd.n292 19.3944
R8648 gnd.n472 gnd.n292 19.3944
R8649 gnd.n472 gnd.n290 19.3944
R8650 gnd.n476 gnd.n290 19.3944
R8651 gnd.n476 gnd.n288 19.3944
R8652 gnd.n482 gnd.n288 19.3944
R8653 gnd.n482 gnd.n286 19.3944
R8654 gnd.n486 gnd.n286 19.3944
R8655 gnd.n392 gnd.n324 19.3944
R8656 gnd.n396 gnd.n324 19.3944
R8657 gnd.n396 gnd.n322 19.3944
R8658 gnd.n402 gnd.n322 19.3944
R8659 gnd.n402 gnd.n320 19.3944
R8660 gnd.n406 gnd.n320 19.3944
R8661 gnd.n406 gnd.n318 19.3944
R8662 gnd.n412 gnd.n318 19.3944
R8663 gnd.n412 gnd.n316 19.3944
R8664 gnd.n416 gnd.n316 19.3944
R8665 gnd.n416 gnd.n314 19.3944
R8666 gnd.n422 gnd.n314 19.3944
R8667 gnd.n422 gnd.n312 19.3944
R8668 gnd.n426 gnd.n312 19.3944
R8669 gnd.n426 gnd.n310 19.3944
R8670 gnd.n432 gnd.n310 19.3944
R8671 gnd.n432 gnd.n308 19.3944
R8672 gnd.n436 gnd.n308 19.3944
R8673 gnd.n346 gnd.n345 19.3944
R8674 gnd.n351 gnd.n346 19.3944
R8675 gnd.n351 gnd.n342 19.3944
R8676 gnd.n355 gnd.n342 19.3944
R8677 gnd.n355 gnd.n340 19.3944
R8678 gnd.n361 gnd.n340 19.3944
R8679 gnd.n361 gnd.n338 19.3944
R8680 gnd.n365 gnd.n338 19.3944
R8681 gnd.n365 gnd.n336 19.3944
R8682 gnd.n371 gnd.n336 19.3944
R8683 gnd.n371 gnd.n334 19.3944
R8684 gnd.n375 gnd.n334 19.3944
R8685 gnd.n375 gnd.n332 19.3944
R8686 gnd.n382 gnd.n332 19.3944
R8687 gnd.n382 gnd.n330 19.3944
R8688 gnd.n386 gnd.n330 19.3944
R8689 gnd.n387 gnd.n386 19.3944
R8690 gnd.n279 gnd.n278 19.3944
R8691 gnd.n278 gnd.n277 19.3944
R8692 gnd.n277 gnd.n171 19.3944
R8693 gnd.n272 gnd.n171 19.3944
R8694 gnd.n272 gnd.n271 19.3944
R8695 gnd.n271 gnd.n270 19.3944
R8696 gnd.n270 gnd.n178 19.3944
R8697 gnd.n265 gnd.n178 19.3944
R8698 gnd.n265 gnd.n264 19.3944
R8699 gnd.n264 gnd.n263 19.3944
R8700 gnd.n263 gnd.n185 19.3944
R8701 gnd.n258 gnd.n185 19.3944
R8702 gnd.n258 gnd.n257 19.3944
R8703 gnd.n257 gnd.n256 19.3944
R8704 gnd.n256 gnd.n192 19.3944
R8705 gnd.n251 gnd.n192 19.3944
R8706 gnd.n5570 gnd.n1744 19.3944
R8707 gnd.n5570 gnd.n1745 19.3944
R8708 gnd.n5566 gnd.n1745 19.3944
R8709 gnd.n5566 gnd.n5565 19.3944
R8710 gnd.n5565 gnd.n5564 19.3944
R8711 gnd.n5564 gnd.n5540 19.3944
R8712 gnd.n5560 gnd.n5540 19.3944
R8713 gnd.n5560 gnd.n5559 19.3944
R8714 gnd.n5559 gnd.n5558 19.3944
R8715 gnd.n5558 gnd.n5553 19.3944
R8716 gnd.n5554 gnd.n5553 19.3944
R8717 gnd.n5554 gnd.n534 19.3944
R8718 gnd.n6877 gnd.n534 19.3944
R8719 gnd.n6877 gnd.n532 19.3944
R8720 gnd.n6881 gnd.n532 19.3944
R8721 gnd.n6881 gnd.n515 19.3944
R8722 gnd.n6904 gnd.n515 19.3944
R8723 gnd.n6904 gnd.n512 19.3944
R8724 gnd.n6908 gnd.n512 19.3944
R8725 gnd.n6908 gnd.n513 19.3944
R8726 gnd.n513 gnd.n64 19.3944
R8727 gnd.n7028 gnd.n64 19.3944
R8728 gnd.n7028 gnd.n7027 19.3944
R8729 gnd.n7027 gnd.n67 19.3944
R8730 gnd.n217 gnd.n67 19.3944
R8731 gnd.n218 gnd.n217 19.3944
R8732 gnd.n218 gnd.n213 19.3944
R8733 gnd.n222 gnd.n213 19.3944
R8734 gnd.n224 gnd.n222 19.3944
R8735 gnd.n225 gnd.n224 19.3944
R8736 gnd.n225 gnd.n210 19.3944
R8737 gnd.n229 gnd.n210 19.3944
R8738 gnd.n231 gnd.n229 19.3944
R8739 gnd.n232 gnd.n231 19.3944
R8740 gnd.n232 gnd.n207 19.3944
R8741 gnd.n236 gnd.n207 19.3944
R8742 gnd.n238 gnd.n236 19.3944
R8743 gnd.n239 gnd.n238 19.3944
R8744 gnd.n239 gnd.n204 19.3944
R8745 gnd.n243 gnd.n204 19.3944
R8746 gnd.n245 gnd.n243 19.3944
R8747 gnd.n246 gnd.n245 19.3944
R8748 gnd.n1683 gnd.n1682 19.3944
R8749 gnd.n5624 gnd.n1682 19.3944
R8750 gnd.n5624 gnd.n5623 19.3944
R8751 gnd.n5623 gnd.n5622 19.3944
R8752 gnd.n5622 gnd.n1689 19.3944
R8753 gnd.n5612 gnd.n1689 19.3944
R8754 gnd.n5612 gnd.n5611 19.3944
R8755 gnd.n5611 gnd.n5610 19.3944
R8756 gnd.n5610 gnd.n1714 19.3944
R8757 gnd.n1714 gnd.n544 19.3944
R8758 gnd.n6866 gnd.n544 19.3944
R8759 gnd.n6866 gnd.n542 19.3944
R8760 gnd.n6873 gnd.n542 19.3944
R8761 gnd.n6873 gnd.n6872 19.3944
R8762 gnd.n6872 gnd.n6871 19.3944
R8763 gnd.n6871 gnd.n521 19.3944
R8764 gnd.n6900 gnd.n6899 19.3944
R8765 gnd.n6916 gnd.n6915 19.3944
R8766 gnd.n6913 gnd.n6912 19.3944
R8767 gnd.n7023 gnd.n7022 19.3944
R8768 gnd.n7019 gnd.n75 19.3944
R8769 gnd.n7019 gnd.n82 19.3944
R8770 gnd.n7009 gnd.n82 19.3944
R8771 gnd.n7009 gnd.n7008 19.3944
R8772 gnd.n7008 gnd.n7007 19.3944
R8773 gnd.n7007 gnd.n104 19.3944
R8774 gnd.n6997 gnd.n104 19.3944
R8775 gnd.n6997 gnd.n6996 19.3944
R8776 gnd.n6996 gnd.n6995 19.3944
R8777 gnd.n6995 gnd.n122 19.3944
R8778 gnd.n6985 gnd.n122 19.3944
R8779 gnd.n6985 gnd.n6984 19.3944
R8780 gnd.n6984 gnd.n6983 19.3944
R8781 gnd.n6983 gnd.n142 19.3944
R8782 gnd.n6973 gnd.n142 19.3944
R8783 gnd.n6973 gnd.n6972 19.3944
R8784 gnd.n6972 gnd.n6971 19.3944
R8785 gnd.n4238 gnd.n4237 19.3944
R8786 gnd.n4237 gnd.n4236 19.3944
R8787 gnd.n4236 gnd.n4235 19.3944
R8788 gnd.n4235 gnd.n4233 19.3944
R8789 gnd.n4233 gnd.n4230 19.3944
R8790 gnd.n4230 gnd.n4229 19.3944
R8791 gnd.n4229 gnd.n4226 19.3944
R8792 gnd.n4226 gnd.n4225 19.3944
R8793 gnd.n4225 gnd.n4222 19.3944
R8794 gnd.n4222 gnd.n4221 19.3944
R8795 gnd.n4221 gnd.n4218 19.3944
R8796 gnd.n4218 gnd.n4217 19.3944
R8797 gnd.n4217 gnd.n4214 19.3944
R8798 gnd.n4214 gnd.n4213 19.3944
R8799 gnd.n4213 gnd.n4210 19.3944
R8800 gnd.n4210 gnd.n4209 19.3944
R8801 gnd.n4209 gnd.n4206 19.3944
R8802 gnd.n4204 gnd.n4201 19.3944
R8803 gnd.n4201 gnd.n4200 19.3944
R8804 gnd.n4200 gnd.n4197 19.3944
R8805 gnd.n4197 gnd.n4196 19.3944
R8806 gnd.n4196 gnd.n4193 19.3944
R8807 gnd.n4193 gnd.n4192 19.3944
R8808 gnd.n4192 gnd.n4189 19.3944
R8809 gnd.n4189 gnd.n4188 19.3944
R8810 gnd.n4188 gnd.n4185 19.3944
R8811 gnd.n4185 gnd.n4184 19.3944
R8812 gnd.n4184 gnd.n4181 19.3944
R8813 gnd.n4181 gnd.n4180 19.3944
R8814 gnd.n4180 gnd.n4177 19.3944
R8815 gnd.n4177 gnd.n4176 19.3944
R8816 gnd.n4176 gnd.n4173 19.3944
R8817 gnd.n4173 gnd.n4172 19.3944
R8818 gnd.n4172 gnd.n4169 19.3944
R8819 gnd.n4169 gnd.n4168 19.3944
R8820 gnd.n4164 gnd.n4161 19.3944
R8821 gnd.n4161 gnd.n4160 19.3944
R8822 gnd.n4160 gnd.n4157 19.3944
R8823 gnd.n4157 gnd.n4156 19.3944
R8824 gnd.n4156 gnd.n4153 19.3944
R8825 gnd.n4153 gnd.n4152 19.3944
R8826 gnd.n4152 gnd.n4149 19.3944
R8827 gnd.n4149 gnd.n4148 19.3944
R8828 gnd.n4148 gnd.n4145 19.3944
R8829 gnd.n4145 gnd.n4144 19.3944
R8830 gnd.n4144 gnd.n4141 19.3944
R8831 gnd.n4141 gnd.n4140 19.3944
R8832 gnd.n4140 gnd.n4137 19.3944
R8833 gnd.n4137 gnd.n4136 19.3944
R8834 gnd.n4136 gnd.n4133 19.3944
R8835 gnd.n4133 gnd.n4132 19.3944
R8836 gnd.n4132 gnd.n4129 19.3944
R8837 gnd.n4129 gnd.n4128 19.3944
R8838 gnd.n4121 gnd.n4119 19.3944
R8839 gnd.n4119 gnd.n4116 19.3944
R8840 gnd.n4116 gnd.n4115 19.3944
R8841 gnd.n4115 gnd.n4112 19.3944
R8842 gnd.n4112 gnd.n4111 19.3944
R8843 gnd.n4111 gnd.n4108 19.3944
R8844 gnd.n4108 gnd.n4107 19.3944
R8845 gnd.n4107 gnd.n4104 19.3944
R8846 gnd.n4104 gnd.n4103 19.3944
R8847 gnd.n4103 gnd.n4100 19.3944
R8848 gnd.n4100 gnd.n4099 19.3944
R8849 gnd.n4099 gnd.n4096 19.3944
R8850 gnd.n4096 gnd.n4095 19.3944
R8851 gnd.n4095 gnd.n4092 19.3944
R8852 gnd.n4092 gnd.n4091 19.3944
R8853 gnd.n4091 gnd.n4088 19.3944
R8854 gnd.n4082 gnd.n4080 19.3944
R8855 gnd.n4080 gnd.n4079 19.3944
R8856 gnd.n4079 gnd.n4077 19.3944
R8857 gnd.n4077 gnd.n4076 19.3944
R8858 gnd.n4076 gnd.n4074 19.3944
R8859 gnd.n4074 gnd.n4073 19.3944
R8860 gnd.n4073 gnd.n4071 19.3944
R8861 gnd.n4071 gnd.n4070 19.3944
R8862 gnd.n4070 gnd.n4068 19.3944
R8863 gnd.n4068 gnd.n4067 19.3944
R8864 gnd.n4067 gnd.n4065 19.3944
R8865 gnd.n4065 gnd.n4064 19.3944
R8866 gnd.n4064 gnd.n4062 19.3944
R8867 gnd.n4062 gnd.n4061 19.3944
R8868 gnd.n4061 gnd.n4059 19.3944
R8869 gnd.n4059 gnd.n4058 19.3944
R8870 gnd.n4058 gnd.n4056 19.3944
R8871 gnd.n4056 gnd.n4055 19.3944
R8872 gnd.n4055 gnd.n4053 19.3944
R8873 gnd.n4053 gnd.n4052 19.3944
R8874 gnd.n4052 gnd.n4050 19.3944
R8875 gnd.n4050 gnd.n4047 19.3944
R8876 gnd.n4047 gnd.n2332 19.3944
R8877 gnd.n4370 gnd.n2332 19.3944
R8878 gnd.n4370 gnd.n2330 19.3944
R8879 gnd.n4374 gnd.n2330 19.3944
R8880 gnd.n4374 gnd.n2325 19.3944
R8881 gnd.n4393 gnd.n2325 19.3944
R8882 gnd.n4393 gnd.n2326 19.3944
R8883 gnd.n4389 gnd.n2326 19.3944
R8884 gnd.n4389 gnd.n2317 19.3944
R8885 gnd.n4424 gnd.n2317 19.3944
R8886 gnd.n4424 gnd.n2315 19.3944
R8887 gnd.n4428 gnd.n2315 19.3944
R8888 gnd.n4428 gnd.n2308 19.3944
R8889 gnd.n4688 gnd.n2308 19.3944
R8890 gnd.n4688 gnd.n2309 19.3944
R8891 gnd.n4684 gnd.n2309 19.3944
R8892 gnd.n4684 gnd.n4683 19.3944
R8893 gnd.n4683 gnd.n4682 19.3944
R8894 gnd.n4682 gnd.n4679 19.3944
R8895 gnd.n4679 gnd.n2295 19.3944
R8896 gnd.n4247 gnd.n4245 19.3944
R8897 gnd.n4247 gnd.n4246 19.3944
R8898 gnd.n4246 gnd.n2419 19.3944
R8899 gnd.n4262 gnd.n2419 19.3944
R8900 gnd.n4263 gnd.n4262 19.3944
R8901 gnd.n4264 gnd.n4263 19.3944
R8902 gnd.n4264 gnd.n2401 19.3944
R8903 gnd.n4282 gnd.n2401 19.3944
R8904 gnd.n4283 gnd.n4282 19.3944
R8905 gnd.n4284 gnd.n4283 19.3944
R8906 gnd.n4284 gnd.n2383 19.3944
R8907 gnd.n4302 gnd.n2383 19.3944
R8908 gnd.n4303 gnd.n4302 19.3944
R8909 gnd.n4304 gnd.n4303 19.3944
R8910 gnd.n4304 gnd.n2365 19.3944
R8911 gnd.n4323 gnd.n2365 19.3944
R8912 gnd.n4324 gnd.n4323 19.3944
R8913 gnd.n4325 gnd.n4324 19.3944
R8914 gnd.n4325 gnd.n2349 19.3944
R8915 gnd.n4343 gnd.n2349 19.3944
R8916 gnd.n4344 gnd.n4343 19.3944
R8917 gnd.n4346 gnd.n4344 19.3944
R8918 gnd.n4347 gnd.n4346 19.3944
R8919 gnd.n4349 gnd.n4347 19.3944
R8920 gnd.n4349 gnd.n2328 19.3944
R8921 gnd.n4378 gnd.n2328 19.3944
R8922 gnd.n4379 gnd.n4378 19.3944
R8923 gnd.n4380 gnd.n4379 19.3944
R8924 gnd.n4381 gnd.n4380 19.3944
R8925 gnd.n4385 gnd.n4381 19.3944
R8926 gnd.n4385 gnd.n4384 19.3944
R8927 gnd.n4384 gnd.n4383 19.3944
R8928 gnd.n4383 gnd.n2313 19.3944
R8929 gnd.n4432 gnd.n2313 19.3944
R8930 gnd.n4433 gnd.n4432 19.3944
R8931 gnd.n4434 gnd.n4433 19.3944
R8932 gnd.n4435 gnd.n4434 19.3944
R8933 gnd.n4439 gnd.n4435 19.3944
R8934 gnd.n4440 gnd.n4439 19.3944
R8935 gnd.n4675 gnd.n4440 19.3944
R8936 gnd.n4675 gnd.n4674 19.3944
R8937 gnd.n4674 gnd.n4673 19.3944
R8938 gnd.n4249 gnd.n2435 19.3944
R8939 gnd.n4249 gnd.n2436 19.3944
R8940 gnd.n2438 gnd.n2436 19.3944
R8941 gnd.n2438 gnd.n2417 19.3944
R8942 gnd.n4269 gnd.n2417 19.3944
R8943 gnd.n4269 gnd.n4268 19.3944
R8944 gnd.n4268 gnd.n4267 19.3944
R8945 gnd.n4267 gnd.n2399 19.3944
R8946 gnd.n4289 gnd.n2399 19.3944
R8947 gnd.n4289 gnd.n4288 19.3944
R8948 gnd.n4288 gnd.n4287 19.3944
R8949 gnd.n4287 gnd.n2381 19.3944
R8950 gnd.n4309 gnd.n2381 19.3944
R8951 gnd.n4309 gnd.n4308 19.3944
R8952 gnd.n4308 gnd.n4307 19.3944
R8953 gnd.n4307 gnd.n2363 19.3944
R8954 gnd.n4330 gnd.n2363 19.3944
R8955 gnd.n4330 gnd.n4329 19.3944
R8956 gnd.n4329 gnd.n4328 19.3944
R8957 gnd.n4328 gnd.n2345 19.3944
R8958 gnd.n4357 gnd.n2345 19.3944
R8959 gnd.n4357 gnd.n4356 19.3944
R8960 gnd.n4356 gnd.n4355 19.3944
R8961 gnd.n4355 gnd.n4354 19.3944
R8962 gnd.n4354 gnd.n4352 19.3944
R8963 gnd.n4352 gnd.n1067 19.3944
R8964 gnd.n6132 gnd.n1067 19.3944
R8965 gnd.n6132 gnd.n6131 19.3944
R8966 gnd.n6131 gnd.n6130 19.3944
R8967 gnd.n6130 gnd.n1071 19.3944
R8968 gnd.n6120 gnd.n1071 19.3944
R8969 gnd.n6120 gnd.n6119 19.3944
R8970 gnd.n6119 gnd.n6118 19.3944
R8971 gnd.n6118 gnd.n1092 19.3944
R8972 gnd.n6108 gnd.n1092 19.3944
R8973 gnd.n6108 gnd.n6107 19.3944
R8974 gnd.n6107 gnd.n6106 19.3944
R8975 gnd.n6106 gnd.n1111 19.3944
R8976 gnd.n6096 gnd.n1111 19.3944
R8977 gnd.n6096 gnd.n6095 19.3944
R8978 gnd.n6095 gnd.n6094 19.3944
R8979 gnd.n6094 gnd.n1132 19.3944
R8980 gnd.n6086 gnd.n1142 19.3944
R8981 gnd.n6081 gnd.n1142 19.3944
R8982 gnd.n6081 gnd.n6080 19.3944
R8983 gnd.n6080 gnd.n6079 19.3944
R8984 gnd.n6079 gnd.n6076 19.3944
R8985 gnd.n6076 gnd.n6075 19.3944
R8986 gnd.n6075 gnd.n6072 19.3944
R8987 gnd.n6072 gnd.n6071 19.3944
R8988 gnd.n6071 gnd.n6068 19.3944
R8989 gnd.n6068 gnd.n6067 19.3944
R8990 gnd.n6067 gnd.n6064 19.3944
R8991 gnd.n6064 gnd.n6063 19.3944
R8992 gnd.n6063 gnd.n6060 19.3944
R8993 gnd.n6060 gnd.n6059 19.3944
R8994 gnd.n6059 gnd.n6056 19.3944
R8995 gnd.n6056 gnd.n6055 19.3944
R8996 gnd.n6055 gnd.n6052 19.3944
R8997 gnd.n4621 gnd.n4587 19.3944
R8998 gnd.n4625 gnd.n4587 19.3944
R8999 gnd.n4628 gnd.n4625 19.3944
R9000 gnd.n4631 gnd.n4628 19.3944
R9001 gnd.n4631 gnd.n4585 19.3944
R9002 gnd.n4635 gnd.n4585 19.3944
R9003 gnd.n4638 gnd.n4635 19.3944
R9004 gnd.n4641 gnd.n4638 19.3944
R9005 gnd.n4641 gnd.n4583 19.3944
R9006 gnd.n4645 gnd.n4583 19.3944
R9007 gnd.n4648 gnd.n4645 19.3944
R9008 gnd.n4651 gnd.n4648 19.3944
R9009 gnd.n4651 gnd.n4581 19.3944
R9010 gnd.n4655 gnd.n4581 19.3944
R9011 gnd.n4658 gnd.n4655 19.3944
R9012 gnd.n4661 gnd.n4658 19.3944
R9013 gnd.n4661 gnd.n4579 19.3944
R9014 gnd.n4666 gnd.n4579 19.3944
R9015 gnd.n4599 gnd.n1211 19.3944
R9016 gnd.n4602 gnd.n4599 19.3944
R9017 gnd.n4602 gnd.n4594 19.3944
R9018 gnd.n4606 gnd.n4594 19.3944
R9019 gnd.n4609 gnd.n4606 19.3944
R9020 gnd.n4612 gnd.n4609 19.3944
R9021 gnd.n4612 gnd.n4592 19.3944
R9022 gnd.n4617 gnd.n4592 19.3944
R9023 gnd.n6050 gnd.n6047 19.3944
R9024 gnd.n6047 gnd.n6046 19.3944
R9025 gnd.n6046 gnd.n6043 19.3944
R9026 gnd.n6043 gnd.n6042 19.3944
R9027 gnd.n6042 gnd.n6039 19.3944
R9028 gnd.n6039 gnd.n6038 19.3944
R9029 gnd.n6038 gnd.n6035 19.3944
R9030 gnd.n4253 gnd.n2428 19.3944
R9031 gnd.n4253 gnd.n2426 19.3944
R9032 gnd.n4257 gnd.n2426 19.3944
R9033 gnd.n4257 gnd.n2409 19.3944
R9034 gnd.n4273 gnd.n2409 19.3944
R9035 gnd.n4273 gnd.n2407 19.3944
R9036 gnd.n4277 gnd.n2407 19.3944
R9037 gnd.n4277 gnd.n2392 19.3944
R9038 gnd.n4293 gnd.n2392 19.3944
R9039 gnd.n4293 gnd.n2390 19.3944
R9040 gnd.n4297 gnd.n2390 19.3944
R9041 gnd.n4297 gnd.n2373 19.3944
R9042 gnd.n4313 gnd.n2373 19.3944
R9043 gnd.n4313 gnd.n2371 19.3944
R9044 gnd.n4318 gnd.n2371 19.3944
R9045 gnd.n4318 gnd.n4317 19.3944
R9046 gnd.n4335 gnd.n4334 19.3944
R9047 gnd.n4338 gnd.n4337 19.3944
R9048 gnd.n4362 gnd.n4361 19.3944
R9049 gnd.n4365 gnd.n4364 19.3944
R9050 gnd.n6138 gnd.n6137 19.3944
R9051 gnd.n6137 gnd.n6136 19.3944
R9052 gnd.n6136 gnd.n1060 19.3944
R9053 gnd.n6126 gnd.n1060 19.3944
R9054 gnd.n6126 gnd.n6125 19.3944
R9055 gnd.n6125 gnd.n6124 19.3944
R9056 gnd.n6124 gnd.n1082 19.3944
R9057 gnd.n6114 gnd.n1082 19.3944
R9058 gnd.n6114 gnd.n6113 19.3944
R9059 gnd.n6113 gnd.n6112 19.3944
R9060 gnd.n6112 gnd.n1102 19.3944
R9061 gnd.n6102 gnd.n1102 19.3944
R9062 gnd.n6102 gnd.n6101 19.3944
R9063 gnd.n6101 gnd.n6100 19.3944
R9064 gnd.n6100 gnd.n1122 19.3944
R9065 gnd.n6090 gnd.n1122 19.3944
R9066 gnd.n6090 gnd.n6089 19.3944
R9067 gnd.n6311 gnd.n882 19.3944
R9068 gnd.n6305 gnd.n882 19.3944
R9069 gnd.n6305 gnd.n6304 19.3944
R9070 gnd.n6304 gnd.n6303 19.3944
R9071 gnd.n6303 gnd.n889 19.3944
R9072 gnd.n6297 gnd.n889 19.3944
R9073 gnd.n6297 gnd.n6296 19.3944
R9074 gnd.n6296 gnd.n6295 19.3944
R9075 gnd.n6295 gnd.n897 19.3944
R9076 gnd.n6289 gnd.n897 19.3944
R9077 gnd.n6289 gnd.n6288 19.3944
R9078 gnd.n6288 gnd.n6287 19.3944
R9079 gnd.n6287 gnd.n905 19.3944
R9080 gnd.n6281 gnd.n905 19.3944
R9081 gnd.n6281 gnd.n6280 19.3944
R9082 gnd.n6280 gnd.n6279 19.3944
R9083 gnd.n6279 gnd.n913 19.3944
R9084 gnd.n6273 gnd.n913 19.3944
R9085 gnd.n6273 gnd.n6272 19.3944
R9086 gnd.n6272 gnd.n6271 19.3944
R9087 gnd.n6271 gnd.n921 19.3944
R9088 gnd.n6265 gnd.n921 19.3944
R9089 gnd.n6265 gnd.n6264 19.3944
R9090 gnd.n6264 gnd.n6263 19.3944
R9091 gnd.n6263 gnd.n929 19.3944
R9092 gnd.n6257 gnd.n929 19.3944
R9093 gnd.n6257 gnd.n6256 19.3944
R9094 gnd.n6256 gnd.n6255 19.3944
R9095 gnd.n6255 gnd.n937 19.3944
R9096 gnd.n6249 gnd.n937 19.3944
R9097 gnd.n6249 gnd.n6248 19.3944
R9098 gnd.n6248 gnd.n6247 19.3944
R9099 gnd.n6247 gnd.n945 19.3944
R9100 gnd.n6241 gnd.n945 19.3944
R9101 gnd.n6241 gnd.n6240 19.3944
R9102 gnd.n6240 gnd.n6239 19.3944
R9103 gnd.n6239 gnd.n953 19.3944
R9104 gnd.n6233 gnd.n953 19.3944
R9105 gnd.n6233 gnd.n6232 19.3944
R9106 gnd.n6232 gnd.n6231 19.3944
R9107 gnd.n6231 gnd.n961 19.3944
R9108 gnd.n6225 gnd.n961 19.3944
R9109 gnd.n6225 gnd.n6224 19.3944
R9110 gnd.n6224 gnd.n6223 19.3944
R9111 gnd.n6223 gnd.n969 19.3944
R9112 gnd.n6217 gnd.n969 19.3944
R9113 gnd.n6217 gnd.n6216 19.3944
R9114 gnd.n6216 gnd.n6215 19.3944
R9115 gnd.n6215 gnd.n977 19.3944
R9116 gnd.n6209 gnd.n977 19.3944
R9117 gnd.n6209 gnd.n6208 19.3944
R9118 gnd.n6208 gnd.n6207 19.3944
R9119 gnd.n6207 gnd.n985 19.3944
R9120 gnd.n6201 gnd.n985 19.3944
R9121 gnd.n6201 gnd.n6200 19.3944
R9122 gnd.n6200 gnd.n6199 19.3944
R9123 gnd.n6199 gnd.n993 19.3944
R9124 gnd.n6193 gnd.n993 19.3944
R9125 gnd.n6193 gnd.n6192 19.3944
R9126 gnd.n6192 gnd.n6191 19.3944
R9127 gnd.n6191 gnd.n1001 19.3944
R9128 gnd.n6185 gnd.n1001 19.3944
R9129 gnd.n6185 gnd.n6184 19.3944
R9130 gnd.n6184 gnd.n6183 19.3944
R9131 gnd.n6183 gnd.n1009 19.3944
R9132 gnd.n6177 gnd.n1009 19.3944
R9133 gnd.n6177 gnd.n6176 19.3944
R9134 gnd.n6176 gnd.n6175 19.3944
R9135 gnd.n6175 gnd.n1017 19.3944
R9136 gnd.n6169 gnd.n1017 19.3944
R9137 gnd.n6169 gnd.n6168 19.3944
R9138 gnd.n6168 gnd.n6167 19.3944
R9139 gnd.n6167 gnd.n1025 19.3944
R9140 gnd.n6161 gnd.n1025 19.3944
R9141 gnd.n6161 gnd.n6160 19.3944
R9142 gnd.n6160 gnd.n6159 19.3944
R9143 gnd.n6159 gnd.n1033 19.3944
R9144 gnd.n6153 gnd.n1033 19.3944
R9145 gnd.n6153 gnd.n6152 19.3944
R9146 gnd.n6152 gnd.n6151 19.3944
R9147 gnd.n6151 gnd.n1041 19.3944
R9148 gnd.n6145 gnd.n1041 19.3944
R9149 gnd.n6145 gnd.n6144 19.3944
R9150 gnd.n6144 gnd.n6143 19.3944
R9151 gnd.n4757 gnd.n2261 19.3944
R9152 gnd.n4761 gnd.n2261 19.3944
R9153 gnd.n4761 gnd.n2259 19.3944
R9154 gnd.n4765 gnd.n2259 19.3944
R9155 gnd.n4765 gnd.n2257 19.3944
R9156 gnd.n4769 gnd.n2257 19.3944
R9157 gnd.n4769 gnd.n2250 19.3944
R9158 gnd.n4790 gnd.n2250 19.3944
R9159 gnd.n4790 gnd.n2248 19.3944
R9160 gnd.n4794 gnd.n2248 19.3944
R9161 gnd.n4825 gnd.n4794 19.3944
R9162 gnd.n4826 gnd.n4825 19.3944
R9163 gnd.n4826 gnd.n2245 19.3944
R9164 gnd.n4835 gnd.n2245 19.3944
R9165 gnd.n4835 gnd.n2246 19.3944
R9166 gnd.n4831 gnd.n2246 19.3944
R9167 gnd.n4831 gnd.n4830 19.3944
R9168 gnd.n4830 gnd.n2219 19.3944
R9169 gnd.n4889 gnd.n2219 19.3944
R9170 gnd.n4889 gnd.n2217 19.3944
R9171 gnd.n4893 gnd.n2217 19.3944
R9172 gnd.n4894 gnd.n4893 19.3944
R9173 gnd.n4897 gnd.n4894 19.3944
R9174 gnd.n4897 gnd.n2214 19.3944
R9175 gnd.n4928 gnd.n2214 19.3944
R9176 gnd.n4928 gnd.n2215 19.3944
R9177 gnd.n4924 gnd.n2215 19.3944
R9178 gnd.n4924 gnd.n4923 19.3944
R9179 gnd.n4923 gnd.n4922 19.3944
R9180 gnd.n4922 gnd.n4903 19.3944
R9181 gnd.n4918 gnd.n4903 19.3944
R9182 gnd.n4918 gnd.n4917 19.3944
R9183 gnd.n4917 gnd.n4916 19.3944
R9184 gnd.n4916 gnd.n4911 19.3944
R9185 gnd.n4912 gnd.n4911 19.3944
R9186 gnd.n4912 gnd.n2119 19.3944
R9187 gnd.n5062 gnd.n2119 19.3944
R9188 gnd.n5062 gnd.n2116 19.3944
R9189 gnd.n5087 gnd.n2116 19.3944
R9190 gnd.n5087 gnd.n2117 19.3944
R9191 gnd.n5083 gnd.n2117 19.3944
R9192 gnd.n5083 gnd.n5082 19.3944
R9193 gnd.n5082 gnd.n5081 19.3944
R9194 gnd.n5081 gnd.n5068 19.3944
R9195 gnd.n5077 gnd.n5068 19.3944
R9196 gnd.n5077 gnd.n5076 19.3944
R9197 gnd.n5076 gnd.n5075 19.3944
R9198 gnd.n5075 gnd.n5072 19.3944
R9199 gnd.n5072 gnd.n2055 19.3944
R9200 gnd.n5187 gnd.n2055 19.3944
R9201 gnd.n5187 gnd.n2052 19.3944
R9202 gnd.n5195 gnd.n2052 19.3944
R9203 gnd.n5195 gnd.n2053 19.3944
R9204 gnd.n5191 gnd.n2053 19.3944
R9205 gnd.n5191 gnd.n2030 19.3944
R9206 gnd.n2030 gnd.n2028 19.3944
R9207 gnd.n5225 gnd.n2028 19.3944
R9208 gnd.n5225 gnd.n2025 19.3944
R9209 gnd.n5258 gnd.n2025 19.3944
R9210 gnd.n5258 gnd.n2026 19.3944
R9211 gnd.n5254 gnd.n2026 19.3944
R9212 gnd.n5254 gnd.n5253 19.3944
R9213 gnd.n5253 gnd.n5252 19.3944
R9214 gnd.n5252 gnd.n5230 19.3944
R9215 gnd.n5248 gnd.n5230 19.3944
R9216 gnd.n5248 gnd.n5247 19.3944
R9217 gnd.n5247 gnd.n5246 19.3944
R9218 gnd.n5246 gnd.n5236 19.3944
R9219 gnd.n5242 gnd.n5236 19.3944
R9220 gnd.n5242 gnd.n5241 19.3944
R9221 gnd.n5241 gnd.n5240 19.3944
R9222 gnd.n5240 gnd.n1929 19.3944
R9223 gnd.n5389 gnd.n1929 19.3944
R9224 gnd.n5389 gnd.n1926 19.3944
R9225 gnd.n5394 gnd.n1926 19.3944
R9226 gnd.n5394 gnd.n1927 19.3944
R9227 gnd.n1927 gnd.n1782 19.3944
R9228 gnd.n5498 gnd.n1782 19.3944
R9229 gnd.n5498 gnd.n1780 19.3944
R9230 gnd.n5502 gnd.n1780 19.3944
R9231 gnd.n5502 gnd.n1493 19.3944
R9232 gnd.n5821 gnd.n1493 19.3944
R9233 gnd.n5818 gnd.n5817 19.3944
R9234 gnd.n5817 gnd.n5816 19.3944
R9235 gnd.n5816 gnd.n1498 19.3944
R9236 gnd.n5812 gnd.n1498 19.3944
R9237 gnd.n5812 gnd.n5811 19.3944
R9238 gnd.n5811 gnd.n5810 19.3944
R9239 gnd.n5810 gnd.n1503 19.3944
R9240 gnd.n5805 gnd.n1503 19.3944
R9241 gnd.n5805 gnd.n5804 19.3944
R9242 gnd.n5804 gnd.n1508 19.3944
R9243 gnd.n5797 gnd.n1508 19.3944
R9244 gnd.n5797 gnd.n5796 19.3944
R9245 gnd.n5796 gnd.n1517 19.3944
R9246 gnd.n5789 gnd.n1517 19.3944
R9247 gnd.n5789 gnd.n5788 19.3944
R9248 gnd.n5788 gnd.n1525 19.3944
R9249 gnd.n5781 gnd.n1525 19.3944
R9250 gnd.n5781 gnd.n5780 19.3944
R9251 gnd.n5780 gnd.n1533 19.3944
R9252 gnd.n5773 gnd.n1533 19.3944
R9253 gnd.n5773 gnd.n5772 19.3944
R9254 gnd.n5772 gnd.n1541 19.3944
R9255 gnd.n5765 gnd.n1541 19.3944
R9256 gnd.n5765 gnd.n5764 19.3944
R9257 gnd.n1769 gnd.n1748 19.3944
R9258 gnd.n5532 gnd.n1748 19.3944
R9259 gnd.n5532 gnd.n5531 19.3944
R9260 gnd.n4953 gnd.t29 19.1199
R9261 gnd.n4973 gnd.n2168 19.1199
R9262 gnd.n5060 gnd.n2122 19.1199
R9263 gnd.n5126 gnd.n2088 19.1199
R9264 gnd.n2043 gnd.n2031 19.1199
R9265 gnd.n5261 gnd.t15 19.1199
R9266 gnd.n5477 gnd.n5476 19.1199
R9267 gnd.n3291 gnd.t60 18.8012
R9268 gnd.n3276 gnd.t46 18.8012
R9269 gnd.n3135 gnd.n3134 18.4825
R9270 gnd.n5367 gnd.t120 18.4825
R9271 gnd.n5703 gnd.n5702 18.4247
R9272 gnd.n6035 gnd.n6034 18.4247
R9273 gnd.n5761 gnd.n5760 18.2308
R9274 gnd.n4526 gnd.n2294 18.2308
R9275 gnd.n251 gnd.n250 18.2308
R9276 gnd.n4088 gnd.n4026 18.2308
R9277 gnd.t8 gnd.n2815 18.1639
R9278 gnd.t306 gnd.n1380 18.1639
R9279 gnd.t22 gnd.n5376 18.1639
R9280 gnd.n4802 gnd.n1394 17.8452
R9281 gnd.n2231 gnd.n2222 17.8452
R9282 gnd.n5050 gnd.n5049 17.8452
R9283 gnd.n5136 gnd.n2074 17.8452
R9284 gnd.n5315 gnd.n5314 17.8452
R9285 gnd.n5348 gnd.n1960 17.8452
R9286 gnd.n2843 gnd.t315 17.5266
R9287 gnd.n4994 gnd.t53 17.5266
R9288 gnd.n5197 gnd.t312 17.5266
R9289 gnd.n3519 gnd.n3518 17.2079
R9290 gnd.n4822 gnd.t305 17.2079
R9291 gnd.t7 gnd.n1939 17.2079
R9292 gnd.n3242 gnd.t184 16.8893
R9293 gnd.n4251 gnd.t74 16.8893
R9294 gnd.t226 gnd.n1084 16.8893
R9295 gnd.t198 gnd.n549 16.8893
R9296 gnd.n162 gnd.t78 16.8893
R9297 gnd.n5685 gnd.n5682 16.6793
R9298 gnd.n436 gnd.n306 16.6793
R9299 gnd.n4168 gnd.n4165 16.6793
R9300 gnd.n4618 gnd.n4617 16.6793
R9301 gnd.n4845 gnd.n2241 16.5706
R9302 gnd.n4865 gnd.n4864 16.5706
R9303 gnd.n5005 gnd.n5004 16.5706
R9304 gnd.n4908 gnd.n2144 16.5706
R9305 gnd.n5174 gnd.n2069 16.5706
R9306 gnd.n5185 gnd.n2058 16.5706
R9307 gnd.n1979 gnd.n1973 16.5706
R9308 gnd.n5340 gnd.n5339 16.5706
R9309 gnd.n3070 gnd.t181 16.2519
R9310 gnd.n2770 gnd.t50 16.2519
R9311 gnd.n2265 gnd.t133 16.2519
R9312 gnd.t113 gnd.n1488 16.2519
R9313 gnd.n4947 gnd.t52 15.9333
R9314 gnd.n5284 gnd.t11 15.9333
R9315 gnd.n3758 gnd.n3756 15.6674
R9316 gnd.n3726 gnd.n3724 15.6674
R9317 gnd.n3694 gnd.n3692 15.6674
R9318 gnd.n3663 gnd.n3661 15.6674
R9319 gnd.n3631 gnd.n3629 15.6674
R9320 gnd.n3599 gnd.n3597 15.6674
R9321 gnd.n3567 gnd.n3565 15.6674
R9322 gnd.n3536 gnd.n3534 15.6674
R9323 gnd.n3061 gnd.t181 15.6146
R9324 gnd.t171 gnd.n2524 15.6146
R9325 gnd.t158 gnd.n2525 15.6146
R9326 gnd.t133 gnd.n1218 15.6146
R9327 gnd.n5504 gnd.t113 15.6146
R9328 gnd.n5642 gnd.n5637 15.3217
R9329 gnd.n491 gnd.n284 15.3217
R9330 gnd.n4126 gnd.n2441 15.3217
R9331 gnd.n4669 gnd.n4667 15.3217
R9332 gnd.n1821 gnd.n1820 15.0827
R9333 gnd.n1262 gnd.n1257 15.0481
R9334 gnd.n1831 gnd.n1830 15.0481
R9335 gnd.n3429 gnd.t314 14.9773
R9336 gnd.t74 gnd.n2422 14.9773
R9337 gnd.n4677 gnd.t106 14.9773
R9338 gnd.n5626 gnd.t82 14.9773
R9339 gnd.n6975 gnd.t78 14.9773
R9340 gnd.n4879 gnd.t0 14.6587
R9341 gnd.n1981 gnd.t21 14.6587
R9342 gnd.t62 gnd.n2567 14.34
R9343 gnd.n3507 gnd.t316 14.34
R9344 gnd.n5933 gnd.n1394 14.0214
R9345 gnd.t6 gnd.n2222 14.0214
R9346 gnd.n4986 gnd.n4984 14.0214
R9347 gnd.n5049 gnd.n2133 14.0214
R9348 gnd.n5136 gnd.n5135 14.0214
R9349 gnd.n5211 gnd.n2040 14.0214
R9350 gnd.n5315 gnd.t45 14.0214
R9351 gnd.n1960 gnd.n1953 14.0214
R9352 gnd.n5403 gnd.t65 14.0214
R9353 gnd.n3217 gnd.t48 13.7027
R9354 gnd.n4846 gnd.t2 13.7027
R9355 gnd.t4 gnd.n1967 13.7027
R9356 gnd.n2927 gnd.n2926 13.5763
R9357 gnd.n3872 gnd.n2481 13.5763
R9358 gnd.n3135 gnd.n2873 13.384
R9359 gnd.n1273 gnd.n1254 13.1884
R9360 gnd.n1268 gnd.n1267 13.1884
R9361 gnd.n1267 gnd.n1266 13.1884
R9362 gnd.n1824 gnd.n1819 13.1884
R9363 gnd.n1825 gnd.n1824 13.1884
R9364 gnd.n1269 gnd.n1256 13.146
R9365 gnd.n1265 gnd.n1256 13.146
R9366 gnd.n1823 gnd.n1822 13.146
R9367 gnd.n1823 gnd.n1818 13.146
R9368 gnd.n3759 gnd.n3755 12.8005
R9369 gnd.n3727 gnd.n3723 12.8005
R9370 gnd.n3695 gnd.n3691 12.8005
R9371 gnd.n3664 gnd.n3660 12.8005
R9372 gnd.n3632 gnd.n3628 12.8005
R9373 gnd.n3600 gnd.n3596 12.8005
R9374 gnd.n3568 gnd.n3564 12.8005
R9375 gnd.n3537 gnd.n3533 12.8005
R9376 gnd.n1361 gnd.n1276 12.7467
R9377 gnd.t96 gnd.t102 12.7467
R9378 gnd.n5939 gnd.n1380 12.7467
R9379 gnd.t24 gnd.n2241 12.7467
R9380 gnd.n4941 gnd.n4940 12.7467
R9381 gnd.n4973 gnd.n2167 12.7467
R9382 gnd.n5016 gnd.n2122 12.7467
R9383 gnd.n5017 gnd.t20 12.7467
R9384 gnd.t27 gnd.n2084 12.7467
R9385 gnd.n5127 gnd.n5126 12.7467
R9386 gnd.n5221 gnd.n2031 12.7467
R9387 gnd.n5296 gnd.n5294 12.7467
R9388 gnd.n5339 gnd.t17 12.7467
R9389 gnd.n5376 gnd.n1942 12.7467
R9390 gnd.n5369 gnd.t149 12.7467
R9391 gnd.n4941 gnd.t13 12.4281
R9392 gnd.n5294 gnd.t321 12.4281
R9393 gnd.n2926 gnd.n2921 12.4126
R9394 gnd.n3875 gnd.n3872 12.4126
R9395 gnd.n6027 gnd.n5964 12.1761
R9396 gnd.n1837 gnd.n1836 12.1761
R9397 gnd.n3763 gnd.n3762 12.0247
R9398 gnd.n3731 gnd.n3730 12.0247
R9399 gnd.n3699 gnd.n3698 12.0247
R9400 gnd.n3668 gnd.n3667 12.0247
R9401 gnd.n3636 gnd.n3635 12.0247
R9402 gnd.n3604 gnd.n3603 12.0247
R9403 gnd.n3572 gnd.n3571 12.0247
R9404 gnd.n3541 gnd.n3540 12.0247
R9405 gnd.n2414 gnd.t196 11.7908
R9406 gnd.t106 gnd.n1134 11.7908
R9407 gnd.n5573 gnd.t82 11.7908
R9408 gnd.n6987 gnd.t231 11.7908
R9409 gnd.n4777 gnd.n1280 11.4721
R9410 gnd.n2184 gnd.n2180 11.4721
R9411 gnd.n4932 gnd.n4930 11.4721
R9412 gnd.n5097 gnd.n2108 11.4721
R9413 gnd.n5105 gnd.n2102 11.4721
R9414 gnd.n5268 gnd.n2019 11.4721
R9415 gnd.n5260 gnd.n2003 11.4721
R9416 gnd.n5369 gnd.n5368 11.4721
R9417 gnd.n5485 gnd.n5484 11.4721
R9418 gnd.n3766 gnd.n3753 11.249
R9419 gnd.n3734 gnd.n3721 11.249
R9420 gnd.n3702 gnd.n3689 11.249
R9421 gnd.n3671 gnd.n3658 11.249
R9422 gnd.n3639 gnd.n3626 11.249
R9423 gnd.n3607 gnd.n3594 11.249
R9424 gnd.n3575 gnd.n3562 11.249
R9425 gnd.n3544 gnd.n3531 11.249
R9426 gnd.n3205 gnd.t48 11.1535
R9427 gnd.n2378 gnd.t244 11.1535
R9428 gnd.n7011 gnd.t213 11.1535
R9429 gnd.n1361 gnd.t137 10.8348
R9430 gnd.n4967 gnd.t44 10.8348
R9431 gnd.t44 gnd.n4966 10.8348
R9432 gnd.n2033 gnd.t32 10.8348
R9433 gnd.t32 gnd.n2032 10.8348
R9434 gnd.n5645 gnd.n5642 10.6672
R9435 gnd.n486 gnd.n284 10.6672
R9436 gnd.n4128 gnd.n4126 10.6672
R9437 gnd.n4667 gnd.n4666 10.6672
R9438 gnd.n5472 gnd.n5471 10.6151
R9439 gnd.n5471 gnd.n5468 10.6151
R9440 gnd.n5466 gnd.n5463 10.6151
R9441 gnd.n5463 gnd.n5462 10.6151
R9442 gnd.n5462 gnd.n5459 10.6151
R9443 gnd.n5459 gnd.n5458 10.6151
R9444 gnd.n5458 gnd.n5455 10.6151
R9445 gnd.n5455 gnd.n5454 10.6151
R9446 gnd.n5454 gnd.n5451 10.6151
R9447 gnd.n5451 gnd.n5450 10.6151
R9448 gnd.n5450 gnd.n5447 10.6151
R9449 gnd.n5447 gnd.n5446 10.6151
R9450 gnd.n5446 gnd.n5443 10.6151
R9451 gnd.n5443 gnd.n5442 10.6151
R9452 gnd.n5442 gnd.n5439 10.6151
R9453 gnd.n5439 gnd.n5438 10.6151
R9454 gnd.n5438 gnd.n5435 10.6151
R9455 gnd.n5435 gnd.n5434 10.6151
R9456 gnd.n5434 gnd.n5431 10.6151
R9457 gnd.n5431 gnd.n5430 10.6151
R9458 gnd.n5430 gnd.n5427 10.6151
R9459 gnd.n5427 gnd.n5426 10.6151
R9460 gnd.n5426 gnd.n5423 10.6151
R9461 gnd.n5423 gnd.n5422 10.6151
R9462 gnd.n5422 gnd.n5419 10.6151
R9463 gnd.n5419 gnd.n5418 10.6151
R9464 gnd.n5418 gnd.n5415 10.6151
R9465 gnd.n5415 gnd.n5414 10.6151
R9466 gnd.n5414 gnd.n5411 10.6151
R9467 gnd.n5411 gnd.n5410 10.6151
R9468 gnd.n1364 gnd.n1363 10.6151
R9469 gnd.n1365 gnd.n1364 10.6151
R9470 gnd.n1367 gnd.n1365 10.6151
R9471 gnd.n1368 gnd.n1367 10.6151
R9472 gnd.n5950 gnd.n1368 10.6151
R9473 gnd.n5950 gnd.n5949 10.6151
R9474 gnd.n5949 gnd.n5948 10.6151
R9475 gnd.n5948 gnd.n1369 10.6151
R9476 gnd.n4805 gnd.n1369 10.6151
R9477 gnd.n4807 gnd.n4805 10.6151
R9478 gnd.n4808 gnd.n4807 10.6151
R9479 gnd.n4810 gnd.n4808 10.6151
R9480 gnd.n4811 gnd.n4810 10.6151
R9481 gnd.n4813 gnd.n4811 10.6151
R9482 gnd.n4813 gnd.n4812 10.6151
R9483 gnd.n4812 gnd.n2239 10.6151
R9484 gnd.n4848 gnd.n2239 10.6151
R9485 gnd.n4849 gnd.n4848 10.6151
R9486 gnd.n4862 gnd.n4849 10.6151
R9487 gnd.n4862 gnd.n4861 10.6151
R9488 gnd.n4861 gnd.n4860 10.6151
R9489 gnd.n4860 gnd.n4850 10.6151
R9490 gnd.n4856 gnd.n4850 10.6151
R9491 gnd.n4856 gnd.n4855 10.6151
R9492 gnd.n4855 gnd.n4854 10.6151
R9493 gnd.n4854 gnd.n2182 10.6151
R9494 gnd.n4949 gnd.n2182 10.6151
R9495 gnd.n4950 gnd.n4949 10.6151
R9496 gnd.n4951 gnd.n4950 10.6151
R9497 gnd.n4951 gnd.n2174 10.6151
R9498 gnd.n4961 gnd.n2174 10.6151
R9499 gnd.n4962 gnd.n4961 10.6151
R9500 gnd.n4964 gnd.n4962 10.6151
R9501 gnd.n4964 gnd.n4963 10.6151
R9502 gnd.n4963 gnd.n2165 10.6151
R9503 gnd.n4976 gnd.n2165 10.6151
R9504 gnd.n4977 gnd.n4976 10.6151
R9505 gnd.n4982 gnd.n4977 10.6151
R9506 gnd.n4982 gnd.n4981 10.6151
R9507 gnd.n4981 gnd.n4980 10.6151
R9508 gnd.n4980 gnd.n4978 10.6151
R9509 gnd.n4978 gnd.n2140 10.6151
R9510 gnd.n5013 gnd.n2140 10.6151
R9511 gnd.n5014 gnd.n5013 10.6151
R9512 gnd.n5036 gnd.n5014 10.6151
R9513 gnd.n5036 gnd.n5035 10.6151
R9514 gnd.n5035 gnd.n5034 10.6151
R9515 gnd.n5034 gnd.n5033 10.6151
R9516 gnd.n5033 gnd.n5015 10.6151
R9517 gnd.n5028 gnd.n5015 10.6151
R9518 gnd.n5028 gnd.n5027 10.6151
R9519 gnd.n5027 gnd.n5026 10.6151
R9520 gnd.n5026 gnd.n5025 10.6151
R9521 gnd.n5025 gnd.n5023 10.6151
R9522 gnd.n5023 gnd.n5022 10.6151
R9523 gnd.n5022 gnd.n5020 10.6151
R9524 gnd.n5020 gnd.n5019 10.6151
R9525 gnd.n5019 gnd.n2092 10.6151
R9526 gnd.n5115 gnd.n2092 10.6151
R9527 gnd.n5116 gnd.n5115 10.6151
R9528 gnd.n5117 gnd.n5116 10.6151
R9529 gnd.n5117 gnd.n2076 10.6151
R9530 gnd.n5138 gnd.n2076 10.6151
R9531 gnd.n5139 gnd.n5138 10.6151
R9532 gnd.n5160 gnd.n5139 10.6151
R9533 gnd.n5160 gnd.n5159 10.6151
R9534 gnd.n5159 gnd.n5158 10.6151
R9535 gnd.n5158 gnd.n5140 10.6151
R9536 gnd.n5153 gnd.n5140 10.6151
R9537 gnd.n5153 gnd.n5152 10.6151
R9538 gnd.n5152 gnd.n5151 10.6151
R9539 gnd.n5151 gnd.n5150 10.6151
R9540 gnd.n5150 gnd.n5148 10.6151
R9541 gnd.n5148 gnd.n5147 10.6151
R9542 gnd.n5147 gnd.n5142 10.6151
R9543 gnd.n5143 gnd.n5142 10.6151
R9544 gnd.n5143 gnd.n2015 10.6151
R9545 gnd.n5270 gnd.n2015 10.6151
R9546 gnd.n5271 gnd.n5270 10.6151
R9547 gnd.n5273 gnd.n5271 10.6151
R9548 gnd.n5273 gnd.n5272 10.6151
R9549 gnd.n5272 gnd.n2001 10.6151
R9550 gnd.n5286 gnd.n2001 10.6151
R9551 gnd.n5287 gnd.n5286 10.6151
R9552 gnd.n5292 gnd.n5287 10.6151
R9553 gnd.n5292 gnd.n5291 10.6151
R9554 gnd.n5291 gnd.n5290 10.6151
R9555 gnd.n5290 gnd.n5288 10.6151
R9556 gnd.n5288 gnd.n1976 10.6151
R9557 gnd.n5323 gnd.n1976 10.6151
R9558 gnd.n5324 gnd.n5323 10.6151
R9559 gnd.n5331 gnd.n5324 10.6151
R9560 gnd.n5331 gnd.n5330 10.6151
R9561 gnd.n5330 gnd.n5329 10.6151
R9562 gnd.n5329 gnd.n5328 10.6151
R9563 gnd.n5328 gnd.n5326 10.6151
R9564 gnd.n5326 gnd.n5325 10.6151
R9565 gnd.n5325 gnd.n1951 10.6151
R9566 gnd.n5358 gnd.n1951 10.6151
R9567 gnd.n5359 gnd.n5358 10.6151
R9568 gnd.n5362 gnd.n5359 10.6151
R9569 gnd.n5363 gnd.n5362 10.6151
R9570 gnd.n5365 gnd.n5363 10.6151
R9571 gnd.n5365 gnd.n5364 10.6151
R9572 gnd.n5364 gnd.n1922 10.6151
R9573 gnd.n5399 gnd.n1922 10.6151
R9574 gnd.n5400 gnd.n5399 10.6151
R9575 gnd.n5401 gnd.n5400 10.6151
R9576 gnd.n5407 gnd.n5401 10.6151
R9577 gnd.n5408 gnd.n5407 10.6151
R9578 gnd.n1298 gnd.n1214 10.6151
R9579 gnd.n1301 gnd.n1298 10.6151
R9580 gnd.n1306 gnd.n1303 10.6151
R9581 gnd.n1307 gnd.n1306 10.6151
R9582 gnd.n1310 gnd.n1307 10.6151
R9583 gnd.n1311 gnd.n1310 10.6151
R9584 gnd.n1314 gnd.n1311 10.6151
R9585 gnd.n1315 gnd.n1314 10.6151
R9586 gnd.n1318 gnd.n1315 10.6151
R9587 gnd.n1319 gnd.n1318 10.6151
R9588 gnd.n1322 gnd.n1319 10.6151
R9589 gnd.n1323 gnd.n1322 10.6151
R9590 gnd.n1326 gnd.n1323 10.6151
R9591 gnd.n1327 gnd.n1326 10.6151
R9592 gnd.n1330 gnd.n1327 10.6151
R9593 gnd.n1331 gnd.n1330 10.6151
R9594 gnd.n1334 gnd.n1331 10.6151
R9595 gnd.n1335 gnd.n1334 10.6151
R9596 gnd.n1338 gnd.n1335 10.6151
R9597 gnd.n1339 gnd.n1338 10.6151
R9598 gnd.n1342 gnd.n1339 10.6151
R9599 gnd.n1343 gnd.n1342 10.6151
R9600 gnd.n1346 gnd.n1343 10.6151
R9601 gnd.n1347 gnd.n1346 10.6151
R9602 gnd.n1350 gnd.n1347 10.6151
R9603 gnd.n1351 gnd.n1350 10.6151
R9604 gnd.n1354 gnd.n1351 10.6151
R9605 gnd.n1355 gnd.n1354 10.6151
R9606 gnd.n1358 gnd.n1355 10.6151
R9607 gnd.n1359 gnd.n1358 10.6151
R9608 gnd.n6027 gnd.n6026 10.6151
R9609 gnd.n6026 gnd.n6025 10.6151
R9610 gnd.n6025 gnd.n6024 10.6151
R9611 gnd.n6024 gnd.n6022 10.6151
R9612 gnd.n6022 gnd.n6019 10.6151
R9613 gnd.n6019 gnd.n6018 10.6151
R9614 gnd.n6018 gnd.n6015 10.6151
R9615 gnd.n6015 gnd.n6014 10.6151
R9616 gnd.n6014 gnd.n6011 10.6151
R9617 gnd.n6011 gnd.n6010 10.6151
R9618 gnd.n6010 gnd.n6007 10.6151
R9619 gnd.n6007 gnd.n6006 10.6151
R9620 gnd.n6006 gnd.n6003 10.6151
R9621 gnd.n6003 gnd.n6002 10.6151
R9622 gnd.n6002 gnd.n5999 10.6151
R9623 gnd.n5999 gnd.n5998 10.6151
R9624 gnd.n5998 gnd.n5995 10.6151
R9625 gnd.n5995 gnd.n5994 10.6151
R9626 gnd.n5994 gnd.n5991 10.6151
R9627 gnd.n5991 gnd.n5990 10.6151
R9628 gnd.n5990 gnd.n5987 10.6151
R9629 gnd.n5987 gnd.n5986 10.6151
R9630 gnd.n5986 gnd.n5983 10.6151
R9631 gnd.n5983 gnd.n5982 10.6151
R9632 gnd.n5982 gnd.n5979 10.6151
R9633 gnd.n5979 gnd.n5978 10.6151
R9634 gnd.n5978 gnd.n5975 10.6151
R9635 gnd.n5975 gnd.n5974 10.6151
R9636 gnd.n5971 gnd.n5970 10.6151
R9637 gnd.n5970 gnd.n1215 10.6151
R9638 gnd.n1838 gnd.n1837 10.6151
R9639 gnd.n1841 gnd.n1838 10.6151
R9640 gnd.n1842 gnd.n1841 10.6151
R9641 gnd.n1845 gnd.n1842 10.6151
R9642 gnd.n1846 gnd.n1845 10.6151
R9643 gnd.n1849 gnd.n1846 10.6151
R9644 gnd.n1850 gnd.n1849 10.6151
R9645 gnd.n1853 gnd.n1850 10.6151
R9646 gnd.n1854 gnd.n1853 10.6151
R9647 gnd.n1857 gnd.n1854 10.6151
R9648 gnd.n1858 gnd.n1857 10.6151
R9649 gnd.n1861 gnd.n1858 10.6151
R9650 gnd.n1862 gnd.n1861 10.6151
R9651 gnd.n1865 gnd.n1862 10.6151
R9652 gnd.n1866 gnd.n1865 10.6151
R9653 gnd.n1869 gnd.n1866 10.6151
R9654 gnd.n1870 gnd.n1869 10.6151
R9655 gnd.n1873 gnd.n1870 10.6151
R9656 gnd.n1874 gnd.n1873 10.6151
R9657 gnd.n1877 gnd.n1874 10.6151
R9658 gnd.n1878 gnd.n1877 10.6151
R9659 gnd.n1881 gnd.n1878 10.6151
R9660 gnd.n1882 gnd.n1881 10.6151
R9661 gnd.n1885 gnd.n1882 10.6151
R9662 gnd.n1886 gnd.n1885 10.6151
R9663 gnd.n1889 gnd.n1886 10.6151
R9664 gnd.n1890 gnd.n1889 10.6151
R9665 gnd.n1893 gnd.n1890 10.6151
R9666 gnd.n1898 gnd.n1895 10.6151
R9667 gnd.n1899 gnd.n1898 10.6151
R9668 gnd.n5963 gnd.n5962 10.6151
R9669 gnd.n5962 gnd.n1274 10.6151
R9670 gnd.n4772 gnd.n1274 10.6151
R9671 gnd.n4774 gnd.n4772 10.6151
R9672 gnd.n4774 gnd.n4773 10.6151
R9673 gnd.n4773 gnd.n1374 10.6151
R9674 gnd.n5944 gnd.n1374 10.6151
R9675 gnd.n5944 gnd.n5943 10.6151
R9676 gnd.n5943 gnd.n5942 10.6151
R9677 gnd.n5942 gnd.n1375 10.6151
R9678 gnd.n4820 gnd.n1375 10.6151
R9679 gnd.n4820 gnd.n4819 10.6151
R9680 gnd.n4819 gnd.n4818 10.6151
R9681 gnd.n4818 gnd.n4797 10.6151
R9682 gnd.n4800 gnd.n4797 10.6151
R9683 gnd.n4800 gnd.n4799 10.6151
R9684 gnd.n4799 gnd.n2235 10.6151
R9685 gnd.n4868 gnd.n2235 10.6151
R9686 gnd.n4869 gnd.n4868 10.6151
R9687 gnd.n4875 gnd.n4869 10.6151
R9688 gnd.n4875 gnd.n4874 10.6151
R9689 gnd.n4874 gnd.n4873 10.6151
R9690 gnd.n4873 gnd.n4870 10.6151
R9691 gnd.n4870 gnd.n2187 10.6151
R9692 gnd.n4943 gnd.n2187 10.6151
R9693 gnd.n4944 gnd.n4943 10.6151
R9694 gnd.n4945 gnd.n4944 10.6151
R9695 gnd.n4945 gnd.n2178 10.6151
R9696 gnd.n4955 gnd.n2178 10.6151
R9697 gnd.n4956 gnd.n4955 10.6151
R9698 gnd.n4957 gnd.n4956 10.6151
R9699 gnd.n4957 gnd.n2170 10.6151
R9700 gnd.n4969 gnd.n2170 10.6151
R9701 gnd.n4970 gnd.n4969 10.6151
R9702 gnd.n4971 gnd.n4970 10.6151
R9703 gnd.n4971 gnd.n2160 10.6151
R9704 gnd.n4989 gnd.n2160 10.6151
R9705 gnd.n4990 gnd.n4989 10.6151
R9706 gnd.n4991 gnd.n4990 10.6151
R9707 gnd.n4991 gnd.n2146 10.6151
R9708 gnd.n5007 gnd.n2146 10.6151
R9709 gnd.n5008 gnd.n5007 10.6151
R9710 gnd.n5009 gnd.n5008 10.6151
R9711 gnd.n5009 gnd.n2136 10.6151
R9712 gnd.n5040 gnd.n2136 10.6151
R9713 gnd.n5041 gnd.n5040 10.6151
R9714 gnd.n5047 gnd.n5041 10.6151
R9715 gnd.n5047 gnd.n5046 10.6151
R9716 gnd.n5046 gnd.n5045 10.6151
R9717 gnd.n5045 gnd.n5042 10.6151
R9718 gnd.n5042 gnd.n2112 10.6151
R9719 gnd.n5092 gnd.n2112 10.6151
R9720 gnd.n5093 gnd.n5092 10.6151
R9721 gnd.n5094 gnd.n5093 10.6151
R9722 gnd.n5094 gnd.n2096 10.6151
R9723 gnd.n5108 gnd.n2096 10.6151
R9724 gnd.n5109 gnd.n5108 10.6151
R9725 gnd.n5110 gnd.n5109 10.6151
R9726 gnd.n5110 gnd.n2091 10.6151
R9727 gnd.n5124 gnd.n2091 10.6151
R9728 gnd.n5124 gnd.n5123 10.6151
R9729 gnd.n5123 gnd.n5122 10.6151
R9730 gnd.n5122 gnd.n2072 10.6151
R9731 gnd.n5165 gnd.n2072 10.6151
R9732 gnd.n5166 gnd.n5165 10.6151
R9733 gnd.n5172 gnd.n5166 10.6151
R9734 gnd.n5172 gnd.n5171 10.6151
R9735 gnd.n5171 gnd.n5170 10.6151
R9736 gnd.n5170 gnd.n5167 10.6151
R9737 gnd.n5167 gnd.n2047 10.6151
R9738 gnd.n5200 gnd.n2047 10.6151
R9739 gnd.n5201 gnd.n5200 10.6151
R9740 gnd.n5207 gnd.n5201 10.6151
R9741 gnd.n5207 gnd.n5206 10.6151
R9742 gnd.n5206 gnd.n5205 10.6151
R9743 gnd.n5205 gnd.n5202 10.6151
R9744 gnd.n5202 gnd.n2022 10.6151
R9745 gnd.n5266 gnd.n2022 10.6151
R9746 gnd.n5266 gnd.n5265 10.6151
R9747 gnd.n5265 gnd.n5264 10.6151
R9748 gnd.n5264 gnd.n5263 10.6151
R9749 gnd.n5263 gnd.n2023 10.6151
R9750 gnd.n2023 gnd.n1997 10.6151
R9751 gnd.n5299 gnd.n1997 10.6151
R9752 gnd.n5300 gnd.n5299 10.6151
R9753 gnd.n5301 gnd.n5300 10.6151
R9754 gnd.n5301 gnd.n1983 10.6151
R9755 gnd.n5317 gnd.n1983 10.6151
R9756 gnd.n5318 gnd.n5317 10.6151
R9757 gnd.n5319 gnd.n5318 10.6151
R9758 gnd.n5319 gnd.n1971 10.6151
R9759 gnd.n5335 gnd.n1971 10.6151
R9760 gnd.n5336 gnd.n5335 10.6151
R9761 gnd.n5337 gnd.n5336 10.6151
R9762 gnd.n5337 gnd.n1955 10.6151
R9763 gnd.n5351 gnd.n1955 10.6151
R9764 gnd.n5352 gnd.n5351 10.6151
R9765 gnd.n5353 gnd.n5352 10.6151
R9766 gnd.n5353 gnd.n1945 10.6151
R9767 gnd.n5374 gnd.n1945 10.6151
R9768 gnd.n5374 gnd.n5373 10.6151
R9769 gnd.n5373 gnd.n5372 10.6151
R9770 gnd.n5372 gnd.n1946 10.6151
R9771 gnd.n1948 gnd.n1946 10.6151
R9772 gnd.n1948 gnd.n1947 10.6151
R9773 gnd.n1947 gnd.n1795 10.6151
R9774 gnd.n5482 gnd.n1795 10.6151
R9775 gnd.n5482 gnd.n5481 10.6151
R9776 gnd.n5481 gnd.n5480 10.6151
R9777 gnd.n5480 gnd.n1796 10.6151
R9778 gnd.n3124 gnd.t317 10.5161
R9779 gnd.n2569 gnd.t62 10.5161
R9780 gnd.n3490 gnd.t316 10.5161
R9781 gnd.t258 gnd.n2339 10.5161
R9782 gnd.n2342 gnd.t246 10.5161
R9783 gnd.n6918 gnd.t216 10.5161
R9784 gnd.n6927 gnd.t237 10.5161
R9785 gnd.n3767 gnd.n3751 10.4732
R9786 gnd.n3735 gnd.n3719 10.4732
R9787 gnd.n3703 gnd.n3687 10.4732
R9788 gnd.n3672 gnd.n3656 10.4732
R9789 gnd.n3640 gnd.n3624 10.4732
R9790 gnd.n3608 gnd.n3592 10.4732
R9791 gnd.n3576 gnd.n3560 10.4732
R9792 gnd.n3545 gnd.n3529 10.4732
R9793 gnd.n4777 gnd.n4776 10.1975
R9794 gnd.n4788 gnd.n1292 10.1975
R9795 gnd.n4953 gnd.n2180 10.1975
R9796 gnd.n5097 gnd.n5096 10.1975
R9797 gnd.n5106 gnd.n5105 10.1975
R9798 gnd.n5261 gnd.n5260 10.1975
R9799 gnd.n5368 gnd.n5367 10.1975
R9800 gnd.n5485 gnd.n1790 10.1975
R9801 gnd.t314 gnd.n2586 9.87883
R9802 gnd.t224 gnd.n2375 9.87883
R9803 gnd.n6141 gnd.n1050 9.87883
R9804 gnd.n4387 gnd.t226 9.87883
R9805 gnd.n1725 gnd.t198 9.87883
R9806 gnd.n6848 gnd.n509 9.87883
R9807 gnd.n7005 gnd.t253 9.87883
R9808 gnd.n3771 gnd.n3770 9.69747
R9809 gnd.n3739 gnd.n3738 9.69747
R9810 gnd.n3707 gnd.n3706 9.69747
R9811 gnd.n3676 gnd.n3675 9.69747
R9812 gnd.n3644 gnd.n3643 9.69747
R9813 gnd.n3612 gnd.n3611 9.69747
R9814 gnd.n3580 gnd.n3579 9.69747
R9815 gnd.n3549 gnd.n3548 9.69747
R9816 gnd.n4905 gnd.t28 9.56018
R9817 gnd.n2060 gnd.t10 9.56018
R9818 gnd.n3777 gnd.n3776 9.45567
R9819 gnd.n3745 gnd.n3744 9.45567
R9820 gnd.n3713 gnd.n3712 9.45567
R9821 gnd.n3682 gnd.n3681 9.45567
R9822 gnd.n3650 gnd.n3649 9.45567
R9823 gnd.n3618 gnd.n3617 9.45567
R9824 gnd.n3586 gnd.n3585 9.45567
R9825 gnd.n3555 gnd.n3554 9.45567
R9826 gnd.n5682 gnd.n5681 9.30959
R9827 gnd.n442 gnd.n306 9.30959
R9828 gnd.n4165 gnd.n4164 9.30959
R9829 gnd.n4621 gnd.n4618 9.30959
R9830 gnd.n3776 gnd.n3775 9.3005
R9831 gnd.n3749 gnd.n3748 9.3005
R9832 gnd.n3770 gnd.n3769 9.3005
R9833 gnd.n3768 gnd.n3767 9.3005
R9834 gnd.n3753 gnd.n3752 9.3005
R9835 gnd.n3762 gnd.n3761 9.3005
R9836 gnd.n3760 gnd.n3759 9.3005
R9837 gnd.n3744 gnd.n3743 9.3005
R9838 gnd.n3717 gnd.n3716 9.3005
R9839 gnd.n3738 gnd.n3737 9.3005
R9840 gnd.n3736 gnd.n3735 9.3005
R9841 gnd.n3721 gnd.n3720 9.3005
R9842 gnd.n3730 gnd.n3729 9.3005
R9843 gnd.n3728 gnd.n3727 9.3005
R9844 gnd.n3712 gnd.n3711 9.3005
R9845 gnd.n3685 gnd.n3684 9.3005
R9846 gnd.n3706 gnd.n3705 9.3005
R9847 gnd.n3704 gnd.n3703 9.3005
R9848 gnd.n3689 gnd.n3688 9.3005
R9849 gnd.n3698 gnd.n3697 9.3005
R9850 gnd.n3696 gnd.n3695 9.3005
R9851 gnd.n3681 gnd.n3680 9.3005
R9852 gnd.n3654 gnd.n3653 9.3005
R9853 gnd.n3675 gnd.n3674 9.3005
R9854 gnd.n3673 gnd.n3672 9.3005
R9855 gnd.n3658 gnd.n3657 9.3005
R9856 gnd.n3667 gnd.n3666 9.3005
R9857 gnd.n3665 gnd.n3664 9.3005
R9858 gnd.n3649 gnd.n3648 9.3005
R9859 gnd.n3622 gnd.n3621 9.3005
R9860 gnd.n3643 gnd.n3642 9.3005
R9861 gnd.n3641 gnd.n3640 9.3005
R9862 gnd.n3626 gnd.n3625 9.3005
R9863 gnd.n3635 gnd.n3634 9.3005
R9864 gnd.n3633 gnd.n3632 9.3005
R9865 gnd.n3617 gnd.n3616 9.3005
R9866 gnd.n3590 gnd.n3589 9.3005
R9867 gnd.n3611 gnd.n3610 9.3005
R9868 gnd.n3609 gnd.n3608 9.3005
R9869 gnd.n3594 gnd.n3593 9.3005
R9870 gnd.n3603 gnd.n3602 9.3005
R9871 gnd.n3601 gnd.n3600 9.3005
R9872 gnd.n3585 gnd.n3584 9.3005
R9873 gnd.n3558 gnd.n3557 9.3005
R9874 gnd.n3579 gnd.n3578 9.3005
R9875 gnd.n3577 gnd.n3576 9.3005
R9876 gnd.n3562 gnd.n3561 9.3005
R9877 gnd.n3571 gnd.n3570 9.3005
R9878 gnd.n3569 gnd.n3568 9.3005
R9879 gnd.n3554 gnd.n3553 9.3005
R9880 gnd.n3527 gnd.n3526 9.3005
R9881 gnd.n3548 gnd.n3547 9.3005
R9882 gnd.n3546 gnd.n3545 9.3005
R9883 gnd.n3531 gnd.n3530 9.3005
R9884 gnd.n3540 gnd.n3539 9.3005
R9885 gnd.n3538 gnd.n3537 9.3005
R9886 gnd.n3902 gnd.n3901 9.3005
R9887 gnd.n3900 gnd.n2469 9.3005
R9888 gnd.n3899 gnd.n3898 9.3005
R9889 gnd.n3895 gnd.n2470 9.3005
R9890 gnd.n3892 gnd.n2471 9.3005
R9891 gnd.n3891 gnd.n2472 9.3005
R9892 gnd.n3888 gnd.n2473 9.3005
R9893 gnd.n3887 gnd.n2474 9.3005
R9894 gnd.n3884 gnd.n2475 9.3005
R9895 gnd.n3883 gnd.n2476 9.3005
R9896 gnd.n3880 gnd.n2477 9.3005
R9897 gnd.n3879 gnd.n2478 9.3005
R9898 gnd.n3876 gnd.n2479 9.3005
R9899 gnd.n3875 gnd.n2480 9.3005
R9900 gnd.n3872 gnd.n3871 9.3005
R9901 gnd.n3870 gnd.n2481 9.3005
R9902 gnd.n3903 gnd.n2468 9.3005
R9903 gnd.n3143 gnd.n3142 9.3005
R9904 gnd.n2847 gnd.n2846 9.3005
R9905 gnd.n3170 gnd.n3169 9.3005
R9906 gnd.n3171 gnd.n2845 9.3005
R9907 gnd.n3175 gnd.n3172 9.3005
R9908 gnd.n3174 gnd.n3173 9.3005
R9909 gnd.n2819 gnd.n2818 9.3005
R9910 gnd.n3200 gnd.n3199 9.3005
R9911 gnd.n3201 gnd.n2817 9.3005
R9912 gnd.n3203 gnd.n3202 9.3005
R9913 gnd.n2797 gnd.n2796 9.3005
R9914 gnd.n3231 gnd.n3230 9.3005
R9915 gnd.n3232 gnd.n2795 9.3005
R9916 gnd.n3240 gnd.n3233 9.3005
R9917 gnd.n3239 gnd.n3234 9.3005
R9918 gnd.n3238 gnd.n3236 9.3005
R9919 gnd.n3235 gnd.n2744 9.3005
R9920 gnd.n3288 gnd.n2745 9.3005
R9921 gnd.n3287 gnd.n2746 9.3005
R9922 gnd.n3286 gnd.n2747 9.3005
R9923 gnd.n2766 gnd.n2748 9.3005
R9924 gnd.n2768 gnd.n2767 9.3005
R9925 gnd.n2666 gnd.n2665 9.3005
R9926 gnd.n3326 gnd.n3325 9.3005
R9927 gnd.n3327 gnd.n2664 9.3005
R9928 gnd.n3331 gnd.n3328 9.3005
R9929 gnd.n3330 gnd.n3329 9.3005
R9930 gnd.n2639 gnd.n2638 9.3005
R9931 gnd.n3366 gnd.n3365 9.3005
R9932 gnd.n3367 gnd.n2637 9.3005
R9933 gnd.n3371 gnd.n3368 9.3005
R9934 gnd.n3370 gnd.n3369 9.3005
R9935 gnd.n2612 gnd.n2611 9.3005
R9936 gnd.n3411 gnd.n3410 9.3005
R9937 gnd.n3412 gnd.n2610 9.3005
R9938 gnd.n3416 gnd.n3413 9.3005
R9939 gnd.n3415 gnd.n3414 9.3005
R9940 gnd.n2584 gnd.n2583 9.3005
R9941 gnd.n3451 gnd.n3450 9.3005
R9942 gnd.n3452 gnd.n2582 9.3005
R9943 gnd.n3456 gnd.n3453 9.3005
R9944 gnd.n3455 gnd.n3454 9.3005
R9945 gnd.n2557 gnd.n2556 9.3005
R9946 gnd.n3500 gnd.n3499 9.3005
R9947 gnd.n3501 gnd.n2555 9.3005
R9948 gnd.n3505 gnd.n3502 9.3005
R9949 gnd.n3504 gnd.n3503 9.3005
R9950 gnd.n2530 gnd.n2529 9.3005
R9951 gnd.n3795 gnd.n3794 9.3005
R9952 gnd.n3796 gnd.n2528 9.3005
R9953 gnd.n3802 gnd.n3797 9.3005
R9954 gnd.n3801 gnd.n3798 9.3005
R9955 gnd.n3800 gnd.n3799 9.3005
R9956 gnd.n3144 gnd.n3141 9.3005
R9957 gnd.n2926 gnd.n2885 9.3005
R9958 gnd.n2921 gnd.n2920 9.3005
R9959 gnd.n2919 gnd.n2886 9.3005
R9960 gnd.n2918 gnd.n2917 9.3005
R9961 gnd.n2914 gnd.n2887 9.3005
R9962 gnd.n2911 gnd.n2910 9.3005
R9963 gnd.n2909 gnd.n2888 9.3005
R9964 gnd.n2908 gnd.n2907 9.3005
R9965 gnd.n2904 gnd.n2889 9.3005
R9966 gnd.n2901 gnd.n2900 9.3005
R9967 gnd.n2899 gnd.n2890 9.3005
R9968 gnd.n2898 gnd.n2897 9.3005
R9969 gnd.n2894 gnd.n2892 9.3005
R9970 gnd.n2891 gnd.n2871 9.3005
R9971 gnd.n3138 gnd.n2870 9.3005
R9972 gnd.n3140 gnd.n3139 9.3005
R9973 gnd.n2928 gnd.n2927 9.3005
R9974 gnd.n3151 gnd.n2857 9.3005
R9975 gnd.n3158 gnd.n2858 9.3005
R9976 gnd.n3160 gnd.n3159 9.3005
R9977 gnd.n3161 gnd.n2838 9.3005
R9978 gnd.n3180 gnd.n3179 9.3005
R9979 gnd.n3182 gnd.n2830 9.3005
R9980 gnd.n3189 gnd.n2832 9.3005
R9981 gnd.n3190 gnd.n2827 9.3005
R9982 gnd.n3192 gnd.n3191 9.3005
R9983 gnd.n2828 gnd.n2813 9.3005
R9984 gnd.n3208 gnd.n2811 9.3005
R9985 gnd.n3212 gnd.n3211 9.3005
R9986 gnd.n3210 gnd.n2787 9.3005
R9987 gnd.n3247 gnd.n2786 9.3005
R9988 gnd.n3250 gnd.n3249 9.3005
R9989 gnd.n2783 gnd.n2782 9.3005
R9990 gnd.n3256 gnd.n2784 9.3005
R9991 gnd.n3258 gnd.n3257 9.3005
R9992 gnd.n3260 gnd.n2781 9.3005
R9993 gnd.n3263 gnd.n3262 9.3005
R9994 gnd.n3266 gnd.n3264 9.3005
R9995 gnd.n3268 gnd.n3267 9.3005
R9996 gnd.n3274 gnd.n3269 9.3005
R9997 gnd.n3273 gnd.n3272 9.3005
R9998 gnd.n2657 gnd.n2656 9.3005
R9999 gnd.n3340 gnd.n3339 9.3005
R10000 gnd.n3341 gnd.n2650 9.3005
R10001 gnd.n3349 gnd.n2649 9.3005
R10002 gnd.n3352 gnd.n3351 9.3005
R10003 gnd.n3354 gnd.n3353 9.3005
R10004 gnd.n3357 gnd.n2632 9.3005
R10005 gnd.n3355 gnd.n2630 9.3005
R10006 gnd.n3377 gnd.n2628 9.3005
R10007 gnd.n3379 gnd.n3378 9.3005
R10008 gnd.n2602 gnd.n2601 9.3005
R10009 gnd.n3425 gnd.n3424 9.3005
R10010 gnd.n3426 gnd.n2595 9.3005
R10011 gnd.n3434 gnd.n2594 9.3005
R10012 gnd.n3437 gnd.n3436 9.3005
R10013 gnd.n3439 gnd.n3438 9.3005
R10014 gnd.n3442 gnd.n2577 9.3005
R10015 gnd.n3440 gnd.n2575 9.3005
R10016 gnd.n3462 gnd.n2573 9.3005
R10017 gnd.n3464 gnd.n3463 9.3005
R10018 gnd.n2548 gnd.n2547 9.3005
R10019 gnd.n3514 gnd.n3513 9.3005
R10020 gnd.n3515 gnd.n2541 9.3005
R10021 gnd.n3524 gnd.n2540 9.3005
R10022 gnd.n3783 gnd.n3782 9.3005
R10023 gnd.n3785 gnd.n3784 9.3005
R10024 gnd.n3786 gnd.n2521 9.3005
R10025 gnd.n3810 gnd.n3809 9.3005
R10026 gnd.n2522 gnd.n2484 9.3005
R10027 gnd.n3149 gnd.n3148 9.3005
R10028 gnd.n3866 gnd.n2485 9.3005
R10029 gnd.n3865 gnd.n2487 9.3005
R10030 gnd.n3862 gnd.n2488 9.3005
R10031 gnd.n3861 gnd.n2489 9.3005
R10032 gnd.n3858 gnd.n2490 9.3005
R10033 gnd.n3857 gnd.n2491 9.3005
R10034 gnd.n3854 gnd.n2492 9.3005
R10035 gnd.n3853 gnd.n2493 9.3005
R10036 gnd.n3850 gnd.n2494 9.3005
R10037 gnd.n3849 gnd.n2495 9.3005
R10038 gnd.n3846 gnd.n2496 9.3005
R10039 gnd.n3845 gnd.n2497 9.3005
R10040 gnd.n3842 gnd.n2498 9.3005
R10041 gnd.n3841 gnd.n2499 9.3005
R10042 gnd.n3838 gnd.n2500 9.3005
R10043 gnd.n3837 gnd.n2501 9.3005
R10044 gnd.n3834 gnd.n2502 9.3005
R10045 gnd.n3833 gnd.n2503 9.3005
R10046 gnd.n3830 gnd.n2504 9.3005
R10047 gnd.n3829 gnd.n2505 9.3005
R10048 gnd.n3826 gnd.n2506 9.3005
R10049 gnd.n3825 gnd.n2507 9.3005
R10050 gnd.n3822 gnd.n2511 9.3005
R10051 gnd.n3821 gnd.n2512 9.3005
R10052 gnd.n3818 gnd.n2513 9.3005
R10053 gnd.n3817 gnd.n2514 9.3005
R10054 gnd.n3868 gnd.n3867 9.3005
R10055 gnd.n3318 gnd.n3302 9.3005
R10056 gnd.n3317 gnd.n3303 9.3005
R10057 gnd.n3316 gnd.n3304 9.3005
R10058 gnd.n3314 gnd.n3305 9.3005
R10059 gnd.n3313 gnd.n3306 9.3005
R10060 gnd.n3311 gnd.n3307 9.3005
R10061 gnd.n3310 gnd.n3308 9.3005
R10062 gnd.n2620 gnd.n2619 9.3005
R10063 gnd.n3387 gnd.n3386 9.3005
R10064 gnd.n3388 gnd.n2618 9.3005
R10065 gnd.n3405 gnd.n3389 9.3005
R10066 gnd.n3404 gnd.n3390 9.3005
R10067 gnd.n3403 gnd.n3391 9.3005
R10068 gnd.n3401 gnd.n3392 9.3005
R10069 gnd.n3400 gnd.n3393 9.3005
R10070 gnd.n3398 gnd.n3394 9.3005
R10071 gnd.n3397 gnd.n3395 9.3005
R10072 gnd.n2564 gnd.n2563 9.3005
R10073 gnd.n3472 gnd.n3471 9.3005
R10074 gnd.n3473 gnd.n2562 9.3005
R10075 gnd.n3494 gnd.n3474 9.3005
R10076 gnd.n3493 gnd.n3475 9.3005
R10077 gnd.n3492 gnd.n3476 9.3005
R10078 gnd.n3489 gnd.n3477 9.3005
R10079 gnd.n3488 gnd.n3478 9.3005
R10080 gnd.n3486 gnd.n3479 9.3005
R10081 gnd.n3485 gnd.n3480 9.3005
R10082 gnd.n3483 gnd.n3482 9.3005
R10083 gnd.n3481 gnd.n2516 9.3005
R10084 gnd.n3059 gnd.n3058 9.3005
R10085 gnd.n2949 gnd.n2948 9.3005
R10086 gnd.n3073 gnd.n3072 9.3005
R10087 gnd.n3074 gnd.n2947 9.3005
R10088 gnd.n3076 gnd.n3075 9.3005
R10089 gnd.n2937 gnd.n2936 9.3005
R10090 gnd.n3089 gnd.n3088 9.3005
R10091 gnd.n3090 gnd.n2935 9.3005
R10092 gnd.n3122 gnd.n3091 9.3005
R10093 gnd.n3121 gnd.n3092 9.3005
R10094 gnd.n3120 gnd.n3093 9.3005
R10095 gnd.n3119 gnd.n3094 9.3005
R10096 gnd.n3116 gnd.n3095 9.3005
R10097 gnd.n3115 gnd.n3096 9.3005
R10098 gnd.n3114 gnd.n3097 9.3005
R10099 gnd.n3112 gnd.n3098 9.3005
R10100 gnd.n3111 gnd.n3099 9.3005
R10101 gnd.n3108 gnd.n3100 9.3005
R10102 gnd.n3107 gnd.n3101 9.3005
R10103 gnd.n3106 gnd.n3102 9.3005
R10104 gnd.n3104 gnd.n3103 9.3005
R10105 gnd.n2803 gnd.n2802 9.3005
R10106 gnd.n3220 gnd.n3219 9.3005
R10107 gnd.n3221 gnd.n2801 9.3005
R10108 gnd.n3225 gnd.n3222 9.3005
R10109 gnd.n3224 gnd.n3223 9.3005
R10110 gnd.n2725 gnd.n2724 9.3005
R10111 gnd.n3300 gnd.n3299 9.3005
R10112 gnd.n3057 gnd.n2958 9.3005
R10113 gnd.n2960 gnd.n2959 9.3005
R10114 gnd.n3004 gnd.n3002 9.3005
R10115 gnd.n3005 gnd.n3001 9.3005
R10116 gnd.n3008 gnd.n2997 9.3005
R10117 gnd.n3009 gnd.n2996 9.3005
R10118 gnd.n3012 gnd.n2995 9.3005
R10119 gnd.n3013 gnd.n2994 9.3005
R10120 gnd.n3016 gnd.n2993 9.3005
R10121 gnd.n3017 gnd.n2992 9.3005
R10122 gnd.n3020 gnd.n2991 9.3005
R10123 gnd.n3021 gnd.n2990 9.3005
R10124 gnd.n3024 gnd.n2989 9.3005
R10125 gnd.n3025 gnd.n2988 9.3005
R10126 gnd.n3028 gnd.n2987 9.3005
R10127 gnd.n3029 gnd.n2986 9.3005
R10128 gnd.n3032 gnd.n2985 9.3005
R10129 gnd.n3033 gnd.n2984 9.3005
R10130 gnd.n3036 gnd.n2983 9.3005
R10131 gnd.n3037 gnd.n2982 9.3005
R10132 gnd.n3040 gnd.n2981 9.3005
R10133 gnd.n3041 gnd.n2980 9.3005
R10134 gnd.n3044 gnd.n2979 9.3005
R10135 gnd.n3046 gnd.n2978 9.3005
R10136 gnd.n3047 gnd.n2977 9.3005
R10137 gnd.n3048 gnd.n2976 9.3005
R10138 gnd.n3049 gnd.n2975 9.3005
R10139 gnd.n3056 gnd.n3055 9.3005
R10140 gnd.n3065 gnd.n3064 9.3005
R10141 gnd.n3066 gnd.n2952 9.3005
R10142 gnd.n3068 gnd.n3067 9.3005
R10143 gnd.n2943 gnd.n2942 9.3005
R10144 gnd.n3081 gnd.n3080 9.3005
R10145 gnd.n3082 gnd.n2941 9.3005
R10146 gnd.n3084 gnd.n3083 9.3005
R10147 gnd.n2930 gnd.n2929 9.3005
R10148 gnd.n3127 gnd.n3126 9.3005
R10149 gnd.n3128 gnd.n2884 9.3005
R10150 gnd.n3132 gnd.n3130 9.3005
R10151 gnd.n3131 gnd.n2863 9.3005
R10152 gnd.n3150 gnd.n2862 9.3005
R10153 gnd.n3153 gnd.n3152 9.3005
R10154 gnd.n2856 gnd.n2855 9.3005
R10155 gnd.n3164 gnd.n3162 9.3005
R10156 gnd.n3163 gnd.n2837 9.3005
R10157 gnd.n3181 gnd.n2836 9.3005
R10158 gnd.n3184 gnd.n3183 9.3005
R10159 gnd.n2831 gnd.n2826 9.3005
R10160 gnd.n3194 gnd.n3193 9.3005
R10161 gnd.n2829 gnd.n2809 9.3005
R10162 gnd.n3215 gnd.n2810 9.3005
R10163 gnd.n3214 gnd.n3213 9.3005
R10164 gnd.n2812 gnd.n2788 9.3005
R10165 gnd.n3246 gnd.n3245 9.3005
R10166 gnd.n3248 gnd.n2733 9.3005
R10167 gnd.n3295 gnd.n2734 9.3005
R10168 gnd.n3294 gnd.n2735 9.3005
R10169 gnd.n3293 gnd.n2736 9.3005
R10170 gnd.n3259 gnd.n2737 9.3005
R10171 gnd.n3261 gnd.n2755 9.3005
R10172 gnd.n3281 gnd.n2756 9.3005
R10173 gnd.n3280 gnd.n2757 9.3005
R10174 gnd.n3279 gnd.n2758 9.3005
R10175 gnd.n3270 gnd.n2759 9.3005
R10176 gnd.n3271 gnd.n2658 9.3005
R10177 gnd.n3337 gnd.n3336 9.3005
R10178 gnd.n3338 gnd.n2651 9.3005
R10179 gnd.n3348 gnd.n3347 9.3005
R10180 gnd.n3350 gnd.n2647 9.3005
R10181 gnd.n3360 gnd.n2648 9.3005
R10182 gnd.n3359 gnd.n3358 9.3005
R10183 gnd.n3356 gnd.n2626 9.3005
R10184 gnd.n3382 gnd.n2627 9.3005
R10185 gnd.n3381 gnd.n3380 9.3005
R10186 gnd.n2629 gnd.n2603 9.3005
R10187 gnd.n3422 gnd.n3421 9.3005
R10188 gnd.n3423 gnd.n2596 9.3005
R10189 gnd.n3433 gnd.n3432 9.3005
R10190 gnd.n3435 gnd.n2592 9.3005
R10191 gnd.n3445 gnd.n2593 9.3005
R10192 gnd.n3444 gnd.n3443 9.3005
R10193 gnd.n3441 gnd.n2571 9.3005
R10194 gnd.n3467 gnd.n2572 9.3005
R10195 gnd.n3466 gnd.n3465 9.3005
R10196 gnd.n2574 gnd.n2549 9.3005
R10197 gnd.n3511 gnd.n3510 9.3005
R10198 gnd.n3512 gnd.n2542 9.3005
R10199 gnd.n3523 gnd.n3522 9.3005
R10200 gnd.n3781 gnd.n2538 9.3005
R10201 gnd.n3789 gnd.n2539 9.3005
R10202 gnd.n3788 gnd.n3787 9.3005
R10203 gnd.n2520 gnd.n2519 9.3005
R10204 gnd.n3812 gnd.n3811 9.3005
R10205 gnd.n2954 gnd.n2953 9.3005
R10206 gnd.n6313 gnd.n880 9.3005
R10207 gnd.n6315 gnd.n6314 9.3005
R10208 gnd.n876 gnd.n875 9.3005
R10209 gnd.n6322 gnd.n6321 9.3005
R10210 gnd.n6323 gnd.n874 9.3005
R10211 gnd.n6325 gnd.n6324 9.3005
R10212 gnd.n870 gnd.n869 9.3005
R10213 gnd.n6332 gnd.n6331 9.3005
R10214 gnd.n6333 gnd.n868 9.3005
R10215 gnd.n6335 gnd.n6334 9.3005
R10216 gnd.n864 gnd.n863 9.3005
R10217 gnd.n6342 gnd.n6341 9.3005
R10218 gnd.n6343 gnd.n862 9.3005
R10219 gnd.n6345 gnd.n6344 9.3005
R10220 gnd.n858 gnd.n857 9.3005
R10221 gnd.n6352 gnd.n6351 9.3005
R10222 gnd.n6353 gnd.n856 9.3005
R10223 gnd.n6355 gnd.n6354 9.3005
R10224 gnd.n852 gnd.n851 9.3005
R10225 gnd.n6362 gnd.n6361 9.3005
R10226 gnd.n6363 gnd.n850 9.3005
R10227 gnd.n6365 gnd.n6364 9.3005
R10228 gnd.n846 gnd.n845 9.3005
R10229 gnd.n6372 gnd.n6371 9.3005
R10230 gnd.n6373 gnd.n844 9.3005
R10231 gnd.n6375 gnd.n6374 9.3005
R10232 gnd.n840 gnd.n839 9.3005
R10233 gnd.n6382 gnd.n6381 9.3005
R10234 gnd.n6383 gnd.n838 9.3005
R10235 gnd.n6385 gnd.n6384 9.3005
R10236 gnd.n834 gnd.n833 9.3005
R10237 gnd.n6392 gnd.n6391 9.3005
R10238 gnd.n6393 gnd.n832 9.3005
R10239 gnd.n6395 gnd.n6394 9.3005
R10240 gnd.n828 gnd.n827 9.3005
R10241 gnd.n6402 gnd.n6401 9.3005
R10242 gnd.n6403 gnd.n826 9.3005
R10243 gnd.n6405 gnd.n6404 9.3005
R10244 gnd.n822 gnd.n821 9.3005
R10245 gnd.n6412 gnd.n6411 9.3005
R10246 gnd.n6413 gnd.n820 9.3005
R10247 gnd.n6415 gnd.n6414 9.3005
R10248 gnd.n816 gnd.n815 9.3005
R10249 gnd.n6422 gnd.n6421 9.3005
R10250 gnd.n6423 gnd.n814 9.3005
R10251 gnd.n6425 gnd.n6424 9.3005
R10252 gnd.n810 gnd.n809 9.3005
R10253 gnd.n6432 gnd.n6431 9.3005
R10254 gnd.n6433 gnd.n808 9.3005
R10255 gnd.n6435 gnd.n6434 9.3005
R10256 gnd.n804 gnd.n803 9.3005
R10257 gnd.n6442 gnd.n6441 9.3005
R10258 gnd.n6443 gnd.n802 9.3005
R10259 gnd.n6445 gnd.n6444 9.3005
R10260 gnd.n798 gnd.n797 9.3005
R10261 gnd.n6452 gnd.n6451 9.3005
R10262 gnd.n6453 gnd.n796 9.3005
R10263 gnd.n6455 gnd.n6454 9.3005
R10264 gnd.n792 gnd.n791 9.3005
R10265 gnd.n6462 gnd.n6461 9.3005
R10266 gnd.n6463 gnd.n790 9.3005
R10267 gnd.n6465 gnd.n6464 9.3005
R10268 gnd.n786 gnd.n785 9.3005
R10269 gnd.n6472 gnd.n6471 9.3005
R10270 gnd.n6473 gnd.n784 9.3005
R10271 gnd.n6475 gnd.n6474 9.3005
R10272 gnd.n780 gnd.n779 9.3005
R10273 gnd.n6482 gnd.n6481 9.3005
R10274 gnd.n6483 gnd.n778 9.3005
R10275 gnd.n6485 gnd.n6484 9.3005
R10276 gnd.n774 gnd.n773 9.3005
R10277 gnd.n6492 gnd.n6491 9.3005
R10278 gnd.n6493 gnd.n772 9.3005
R10279 gnd.n6495 gnd.n6494 9.3005
R10280 gnd.n768 gnd.n767 9.3005
R10281 gnd.n6502 gnd.n6501 9.3005
R10282 gnd.n6503 gnd.n766 9.3005
R10283 gnd.n6505 gnd.n6504 9.3005
R10284 gnd.n762 gnd.n761 9.3005
R10285 gnd.n6512 gnd.n6511 9.3005
R10286 gnd.n6513 gnd.n760 9.3005
R10287 gnd.n6515 gnd.n6514 9.3005
R10288 gnd.n756 gnd.n755 9.3005
R10289 gnd.n6522 gnd.n6521 9.3005
R10290 gnd.n6523 gnd.n754 9.3005
R10291 gnd.n6525 gnd.n6524 9.3005
R10292 gnd.n750 gnd.n749 9.3005
R10293 gnd.n6532 gnd.n6531 9.3005
R10294 gnd.n6533 gnd.n748 9.3005
R10295 gnd.n6535 gnd.n6534 9.3005
R10296 gnd.n744 gnd.n743 9.3005
R10297 gnd.n6542 gnd.n6541 9.3005
R10298 gnd.n6543 gnd.n742 9.3005
R10299 gnd.n6545 gnd.n6544 9.3005
R10300 gnd.n738 gnd.n737 9.3005
R10301 gnd.n6552 gnd.n6551 9.3005
R10302 gnd.n6553 gnd.n736 9.3005
R10303 gnd.n6555 gnd.n6554 9.3005
R10304 gnd.n732 gnd.n731 9.3005
R10305 gnd.n6562 gnd.n6561 9.3005
R10306 gnd.n6563 gnd.n730 9.3005
R10307 gnd.n6565 gnd.n6564 9.3005
R10308 gnd.n726 gnd.n725 9.3005
R10309 gnd.n6572 gnd.n6571 9.3005
R10310 gnd.n6573 gnd.n724 9.3005
R10311 gnd.n6575 gnd.n6574 9.3005
R10312 gnd.n720 gnd.n719 9.3005
R10313 gnd.n6582 gnd.n6581 9.3005
R10314 gnd.n6583 gnd.n718 9.3005
R10315 gnd.n6585 gnd.n6584 9.3005
R10316 gnd.n714 gnd.n713 9.3005
R10317 gnd.n6592 gnd.n6591 9.3005
R10318 gnd.n6593 gnd.n712 9.3005
R10319 gnd.n6595 gnd.n6594 9.3005
R10320 gnd.n708 gnd.n707 9.3005
R10321 gnd.n6602 gnd.n6601 9.3005
R10322 gnd.n6603 gnd.n706 9.3005
R10323 gnd.n6605 gnd.n6604 9.3005
R10324 gnd.n702 gnd.n701 9.3005
R10325 gnd.n6612 gnd.n6611 9.3005
R10326 gnd.n6613 gnd.n700 9.3005
R10327 gnd.n6615 gnd.n6614 9.3005
R10328 gnd.n696 gnd.n695 9.3005
R10329 gnd.n6622 gnd.n6621 9.3005
R10330 gnd.n6623 gnd.n694 9.3005
R10331 gnd.n6626 gnd.n6625 9.3005
R10332 gnd.n6624 gnd.n690 9.3005
R10333 gnd.n6632 gnd.n689 9.3005
R10334 gnd.n6634 gnd.n6633 9.3005
R10335 gnd.n685 gnd.n684 9.3005
R10336 gnd.n6643 gnd.n6642 9.3005
R10337 gnd.n6644 gnd.n683 9.3005
R10338 gnd.n6646 gnd.n6645 9.3005
R10339 gnd.n679 gnd.n678 9.3005
R10340 gnd.n6653 gnd.n6652 9.3005
R10341 gnd.n6654 gnd.n677 9.3005
R10342 gnd.n6656 gnd.n6655 9.3005
R10343 gnd.n673 gnd.n672 9.3005
R10344 gnd.n6663 gnd.n6662 9.3005
R10345 gnd.n6664 gnd.n671 9.3005
R10346 gnd.n6666 gnd.n6665 9.3005
R10347 gnd.n667 gnd.n666 9.3005
R10348 gnd.n6673 gnd.n6672 9.3005
R10349 gnd.n6674 gnd.n665 9.3005
R10350 gnd.n6676 gnd.n6675 9.3005
R10351 gnd.n661 gnd.n660 9.3005
R10352 gnd.n6683 gnd.n6682 9.3005
R10353 gnd.n6684 gnd.n659 9.3005
R10354 gnd.n6686 gnd.n6685 9.3005
R10355 gnd.n655 gnd.n654 9.3005
R10356 gnd.n6693 gnd.n6692 9.3005
R10357 gnd.n6694 gnd.n653 9.3005
R10358 gnd.n6696 gnd.n6695 9.3005
R10359 gnd.n649 gnd.n648 9.3005
R10360 gnd.n6703 gnd.n6702 9.3005
R10361 gnd.n6704 gnd.n647 9.3005
R10362 gnd.n6706 gnd.n6705 9.3005
R10363 gnd.n643 gnd.n642 9.3005
R10364 gnd.n6713 gnd.n6712 9.3005
R10365 gnd.n6714 gnd.n641 9.3005
R10366 gnd.n6716 gnd.n6715 9.3005
R10367 gnd.n637 gnd.n636 9.3005
R10368 gnd.n6723 gnd.n6722 9.3005
R10369 gnd.n6724 gnd.n635 9.3005
R10370 gnd.n6726 gnd.n6725 9.3005
R10371 gnd.n631 gnd.n630 9.3005
R10372 gnd.n6733 gnd.n6732 9.3005
R10373 gnd.n6734 gnd.n629 9.3005
R10374 gnd.n6736 gnd.n6735 9.3005
R10375 gnd.n625 gnd.n624 9.3005
R10376 gnd.n6743 gnd.n6742 9.3005
R10377 gnd.n6744 gnd.n623 9.3005
R10378 gnd.n6746 gnd.n6745 9.3005
R10379 gnd.n619 gnd.n618 9.3005
R10380 gnd.n6753 gnd.n6752 9.3005
R10381 gnd.n6754 gnd.n617 9.3005
R10382 gnd.n6756 gnd.n6755 9.3005
R10383 gnd.n613 gnd.n612 9.3005
R10384 gnd.n6763 gnd.n6762 9.3005
R10385 gnd.n6764 gnd.n611 9.3005
R10386 gnd.n6766 gnd.n6765 9.3005
R10387 gnd.n607 gnd.n606 9.3005
R10388 gnd.n6773 gnd.n6772 9.3005
R10389 gnd.n6774 gnd.n605 9.3005
R10390 gnd.n6776 gnd.n6775 9.3005
R10391 gnd.n601 gnd.n600 9.3005
R10392 gnd.n6783 gnd.n6782 9.3005
R10393 gnd.n6784 gnd.n599 9.3005
R10394 gnd.n6786 gnd.n6785 9.3005
R10395 gnd.n595 gnd.n594 9.3005
R10396 gnd.n6793 gnd.n6792 9.3005
R10397 gnd.n6794 gnd.n593 9.3005
R10398 gnd.n6796 gnd.n6795 9.3005
R10399 gnd.n589 gnd.n588 9.3005
R10400 gnd.n6803 gnd.n6802 9.3005
R10401 gnd.n6804 gnd.n587 9.3005
R10402 gnd.n6806 gnd.n6805 9.3005
R10403 gnd.n583 gnd.n582 9.3005
R10404 gnd.n6813 gnd.n6812 9.3005
R10405 gnd.n6814 gnd.n581 9.3005
R10406 gnd.n6816 gnd.n6815 9.3005
R10407 gnd.n577 gnd.n576 9.3005
R10408 gnd.n6823 gnd.n6822 9.3005
R10409 gnd.n6824 gnd.n575 9.3005
R10410 gnd.n6826 gnd.n6825 9.3005
R10411 gnd.n571 gnd.n570 9.3005
R10412 gnd.n6833 gnd.n6832 9.3005
R10413 gnd.n6834 gnd.n569 9.3005
R10414 gnd.n6836 gnd.n6835 9.3005
R10415 gnd.n565 gnd.n564 9.3005
R10416 gnd.n6844 gnd.n6843 9.3005
R10417 gnd.n6845 gnd.n563 9.3005
R10418 gnd.n6847 gnd.n6846 9.3005
R10419 gnd.n6636 gnd.n6635 9.3005
R10420 gnd.n7029 gnd.n7028 9.3005
R10421 gnd.n7027 gnd.n65 9.3005
R10422 gnd.n214 gnd.n67 9.3005
R10423 gnd.n217 gnd.n215 9.3005
R10424 gnd.n219 gnd.n218 9.3005
R10425 gnd.n220 gnd.n213 9.3005
R10426 gnd.n222 gnd.n221 9.3005
R10427 gnd.n224 gnd.n211 9.3005
R10428 gnd.n226 gnd.n225 9.3005
R10429 gnd.n227 gnd.n210 9.3005
R10430 gnd.n229 gnd.n228 9.3005
R10431 gnd.n231 gnd.n208 9.3005
R10432 gnd.n233 gnd.n232 9.3005
R10433 gnd.n234 gnd.n207 9.3005
R10434 gnd.n236 gnd.n235 9.3005
R10435 gnd.n238 gnd.n205 9.3005
R10436 gnd.n240 gnd.n239 9.3005
R10437 gnd.n241 gnd.n204 9.3005
R10438 gnd.n243 gnd.n242 9.3005
R10439 gnd.n245 gnd.n202 9.3005
R10440 gnd.n247 gnd.n246 9.3005
R10441 gnd.n278 gnd.n168 9.3005
R10442 gnd.n277 gnd.n170 9.3005
R10443 gnd.n174 gnd.n171 9.3005
R10444 gnd.n272 gnd.n175 9.3005
R10445 gnd.n271 gnd.n176 9.3005
R10446 gnd.n270 gnd.n177 9.3005
R10447 gnd.n181 gnd.n178 9.3005
R10448 gnd.n265 gnd.n182 9.3005
R10449 gnd.n264 gnd.n183 9.3005
R10450 gnd.n263 gnd.n184 9.3005
R10451 gnd.n188 gnd.n185 9.3005
R10452 gnd.n258 gnd.n189 9.3005
R10453 gnd.n257 gnd.n190 9.3005
R10454 gnd.n256 gnd.n191 9.3005
R10455 gnd.n195 gnd.n192 9.3005
R10456 gnd.n251 gnd.n196 9.3005
R10457 gnd.n250 gnd.n249 9.3005
R10458 gnd.n248 gnd.n199 9.3005
R10459 gnd.n280 gnd.n279 9.3005
R10460 gnd.n346 gnd.n343 9.3005
R10461 gnd.n352 gnd.n351 9.3005
R10462 gnd.n353 gnd.n342 9.3005
R10463 gnd.n355 gnd.n354 9.3005
R10464 gnd.n340 gnd.n339 9.3005
R10465 gnd.n362 gnd.n361 9.3005
R10466 gnd.n363 gnd.n338 9.3005
R10467 gnd.n365 gnd.n364 9.3005
R10468 gnd.n336 gnd.n335 9.3005
R10469 gnd.n372 gnd.n371 9.3005
R10470 gnd.n373 gnd.n334 9.3005
R10471 gnd.n375 gnd.n374 9.3005
R10472 gnd.n332 gnd.n331 9.3005
R10473 gnd.n383 gnd.n382 9.3005
R10474 gnd.n384 gnd.n330 9.3005
R10475 gnd.n386 gnd.n385 9.3005
R10476 gnd.n387 gnd.n325 9.3005
R10477 gnd.n393 gnd.n392 9.3005
R10478 gnd.n394 gnd.n324 9.3005
R10479 gnd.n396 gnd.n395 9.3005
R10480 gnd.n322 gnd.n321 9.3005
R10481 gnd.n403 gnd.n402 9.3005
R10482 gnd.n404 gnd.n320 9.3005
R10483 gnd.n406 gnd.n405 9.3005
R10484 gnd.n318 gnd.n317 9.3005
R10485 gnd.n413 gnd.n412 9.3005
R10486 gnd.n414 gnd.n316 9.3005
R10487 gnd.n416 gnd.n415 9.3005
R10488 gnd.n314 gnd.n313 9.3005
R10489 gnd.n423 gnd.n422 9.3005
R10490 gnd.n424 gnd.n312 9.3005
R10491 gnd.n426 gnd.n425 9.3005
R10492 gnd.n310 gnd.n309 9.3005
R10493 gnd.n433 gnd.n432 9.3005
R10494 gnd.n434 gnd.n308 9.3005
R10495 gnd.n436 gnd.n435 9.3005
R10496 gnd.n306 gnd.n303 9.3005
R10497 gnd.n443 gnd.n442 9.3005
R10498 gnd.n444 gnd.n302 9.3005
R10499 gnd.n446 gnd.n445 9.3005
R10500 gnd.n300 gnd.n299 9.3005
R10501 gnd.n453 gnd.n452 9.3005
R10502 gnd.n454 gnd.n298 9.3005
R10503 gnd.n456 gnd.n455 9.3005
R10504 gnd.n296 gnd.n295 9.3005
R10505 gnd.n463 gnd.n462 9.3005
R10506 gnd.n464 gnd.n294 9.3005
R10507 gnd.n466 gnd.n465 9.3005
R10508 gnd.n292 gnd.n291 9.3005
R10509 gnd.n473 gnd.n472 9.3005
R10510 gnd.n474 gnd.n290 9.3005
R10511 gnd.n476 gnd.n475 9.3005
R10512 gnd.n288 gnd.n287 9.3005
R10513 gnd.n483 gnd.n482 9.3005
R10514 gnd.n484 gnd.n286 9.3005
R10515 gnd.n486 gnd.n485 9.3005
R10516 gnd.n284 gnd.n281 9.3005
R10517 gnd.n492 gnd.n491 9.3005
R10518 gnd.n345 gnd.n344 9.3005
R10519 gnd.n5631 gnd.n5630 9.3005
R10520 gnd.n1674 gnd.n1673 9.3005
R10521 gnd.n1698 gnd.n1697 9.3005
R10522 gnd.n5618 gnd.n1699 9.3005
R10523 gnd.n5617 gnd.n1700 9.3005
R10524 gnd.n5616 gnd.n1701 9.3005
R10525 gnd.n5547 gnd.n1702 9.3005
R10526 gnd.n5606 gnd.n1721 9.3005
R10527 gnd.n5605 gnd.n5604 9.3005
R10528 gnd.n1722 gnd.n552 9.3005
R10529 gnd.n6862 gnd.n553 9.3005
R10530 gnd.n6861 gnd.n554 9.3005
R10531 gnd.n6860 gnd.n555 9.3005
R10532 gnd.n6859 gnd.n556 9.3005
R10533 gnd.n529 gnd.n525 9.3005
R10534 gnd.n6895 gnd.n526 9.3005
R10535 gnd.n6894 gnd.n527 9.3005
R10536 gnd.n6893 gnd.n6891 9.3005
R10537 gnd.n503 gnd.n502 9.3005
R10538 gnd.n6921 gnd.n6920 9.3005
R10539 gnd.n6922 gnd.n496 9.3005
R10540 gnd.n6929 gnd.n497 9.3005
R10541 gnd.n6930 gnd.n495 9.3005
R10542 gnd.n6933 gnd.n6932 9.3005
R10543 gnd.n6934 gnd.n91 9.3005
R10544 gnd.n7015 gnd.n92 9.3005
R10545 gnd.n7014 gnd.n93 9.3005
R10546 gnd.n7013 gnd.n94 9.3005
R10547 gnd.n6942 gnd.n95 9.3005
R10548 gnd.n7003 gnd.n109 9.3005
R10549 gnd.n7002 gnd.n110 9.3005
R10550 gnd.n7001 gnd.n111 9.3005
R10551 gnd.n6949 gnd.n112 9.3005
R10552 gnd.n6991 gnd.n129 9.3005
R10553 gnd.n6990 gnd.n130 9.3005
R10554 gnd.n6989 gnd.n131 9.3005
R10555 gnd.n6956 gnd.n132 9.3005
R10556 gnd.n6979 gnd.n149 9.3005
R10557 gnd.n6978 gnd.n150 9.3005
R10558 gnd.n6977 gnd.n151 9.3005
R10559 gnd.n167 gnd.n152 9.3005
R10560 gnd.n6967 gnd.n6966 9.3005
R10561 gnd.n5632 gnd.n1672 9.3005
R10562 gnd.n5630 gnd.n5629 9.3005
R10563 gnd.n5628 gnd.n1674 9.3005
R10564 gnd.n1698 gnd.n1675 9.3005
R10565 gnd.n5542 gnd.n1699 9.3005
R10566 gnd.n5545 gnd.n1700 9.3005
R10567 gnd.n5546 gnd.n1701 9.3005
R10568 gnd.n5548 gnd.n5547 9.3005
R10569 gnd.n1723 gnd.n1721 9.3005
R10570 gnd.n5604 gnd.n5603 9.3005
R10571 gnd.n1729 gnd.n1722 9.3005
R10572 gnd.n1728 gnd.n553 9.3005
R10573 gnd.n1727 gnd.n554 9.3005
R10574 gnd.n1724 gnd.n555 9.3005
R10575 gnd.n556 gnd.n528 9.3005
R10576 gnd.n6885 gnd.n529 9.3005
R10577 gnd.n6886 gnd.n526 9.3005
R10578 gnd.n6887 gnd.n527 9.3005
R10579 gnd.n6891 gnd.n6890 9.3005
R10580 gnd.n6888 gnd.n502 9.3005
R10581 gnd.n6921 gnd.n501 9.3005
R10582 gnd.n6923 gnd.n6922 9.3005
R10583 gnd.n6925 gnd.n497 9.3005
R10584 gnd.n6924 gnd.n495 9.3005
R10585 gnd.n6933 gnd.n494 9.3005
R10586 gnd.n6937 gnd.n6934 9.3005
R10587 gnd.n6938 gnd.n92 9.3005
R10588 gnd.n6940 gnd.n93 9.3005
R10589 gnd.n6941 gnd.n94 9.3005
R10590 gnd.n6944 gnd.n6942 9.3005
R10591 gnd.n6945 gnd.n109 9.3005
R10592 gnd.n6947 gnd.n110 9.3005
R10593 gnd.n6948 gnd.n111 9.3005
R10594 gnd.n6951 gnd.n6949 9.3005
R10595 gnd.n6952 gnd.n129 9.3005
R10596 gnd.n6954 gnd.n130 9.3005
R10597 gnd.n6955 gnd.n131 9.3005
R10598 gnd.n6958 gnd.n6956 9.3005
R10599 gnd.n6959 gnd.n149 9.3005
R10600 gnd.n6961 gnd.n150 9.3005
R10601 gnd.n6962 gnd.n151 9.3005
R10602 gnd.n6964 gnd.n167 9.3005
R10603 gnd.n6966 gnd.n6965 9.3005
R10604 gnd.n1672 gnd.n1666 9.3005
R10605 gnd.n5642 gnd.n5641 9.3005
R10606 gnd.n5645 gnd.n1664 9.3005
R10607 gnd.n5646 gnd.n1663 9.3005
R10608 gnd.n5649 gnd.n1662 9.3005
R10609 gnd.n5650 gnd.n1661 9.3005
R10610 gnd.n5653 gnd.n1660 9.3005
R10611 gnd.n5654 gnd.n1659 9.3005
R10612 gnd.n5657 gnd.n1658 9.3005
R10613 gnd.n5658 gnd.n1657 9.3005
R10614 gnd.n5661 gnd.n1656 9.3005
R10615 gnd.n5662 gnd.n1655 9.3005
R10616 gnd.n5665 gnd.n1654 9.3005
R10617 gnd.n5666 gnd.n1653 9.3005
R10618 gnd.n5669 gnd.n1652 9.3005
R10619 gnd.n5670 gnd.n1651 9.3005
R10620 gnd.n5673 gnd.n1650 9.3005
R10621 gnd.n5674 gnd.n1649 9.3005
R10622 gnd.n5677 gnd.n1648 9.3005
R10623 gnd.n5678 gnd.n1647 9.3005
R10624 gnd.n5681 gnd.n1646 9.3005
R10625 gnd.n5685 gnd.n1642 9.3005
R10626 gnd.n5686 gnd.n1641 9.3005
R10627 gnd.n5689 gnd.n1640 9.3005
R10628 gnd.n5690 gnd.n1639 9.3005
R10629 gnd.n5693 gnd.n1638 9.3005
R10630 gnd.n5694 gnd.n1637 9.3005
R10631 gnd.n5697 gnd.n1636 9.3005
R10632 gnd.n5698 gnd.n1635 9.3005
R10633 gnd.n5701 gnd.n1634 9.3005
R10634 gnd.n5703 gnd.n1630 9.3005
R10635 gnd.n5706 gnd.n1629 9.3005
R10636 gnd.n5707 gnd.n1628 9.3005
R10637 gnd.n5710 gnd.n1627 9.3005
R10638 gnd.n5711 gnd.n1626 9.3005
R10639 gnd.n5714 gnd.n1625 9.3005
R10640 gnd.n5715 gnd.n1624 9.3005
R10641 gnd.n5718 gnd.n1623 9.3005
R10642 gnd.n5720 gnd.n1620 9.3005
R10643 gnd.n5723 gnd.n1619 9.3005
R10644 gnd.n5724 gnd.n1618 9.3005
R10645 gnd.n5727 gnd.n1617 9.3005
R10646 gnd.n5728 gnd.n1616 9.3005
R10647 gnd.n5731 gnd.n1615 9.3005
R10648 gnd.n5732 gnd.n1614 9.3005
R10649 gnd.n5735 gnd.n1613 9.3005
R10650 gnd.n5736 gnd.n1612 9.3005
R10651 gnd.n5739 gnd.n1611 9.3005
R10652 gnd.n5740 gnd.n1610 9.3005
R10653 gnd.n5743 gnd.n1609 9.3005
R10654 gnd.n5744 gnd.n1608 9.3005
R10655 gnd.n5747 gnd.n1607 9.3005
R10656 gnd.n5749 gnd.n1606 9.3005
R10657 gnd.n5750 gnd.n1605 9.3005
R10658 gnd.n5751 gnd.n1604 9.3005
R10659 gnd.n5752 gnd.n1603 9.3005
R10660 gnd.n5682 gnd.n1643 9.3005
R10661 gnd.n5640 gnd.n5637 9.3005
R10662 gnd.n1685 gnd.n1682 9.3005
R10663 gnd.n5624 gnd.n1686 9.3005
R10664 gnd.n5623 gnd.n1687 9.3005
R10665 gnd.n5622 gnd.n1688 9.3005
R10666 gnd.n1709 gnd.n1689 9.3005
R10667 gnd.n5612 gnd.n1710 9.3005
R10668 gnd.n5611 gnd.n1711 9.3005
R10669 gnd.n5610 gnd.n1712 9.3005
R10670 gnd.n1714 gnd.n1713 9.3005
R10671 gnd.n544 gnd.n543 9.3005
R10672 gnd.n6867 gnd.n6866 9.3005
R10673 gnd.n6868 gnd.n542 9.3005
R10674 gnd.n6873 gnd.n6869 9.3005
R10675 gnd.n6872 gnd.n6870 9.3005
R10676 gnd.n6871 gnd.n77 9.3005
R10677 gnd.n82 gnd.n76 9.3005
R10678 gnd.n7009 gnd.n101 9.3005
R10679 gnd.n7008 gnd.n102 9.3005
R10680 gnd.n7007 gnd.n103 9.3005
R10681 gnd.n118 gnd.n104 9.3005
R10682 gnd.n6997 gnd.n119 9.3005
R10683 gnd.n6996 gnd.n120 9.3005
R10684 gnd.n6995 gnd.n121 9.3005
R10685 gnd.n138 gnd.n122 9.3005
R10686 gnd.n6985 gnd.n139 9.3005
R10687 gnd.n6984 gnd.n140 9.3005
R10688 gnd.n6983 gnd.n141 9.3005
R10689 gnd.n157 gnd.n142 9.3005
R10690 gnd.n6973 gnd.n158 9.3005
R10691 gnd.n6972 gnd.n159 9.3005
R10692 gnd.n6971 gnd.n160 9.3005
R10693 gnd.n1684 gnd.n1683 9.3005
R10694 gnd.n7020 gnd.n7019 9.3005
R10695 gnd.n6852 gnd.n6851 9.3005
R10696 gnd.n4404 gnd.n4403 9.3005
R10697 gnd.n4405 gnd.n4398 9.3005
R10698 gnd.n4407 gnd.n4406 9.3005
R10699 gnd.n2323 gnd.n2322 9.3005
R10700 gnd.n4412 gnd.n4411 9.3005
R10701 gnd.n4413 gnd.n2321 9.3005
R10702 gnd.n4419 gnd.n4414 9.3005
R10703 gnd.n4418 gnd.n4415 9.3005
R10704 gnd.n4417 gnd.n4416 9.3005
R10705 gnd.n2305 gnd.n2304 9.3005
R10706 gnd.n4695 gnd.n4694 9.3005
R10707 gnd.n4696 gnd.n2303 9.3005
R10708 gnd.n4698 gnd.n4697 9.3005
R10709 gnd.n2301 gnd.n2300 9.3005
R10710 gnd.n4703 gnd.n4702 9.3005
R10711 gnd.n4704 gnd.n2299 9.3005
R10712 gnd.n4711 gnd.n4705 9.3005
R10713 gnd.n4710 gnd.n4706 9.3005
R10714 gnd.n4709 gnd.n4707 9.3005
R10715 gnd.n2271 gnd.n2270 9.3005
R10716 gnd.n4741 gnd.n4740 9.3005
R10717 gnd.n4742 gnd.n2269 9.3005
R10718 gnd.n4753 gnd.n4743 9.3005
R10719 gnd.n4752 gnd.n4744 9.3005
R10720 gnd.n4751 gnd.n4745 9.3005
R10721 gnd.n4748 gnd.n4747 9.3005
R10722 gnd.n4746 gnd.n1284 9.3005
R10723 gnd.n5956 gnd.n1285 9.3005
R10724 gnd.n5955 gnd.n1286 9.3005
R10725 gnd.n5954 gnd.n1287 9.3005
R10726 gnd.n1385 gnd.n1288 9.3005
R10727 gnd.n1386 gnd.n1384 9.3005
R10728 gnd.n5937 gnd.n1387 9.3005
R10729 gnd.n5936 gnd.n1388 9.3005
R10730 gnd.n5935 gnd.n1389 9.3005
R10731 gnd.n4840 gnd.n1390 9.3005
R10732 gnd.n4841 gnd.n4839 9.3005
R10733 gnd.n4843 gnd.n4842 9.3005
R10734 gnd.n2227 gnd.n2226 9.3005
R10735 gnd.n4882 gnd.n4881 9.3005
R10736 gnd.n4883 gnd.n2225 9.3005
R10737 gnd.n4886 gnd.n4885 9.3005
R10738 gnd.n4884 gnd.n2195 9.3005
R10739 gnd.n4938 gnd.n2196 9.3005
R10740 gnd.n4937 gnd.n2197 9.3005
R10741 gnd.n4936 gnd.n2198 9.3005
R10742 gnd.n2201 gnd.n2199 9.3005
R10743 gnd.n2211 gnd.n2202 9.3005
R10744 gnd.n2210 gnd.n2203 9.3005
R10745 gnd.n2209 gnd.n2204 9.3005
R10746 gnd.n2206 gnd.n2205 9.3005
R10747 gnd.n2154 gnd.n2153 9.3005
R10748 gnd.n4997 gnd.n4996 9.3005
R10749 gnd.n4998 gnd.n2152 9.3005
R10750 gnd.n5002 gnd.n4999 9.3005
R10751 gnd.n5001 gnd.n5000 9.3005
R10752 gnd.n2128 gnd.n2127 9.3005
R10753 gnd.n5053 gnd.n5052 9.3005
R10754 gnd.n5054 gnd.n2126 9.3005
R10755 gnd.n5058 gnd.n5055 9.3005
R10756 gnd.n5057 gnd.n5056 9.3005
R10757 gnd.n2106 gnd.n2105 9.3005
R10758 gnd.n5100 gnd.n5099 9.3005
R10759 gnd.n5101 gnd.n2104 9.3005
R10760 gnd.n5103 gnd.n5102 9.3005
R10761 gnd.n2082 gnd.n2081 9.3005
R10762 gnd.n5130 gnd.n5129 9.3005
R10763 gnd.n5131 gnd.n2080 9.3005
R10764 gnd.n5133 gnd.n5132 9.3005
R10765 gnd.n2064 gnd.n2063 9.3005
R10766 gnd.n5178 gnd.n5177 9.3005
R10767 gnd.n5179 gnd.n2062 9.3005
R10768 gnd.n5183 gnd.n5180 9.3005
R10769 gnd.n5182 gnd.n5181 9.3005
R10770 gnd.n2038 gnd.n2037 9.3005
R10771 gnd.n5214 gnd.n5213 9.3005
R10772 gnd.n5215 gnd.n2036 9.3005
R10773 gnd.n5219 gnd.n5216 9.3005
R10774 gnd.n5218 gnd.n5217 9.3005
R10775 gnd.n2008 gnd.n2007 9.3005
R10776 gnd.n5278 gnd.n5277 9.3005
R10777 gnd.n5279 gnd.n2006 9.3005
R10778 gnd.n5281 gnd.n5280 9.3005
R10779 gnd.n1991 gnd.n1990 9.3005
R10780 gnd.n5307 gnd.n5306 9.3005
R10781 gnd.n5308 gnd.n1989 9.3005
R10782 gnd.n5312 gnd.n5309 9.3005
R10783 gnd.n5311 gnd.n5310 9.3005
R10784 gnd.n1965 gnd.n1964 9.3005
R10785 gnd.n5343 gnd.n5342 9.3005
R10786 gnd.n5344 gnd.n1963 9.3005
R10787 gnd.n5346 gnd.n5345 9.3005
R10788 gnd.n1937 gnd.n1936 9.3005
R10789 gnd.n5380 gnd.n5379 9.3005
R10790 gnd.n5381 gnd.n1935 9.3005
R10791 gnd.n5385 gnd.n5382 9.3005
R10792 gnd.n5384 gnd.n5383 9.3005
R10793 gnd.n1788 gnd.n1787 9.3005
R10794 gnd.n5488 gnd.n5487 9.3005
R10795 gnd.n5489 gnd.n1786 9.3005
R10796 gnd.n5494 gnd.n5490 9.3005
R10797 gnd.n5493 gnd.n5492 9.3005
R10798 gnd.n5491 gnd.n1777 9.3005
R10799 gnd.n5507 gnd.n1776 9.3005
R10800 gnd.n5509 gnd.n5508 9.3005
R10801 gnd.n5510 gnd.n1775 9.3005
R10802 gnd.n5526 gnd.n5511 9.3005
R10803 gnd.n5525 gnd.n5512 9.3005
R10804 gnd.n5524 gnd.n5513 9.3005
R10805 gnd.n5515 gnd.n5514 9.3005
R10806 gnd.n5520 gnd.n5516 9.3005
R10807 gnd.n5519 gnd.n5518 9.3005
R10808 gnd.n5517 gnd.n1743 9.3005
R10809 gnd.n1741 gnd.n1740 9.3005
R10810 gnd.n5578 gnd.n5577 9.3005
R10811 gnd.n5579 gnd.n1739 9.3005
R10812 gnd.n5581 gnd.n5580 9.3005
R10813 gnd.n1737 gnd.n1736 9.3005
R10814 gnd.n5586 gnd.n5585 9.3005
R10815 gnd.n5587 gnd.n1735 9.3005
R10816 gnd.n5598 gnd.n5588 9.3005
R10817 gnd.n5597 gnd.n5589 9.3005
R10818 gnd.n5596 gnd.n5590 9.3005
R10819 gnd.n5593 gnd.n5592 9.3005
R10820 gnd.n5591 gnd.n559 9.3005
R10821 gnd.n6854 gnd.n560 9.3005
R10822 gnd.n6853 gnd.n561 9.3005
R10823 gnd.n4050 gnd.n4049 9.3005
R10824 gnd.n4080 gnd.n4027 9.3005
R10825 gnd.n4079 gnd.n4028 9.3005
R10826 gnd.n4077 gnd.n4029 9.3005
R10827 gnd.n4076 gnd.n4030 9.3005
R10828 gnd.n4074 gnd.n4031 9.3005
R10829 gnd.n4073 gnd.n4032 9.3005
R10830 gnd.n4071 gnd.n4033 9.3005
R10831 gnd.n4070 gnd.n4034 9.3005
R10832 gnd.n4068 gnd.n4035 9.3005
R10833 gnd.n4067 gnd.n4036 9.3005
R10834 gnd.n4065 gnd.n4037 9.3005
R10835 gnd.n4064 gnd.n4038 9.3005
R10836 gnd.n4062 gnd.n4039 9.3005
R10837 gnd.n4061 gnd.n4040 9.3005
R10838 gnd.n4059 gnd.n4041 9.3005
R10839 gnd.n4058 gnd.n4042 9.3005
R10840 gnd.n4056 gnd.n4043 9.3005
R10841 gnd.n4055 gnd.n4044 9.3005
R10842 gnd.n4053 gnd.n4045 9.3005
R10843 gnd.n4052 gnd.n4046 9.3005
R10844 gnd.n4083 gnd.n4082 9.3005
R10845 gnd.n4088 gnd.n4087 9.3005
R10846 gnd.n4091 gnd.n4022 9.3005
R10847 gnd.n4092 gnd.n4021 9.3005
R10848 gnd.n4095 gnd.n4020 9.3005
R10849 gnd.n4096 gnd.n4019 9.3005
R10850 gnd.n4099 gnd.n4018 9.3005
R10851 gnd.n4100 gnd.n4017 9.3005
R10852 gnd.n4103 gnd.n4016 9.3005
R10853 gnd.n4104 gnd.n4015 9.3005
R10854 gnd.n4107 gnd.n4014 9.3005
R10855 gnd.n4108 gnd.n4013 9.3005
R10856 gnd.n4111 gnd.n4012 9.3005
R10857 gnd.n4112 gnd.n4011 9.3005
R10858 gnd.n4115 gnd.n4010 9.3005
R10859 gnd.n4116 gnd.n4009 9.3005
R10860 gnd.n4119 gnd.n4008 9.3005
R10861 gnd.n4122 gnd.n4121 9.3005
R10862 gnd.n4086 gnd.n4026 9.3005
R10863 gnd.n4085 gnd.n4084 9.3005
R10864 gnd.n6035 gnd.n1210 9.3005
R10865 gnd.n6038 gnd.n1209 9.3005
R10866 gnd.n6039 gnd.n1208 9.3005
R10867 gnd.n6042 gnd.n1207 9.3005
R10868 gnd.n6043 gnd.n1206 9.3005
R10869 gnd.n6046 gnd.n1205 9.3005
R10870 gnd.n6047 gnd.n1204 9.3005
R10871 gnd.n6050 gnd.n1203 9.3005
R10872 gnd.n6052 gnd.n1200 9.3005
R10873 gnd.n6055 gnd.n1199 9.3005
R10874 gnd.n6056 gnd.n1198 9.3005
R10875 gnd.n6059 gnd.n1197 9.3005
R10876 gnd.n6060 gnd.n1196 9.3005
R10877 gnd.n6063 gnd.n1195 9.3005
R10878 gnd.n6064 gnd.n1194 9.3005
R10879 gnd.n6067 gnd.n1193 9.3005
R10880 gnd.n6068 gnd.n1192 9.3005
R10881 gnd.n6071 gnd.n1191 9.3005
R10882 gnd.n6072 gnd.n1190 9.3005
R10883 gnd.n6075 gnd.n1189 9.3005
R10884 gnd.n6076 gnd.n1188 9.3005
R10885 gnd.n6079 gnd.n1187 9.3005
R10886 gnd.n6080 gnd.n1186 9.3005
R10887 gnd.n6081 gnd.n1185 9.3005
R10888 gnd.n1142 gnd.n1141 9.3005
R10889 gnd.n6087 gnd.n6086 9.3005
R10890 gnd.n4599 gnd.n4596 9.3005
R10891 gnd.n4603 gnd.n4602 9.3005
R10892 gnd.n4604 gnd.n4594 9.3005
R10893 gnd.n4606 gnd.n4605 9.3005
R10894 gnd.n4609 gnd.n4593 9.3005
R10895 gnd.n4613 gnd.n4612 9.3005
R10896 gnd.n4614 gnd.n4592 9.3005
R10897 gnd.n4617 gnd.n4615 9.3005
R10898 gnd.n4618 gnd.n4588 9.3005
R10899 gnd.n4622 gnd.n4621 9.3005
R10900 gnd.n4623 gnd.n4587 9.3005
R10901 gnd.n4625 gnd.n4624 9.3005
R10902 gnd.n4628 gnd.n4586 9.3005
R10903 gnd.n4632 gnd.n4631 9.3005
R10904 gnd.n4633 gnd.n4585 9.3005
R10905 gnd.n4635 gnd.n4634 9.3005
R10906 gnd.n4638 gnd.n4584 9.3005
R10907 gnd.n4642 gnd.n4641 9.3005
R10908 gnd.n4643 gnd.n4583 9.3005
R10909 gnd.n4645 gnd.n4644 9.3005
R10910 gnd.n4648 gnd.n4582 9.3005
R10911 gnd.n4652 gnd.n4651 9.3005
R10912 gnd.n4653 gnd.n4581 9.3005
R10913 gnd.n4655 gnd.n4654 9.3005
R10914 gnd.n4658 gnd.n4580 9.3005
R10915 gnd.n4662 gnd.n4661 9.3005
R10916 gnd.n4663 gnd.n4579 9.3005
R10917 gnd.n4666 gnd.n4664 9.3005
R10918 gnd.n4667 gnd.n4575 9.3005
R10919 gnd.n4670 gnd.n4669 9.3005
R10920 gnd.n4595 gnd.n1211 9.3005
R10921 gnd.n4249 gnd.n4248 9.3005
R10922 gnd.n2440 gnd.n2436 9.3005
R10923 gnd.n2439 gnd.n2438 9.3005
R10924 gnd.n2420 gnd.n2417 9.3005
R10925 gnd.n4269 gnd.n2418 9.3005
R10926 gnd.n4268 gnd.n4265 9.3005
R10927 gnd.n4267 gnd.n4266 9.3005
R10928 gnd.n2402 gnd.n2399 9.3005
R10929 gnd.n4289 gnd.n2400 9.3005
R10930 gnd.n4288 gnd.n4285 9.3005
R10931 gnd.n4287 gnd.n4286 9.3005
R10932 gnd.n2384 gnd.n2381 9.3005
R10933 gnd.n4309 gnd.n2382 9.3005
R10934 gnd.n4308 gnd.n4305 9.3005
R10935 gnd.n4307 gnd.n4306 9.3005
R10936 gnd.n2366 gnd.n2363 9.3005
R10937 gnd.n4330 gnd.n2364 9.3005
R10938 gnd.n4329 gnd.n4326 9.3005
R10939 gnd.n4328 gnd.n4327 9.3005
R10940 gnd.n2350 gnd.n2345 9.3005
R10941 gnd.n4357 gnd.n2346 9.3005
R10942 gnd.n4356 gnd.n2347 9.3005
R10943 gnd.n4355 gnd.n2348 9.3005
R10944 gnd.n4354 gnd.n4350 9.3005
R10945 gnd.n4352 gnd.n4351 9.3005
R10946 gnd.n2329 gnd.n1067 9.3005
R10947 gnd.n6132 gnd.n1068 9.3005
R10948 gnd.n6131 gnd.n1069 9.3005
R10949 gnd.n6130 gnd.n1070 9.3005
R10950 gnd.n4382 gnd.n1071 9.3005
R10951 gnd.n6120 gnd.n1089 9.3005
R10952 gnd.n6119 gnd.n1090 9.3005
R10953 gnd.n6118 gnd.n1091 9.3005
R10954 gnd.n2314 gnd.n1092 9.3005
R10955 gnd.n6108 gnd.n1108 9.3005
R10956 gnd.n6107 gnd.n1109 9.3005
R10957 gnd.n6106 gnd.n1110 9.3005
R10958 gnd.n4436 gnd.n1111 9.3005
R10959 gnd.n6096 gnd.n1129 9.3005
R10960 gnd.n6095 gnd.n1130 9.3005
R10961 gnd.n6094 gnd.n1131 9.3005
R10962 gnd.n4672 gnd.n1132 9.3005
R10963 gnd.n2437 gnd.n2435 9.3005
R10964 gnd.n4248 gnd.n4247 9.3005
R10965 gnd.n4246 gnd.n2440 9.3005
R10966 gnd.n2439 gnd.n2419 9.3005
R10967 gnd.n4262 gnd.n2420 9.3005
R10968 gnd.n4263 gnd.n2418 9.3005
R10969 gnd.n4265 gnd.n4264 9.3005
R10970 gnd.n4266 gnd.n2401 9.3005
R10971 gnd.n4282 gnd.n2402 9.3005
R10972 gnd.n4283 gnd.n2400 9.3005
R10973 gnd.n4285 gnd.n4284 9.3005
R10974 gnd.n4286 gnd.n2383 9.3005
R10975 gnd.n4302 gnd.n2384 9.3005
R10976 gnd.n4303 gnd.n2382 9.3005
R10977 gnd.n4305 gnd.n4304 9.3005
R10978 gnd.n4306 gnd.n2365 9.3005
R10979 gnd.n4323 gnd.n2366 9.3005
R10980 gnd.n4324 gnd.n2364 9.3005
R10981 gnd.n4326 gnd.n4325 9.3005
R10982 gnd.n4327 gnd.n2349 9.3005
R10983 gnd.n4343 gnd.n2350 9.3005
R10984 gnd.n4344 gnd.n2346 9.3005
R10985 gnd.n4346 gnd.n2347 9.3005
R10986 gnd.n4347 gnd.n2348 9.3005
R10987 gnd.n4350 gnd.n4349 9.3005
R10988 gnd.n4351 gnd.n2328 9.3005
R10989 gnd.n4378 gnd.n2329 9.3005
R10990 gnd.n4379 gnd.n1068 9.3005
R10991 gnd.n4380 gnd.n1069 9.3005
R10992 gnd.n4381 gnd.n1070 9.3005
R10993 gnd.n4385 gnd.n4382 9.3005
R10994 gnd.n4384 gnd.n1089 9.3005
R10995 gnd.n4383 gnd.n1090 9.3005
R10996 gnd.n2313 gnd.n1091 9.3005
R10997 gnd.n4432 gnd.n2314 9.3005
R10998 gnd.n4433 gnd.n1108 9.3005
R10999 gnd.n4434 gnd.n1109 9.3005
R11000 gnd.n4435 gnd.n1110 9.3005
R11001 gnd.n4439 gnd.n4436 9.3005
R11002 gnd.n4440 gnd.n1129 9.3005
R11003 gnd.n4675 gnd.n1130 9.3005
R11004 gnd.n4674 gnd.n1131 9.3005
R11005 gnd.n4673 gnd.n4672 9.3005
R11006 gnd.n4245 gnd.n2437 9.3005
R11007 gnd.n4126 gnd.n4125 9.3005
R11008 gnd.n4128 gnd.n4005 9.3005
R11009 gnd.n4129 gnd.n4004 9.3005
R11010 gnd.n4132 gnd.n4003 9.3005
R11011 gnd.n4133 gnd.n4002 9.3005
R11012 gnd.n4136 gnd.n4001 9.3005
R11013 gnd.n4137 gnd.n4000 9.3005
R11014 gnd.n4140 gnd.n3999 9.3005
R11015 gnd.n4141 gnd.n3998 9.3005
R11016 gnd.n4144 gnd.n3997 9.3005
R11017 gnd.n4145 gnd.n3996 9.3005
R11018 gnd.n4148 gnd.n3995 9.3005
R11019 gnd.n4149 gnd.n3994 9.3005
R11020 gnd.n4152 gnd.n3993 9.3005
R11021 gnd.n4153 gnd.n3992 9.3005
R11022 gnd.n4156 gnd.n3991 9.3005
R11023 gnd.n4157 gnd.n3990 9.3005
R11024 gnd.n4160 gnd.n3989 9.3005
R11025 gnd.n4161 gnd.n3988 9.3005
R11026 gnd.n4164 gnd.n3987 9.3005
R11027 gnd.n4168 gnd.n3983 9.3005
R11028 gnd.n4169 gnd.n3982 9.3005
R11029 gnd.n4172 gnd.n3981 9.3005
R11030 gnd.n4173 gnd.n3980 9.3005
R11031 gnd.n4176 gnd.n3979 9.3005
R11032 gnd.n4177 gnd.n3978 9.3005
R11033 gnd.n4180 gnd.n3977 9.3005
R11034 gnd.n4181 gnd.n3976 9.3005
R11035 gnd.n4184 gnd.n3975 9.3005
R11036 gnd.n4185 gnd.n3974 9.3005
R11037 gnd.n4188 gnd.n3973 9.3005
R11038 gnd.n4189 gnd.n3972 9.3005
R11039 gnd.n4192 gnd.n3971 9.3005
R11040 gnd.n4193 gnd.n3970 9.3005
R11041 gnd.n4196 gnd.n3969 9.3005
R11042 gnd.n4197 gnd.n3968 9.3005
R11043 gnd.n4200 gnd.n3967 9.3005
R11044 gnd.n4201 gnd.n3966 9.3005
R11045 gnd.n4204 gnd.n3965 9.3005
R11046 gnd.n4206 gnd.n3962 9.3005
R11047 gnd.n4209 gnd.n3961 9.3005
R11048 gnd.n4210 gnd.n3960 9.3005
R11049 gnd.n4213 gnd.n3959 9.3005
R11050 gnd.n4214 gnd.n3958 9.3005
R11051 gnd.n4217 gnd.n3957 9.3005
R11052 gnd.n4218 gnd.n3956 9.3005
R11053 gnd.n4221 gnd.n3955 9.3005
R11054 gnd.n4222 gnd.n3954 9.3005
R11055 gnd.n4225 gnd.n3953 9.3005
R11056 gnd.n4226 gnd.n3952 9.3005
R11057 gnd.n4229 gnd.n3951 9.3005
R11058 gnd.n4230 gnd.n3950 9.3005
R11059 gnd.n4233 gnd.n3949 9.3005
R11060 gnd.n4235 gnd.n3948 9.3005
R11061 gnd.n4236 gnd.n3947 9.3005
R11062 gnd.n4237 gnd.n3946 9.3005
R11063 gnd.n4238 gnd.n3945 9.3005
R11064 gnd.n4165 gnd.n3984 9.3005
R11065 gnd.n4124 gnd.n2441 9.3005
R11066 gnd.n4254 gnd.n4253 9.3005
R11067 gnd.n4255 gnd.n2426 9.3005
R11068 gnd.n4257 gnd.n4256 9.3005
R11069 gnd.n2409 gnd.n2408 9.3005
R11070 gnd.n4274 gnd.n4273 9.3005
R11071 gnd.n4275 gnd.n2407 9.3005
R11072 gnd.n4277 gnd.n4276 9.3005
R11073 gnd.n2392 gnd.n2391 9.3005
R11074 gnd.n4294 gnd.n4293 9.3005
R11075 gnd.n4295 gnd.n2390 9.3005
R11076 gnd.n4297 gnd.n4296 9.3005
R11077 gnd.n2373 gnd.n2372 9.3005
R11078 gnd.n4314 gnd.n4313 9.3005
R11079 gnd.n4315 gnd.n2371 9.3005
R11080 gnd.n4318 gnd.n4316 9.3005
R11081 gnd.n6136 gnd.n1059 9.3005
R11082 gnd.n1078 gnd.n1060 9.3005
R11083 gnd.n6126 gnd.n1079 9.3005
R11084 gnd.n6125 gnd.n1080 9.3005
R11085 gnd.n6124 gnd.n1081 9.3005
R11086 gnd.n1098 gnd.n1082 9.3005
R11087 gnd.n6114 gnd.n1099 9.3005
R11088 gnd.n6113 gnd.n1100 9.3005
R11089 gnd.n6112 gnd.n1101 9.3005
R11090 gnd.n1118 gnd.n1102 9.3005
R11091 gnd.n6102 gnd.n1119 9.3005
R11092 gnd.n6101 gnd.n1120 9.3005
R11093 gnd.n6100 gnd.n1121 9.3005
R11094 gnd.n1139 gnd.n1122 9.3005
R11095 gnd.n6090 gnd.n1140 9.3005
R11096 gnd.n6089 gnd.n6088 9.3005
R11097 gnd.n2428 gnd.n2427 9.3005
R11098 gnd.n6137 gnd.n1058 9.3005
R11099 gnd.n4401 gnd.n4400 9.3005
R11100 gnd.n6144 gnd.n1047 9.3005
R11101 gnd.n6145 gnd.n1046 9.3005
R11102 gnd.n1045 gnd.n1041 9.3005
R11103 gnd.n6151 gnd.n1040 9.3005
R11104 gnd.n6152 gnd.n1039 9.3005
R11105 gnd.n6153 gnd.n1038 9.3005
R11106 gnd.n1037 gnd.n1033 9.3005
R11107 gnd.n6159 gnd.n1032 9.3005
R11108 gnd.n6160 gnd.n1031 9.3005
R11109 gnd.n6161 gnd.n1030 9.3005
R11110 gnd.n1029 gnd.n1025 9.3005
R11111 gnd.n6167 gnd.n1024 9.3005
R11112 gnd.n6168 gnd.n1023 9.3005
R11113 gnd.n6169 gnd.n1022 9.3005
R11114 gnd.n1021 gnd.n1017 9.3005
R11115 gnd.n6175 gnd.n1016 9.3005
R11116 gnd.n6176 gnd.n1015 9.3005
R11117 gnd.n6177 gnd.n1014 9.3005
R11118 gnd.n1013 gnd.n1009 9.3005
R11119 gnd.n6183 gnd.n1008 9.3005
R11120 gnd.n6184 gnd.n1007 9.3005
R11121 gnd.n6185 gnd.n1006 9.3005
R11122 gnd.n1005 gnd.n1001 9.3005
R11123 gnd.n6191 gnd.n1000 9.3005
R11124 gnd.n6192 gnd.n999 9.3005
R11125 gnd.n6193 gnd.n998 9.3005
R11126 gnd.n997 gnd.n993 9.3005
R11127 gnd.n6199 gnd.n992 9.3005
R11128 gnd.n6200 gnd.n991 9.3005
R11129 gnd.n6201 gnd.n990 9.3005
R11130 gnd.n989 gnd.n985 9.3005
R11131 gnd.n6207 gnd.n984 9.3005
R11132 gnd.n6208 gnd.n983 9.3005
R11133 gnd.n6209 gnd.n982 9.3005
R11134 gnd.n981 gnd.n977 9.3005
R11135 gnd.n6215 gnd.n976 9.3005
R11136 gnd.n6216 gnd.n975 9.3005
R11137 gnd.n6217 gnd.n974 9.3005
R11138 gnd.n973 gnd.n969 9.3005
R11139 gnd.n6223 gnd.n968 9.3005
R11140 gnd.n6224 gnd.n967 9.3005
R11141 gnd.n6225 gnd.n966 9.3005
R11142 gnd.n965 gnd.n961 9.3005
R11143 gnd.n6231 gnd.n960 9.3005
R11144 gnd.n6232 gnd.n959 9.3005
R11145 gnd.n6233 gnd.n958 9.3005
R11146 gnd.n957 gnd.n953 9.3005
R11147 gnd.n6239 gnd.n952 9.3005
R11148 gnd.n6240 gnd.n951 9.3005
R11149 gnd.n6241 gnd.n950 9.3005
R11150 gnd.n949 gnd.n945 9.3005
R11151 gnd.n6247 gnd.n944 9.3005
R11152 gnd.n6248 gnd.n943 9.3005
R11153 gnd.n6249 gnd.n942 9.3005
R11154 gnd.n941 gnd.n937 9.3005
R11155 gnd.n6255 gnd.n936 9.3005
R11156 gnd.n6256 gnd.n935 9.3005
R11157 gnd.n6257 gnd.n934 9.3005
R11158 gnd.n933 gnd.n929 9.3005
R11159 gnd.n6263 gnd.n928 9.3005
R11160 gnd.n6264 gnd.n927 9.3005
R11161 gnd.n6265 gnd.n926 9.3005
R11162 gnd.n925 gnd.n921 9.3005
R11163 gnd.n6271 gnd.n920 9.3005
R11164 gnd.n6272 gnd.n919 9.3005
R11165 gnd.n6273 gnd.n918 9.3005
R11166 gnd.n917 gnd.n913 9.3005
R11167 gnd.n6279 gnd.n912 9.3005
R11168 gnd.n6280 gnd.n911 9.3005
R11169 gnd.n6281 gnd.n910 9.3005
R11170 gnd.n909 gnd.n905 9.3005
R11171 gnd.n6287 gnd.n904 9.3005
R11172 gnd.n6288 gnd.n903 9.3005
R11173 gnd.n6289 gnd.n902 9.3005
R11174 gnd.n901 gnd.n897 9.3005
R11175 gnd.n6295 gnd.n896 9.3005
R11176 gnd.n6296 gnd.n895 9.3005
R11177 gnd.n6297 gnd.n894 9.3005
R11178 gnd.n893 gnd.n889 9.3005
R11179 gnd.n6303 gnd.n888 9.3005
R11180 gnd.n6304 gnd.n887 9.3005
R11181 gnd.n6305 gnd.n886 9.3005
R11182 gnd.n882 gnd.n881 9.3005
R11183 gnd.n6312 gnd.n6311 9.3005
R11184 gnd.n6143 gnd.n1048 9.3005
R11185 gnd.n5531 gnd.n1485 9.3005
R11186 gnd.n4732 gnd.n4721 9.3005
R11187 gnd.n4731 gnd.n4730 9.3005
R11188 gnd.n4729 gnd.n4724 9.3005
R11189 gnd.n4728 gnd.n4727 9.3005
R11190 gnd.n2256 gnd.n2255 9.3005
R11191 gnd.n4780 gnd.n4779 9.3005
R11192 gnd.n4781 gnd.n2253 9.3005
R11193 gnd.n4786 gnd.n4785 9.3005
R11194 gnd.n4784 gnd.n2254 9.3005
R11195 gnd.n4783 gnd.n4782 9.3005
R11196 gnd.n1399 gnd.n1397 9.3005
R11197 gnd.n5931 gnd.n5930 9.3005
R11198 gnd.n5929 gnd.n1398 9.3005
R11199 gnd.n5928 gnd.n5927 9.3005
R11200 gnd.n5926 gnd.n1400 9.3005
R11201 gnd.n5925 gnd.n5924 9.3005
R11202 gnd.n5923 gnd.n1404 9.3005
R11203 gnd.n5922 gnd.n5921 9.3005
R11204 gnd.n5920 gnd.n1405 9.3005
R11205 gnd.n5919 gnd.n5918 9.3005
R11206 gnd.n5917 gnd.n1409 9.3005
R11207 gnd.n5916 gnd.n5915 9.3005
R11208 gnd.n5914 gnd.n1410 9.3005
R11209 gnd.n5913 gnd.n5912 9.3005
R11210 gnd.n5911 gnd.n1414 9.3005
R11211 gnd.n5910 gnd.n5909 9.3005
R11212 gnd.n5908 gnd.n1415 9.3005
R11213 gnd.n5907 gnd.n5906 9.3005
R11214 gnd.n5905 gnd.n1419 9.3005
R11215 gnd.n5904 gnd.n5903 9.3005
R11216 gnd.n5902 gnd.n1420 9.3005
R11217 gnd.n5901 gnd.n5900 9.3005
R11218 gnd.n5899 gnd.n1424 9.3005
R11219 gnd.n5898 gnd.n5897 9.3005
R11220 gnd.n5896 gnd.n1425 9.3005
R11221 gnd.n5895 gnd.n5894 9.3005
R11222 gnd.n5893 gnd.n1429 9.3005
R11223 gnd.n5892 gnd.n5891 9.3005
R11224 gnd.n5890 gnd.n1430 9.3005
R11225 gnd.n5889 gnd.n5888 9.3005
R11226 gnd.n5887 gnd.n1434 9.3005
R11227 gnd.n5886 gnd.n5885 9.3005
R11228 gnd.n5884 gnd.n1435 9.3005
R11229 gnd.n5883 gnd.n5882 9.3005
R11230 gnd.n5881 gnd.n1439 9.3005
R11231 gnd.n5880 gnd.n5879 9.3005
R11232 gnd.n5878 gnd.n1440 9.3005
R11233 gnd.n5877 gnd.n5876 9.3005
R11234 gnd.n5875 gnd.n1444 9.3005
R11235 gnd.n5874 gnd.n5873 9.3005
R11236 gnd.n5872 gnd.n1445 9.3005
R11237 gnd.n5871 gnd.n5870 9.3005
R11238 gnd.n5869 gnd.n1449 9.3005
R11239 gnd.n5868 gnd.n5867 9.3005
R11240 gnd.n5866 gnd.n1450 9.3005
R11241 gnd.n5865 gnd.n5864 9.3005
R11242 gnd.n5863 gnd.n1454 9.3005
R11243 gnd.n5862 gnd.n5861 9.3005
R11244 gnd.n5860 gnd.n1455 9.3005
R11245 gnd.n5859 gnd.n5858 9.3005
R11246 gnd.n5857 gnd.n1459 9.3005
R11247 gnd.n5856 gnd.n5855 9.3005
R11248 gnd.n5854 gnd.n1460 9.3005
R11249 gnd.n5853 gnd.n5852 9.3005
R11250 gnd.n5851 gnd.n1464 9.3005
R11251 gnd.n5850 gnd.n5849 9.3005
R11252 gnd.n5848 gnd.n1465 9.3005
R11253 gnd.n5847 gnd.n5846 9.3005
R11254 gnd.n5845 gnd.n1469 9.3005
R11255 gnd.n5844 gnd.n5843 9.3005
R11256 gnd.n5842 gnd.n1470 9.3005
R11257 gnd.n5841 gnd.n5840 9.3005
R11258 gnd.n5839 gnd.n1474 9.3005
R11259 gnd.n5838 gnd.n5837 9.3005
R11260 gnd.n5836 gnd.n1475 9.3005
R11261 gnd.n5835 gnd.n5834 9.3005
R11262 gnd.n5833 gnd.n1479 9.3005
R11263 gnd.n5832 gnd.n5831 9.3005
R11264 gnd.n5830 gnd.n1480 9.3005
R11265 gnd.n5829 gnd.n5828 9.3005
R11266 gnd.n5827 gnd.n1484 9.3005
R11267 gnd.n5826 gnd.n5825 9.3005
R11268 gnd.n4734 gnd.n4733 9.3005
R11269 gnd.n4736 gnd.n4735 9.3005
R11270 gnd.n4048 gnd.n4047 9.3005
R11271 gnd.n2332 gnd.n2331 9.3005
R11272 gnd.n4371 gnd.n4370 9.3005
R11273 gnd.n4372 gnd.n2330 9.3005
R11274 gnd.n4374 gnd.n4373 9.3005
R11275 gnd.n2327 gnd.n2325 9.3005
R11276 gnd.n4393 gnd.n4392 9.3005
R11277 gnd.n4391 gnd.n2326 9.3005
R11278 gnd.n4390 gnd.n4389 9.3005
R11279 gnd.n2317 gnd.n2316 9.3005
R11280 gnd.n4425 gnd.n4424 9.3005
R11281 gnd.n4426 gnd.n2315 9.3005
R11282 gnd.n4428 gnd.n4427 9.3005
R11283 gnd.n2310 gnd.n2308 9.3005
R11284 gnd.n4688 gnd.n4687 9.3005
R11285 gnd.n4686 gnd.n2309 9.3005
R11286 gnd.n4685 gnd.n4684 9.3005
R11287 gnd.n4683 gnd.n2311 9.3005
R11288 gnd.n4682 gnd.n4681 9.3005
R11289 gnd.n4680 gnd.n4679 9.3005
R11290 gnd.n2295 gnd.n2290 9.3005
R11291 gnd.n4566 gnd.n4565 9.3005
R11292 gnd.n4465 gnd.n4464 9.3005
R11293 gnd.n4560 gnd.n4559 9.3005
R11294 gnd.n4558 gnd.n4557 9.3005
R11295 gnd.n4477 gnd.n4476 9.3005
R11296 gnd.n4552 gnd.n4551 9.3005
R11297 gnd.n4550 gnd.n4549 9.3005
R11298 gnd.n4485 gnd.n4484 9.3005
R11299 gnd.n4544 gnd.n4543 9.3005
R11300 gnd.n4542 gnd.n4541 9.3005
R11301 gnd.n4497 gnd.n4496 9.3005
R11302 gnd.n4536 gnd.n4535 9.3005
R11303 gnd.n4534 gnd.n4533 9.3005
R11304 gnd.n4505 gnd.n4504 9.3005
R11305 gnd.n4528 gnd.n4527 9.3005
R11306 gnd.n4526 gnd.n4525 9.3005
R11307 gnd.n4516 gnd.n2294 9.3005
R11308 gnd.n4718 gnd.n4717 9.3005
R11309 gnd.n4568 gnd.n4567 9.3005
R11310 gnd.n4719 gnd.n2289 9.3005
R11311 gnd.n4522 gnd.n2291 9.3005
R11312 gnd.n4524 gnd.n4523 9.3005
R11313 gnd.n4511 gnd.n4510 9.3005
R11314 gnd.n4530 gnd.n4529 9.3005
R11315 gnd.n4532 gnd.n4531 9.3005
R11316 gnd.n4501 gnd.n4500 9.3005
R11317 gnd.n4538 gnd.n4537 9.3005
R11318 gnd.n4540 gnd.n4539 9.3005
R11319 gnd.n4491 gnd.n4490 9.3005
R11320 gnd.n4546 gnd.n4545 9.3005
R11321 gnd.n4548 gnd.n4547 9.3005
R11322 gnd.n4481 gnd.n4480 9.3005
R11323 gnd.n4554 gnd.n4553 9.3005
R11324 gnd.n4556 gnd.n4555 9.3005
R11325 gnd.n4471 gnd.n4470 9.3005
R11326 gnd.n4562 gnd.n4561 9.3005
R11327 gnd.n4564 gnd.n4563 9.3005
R11328 gnd.n4462 gnd.n4461 9.3005
R11329 gnd.n4570 gnd.n4569 9.3005
R11330 gnd.n4571 gnd.n4441 9.3005
R11331 gnd.n4573 gnd.n4572 9.3005
R11332 gnd.n4456 gnd.n4442 9.3005
R11333 gnd.n4455 gnd.n4454 9.3005
R11334 gnd.n4453 gnd.n4443 9.3005
R11335 gnd.n4452 gnd.n4451 9.3005
R11336 gnd.n4448 gnd.n4446 9.3005
R11337 gnd.n4447 gnd.n2262 9.3005
R11338 gnd.n4759 gnd.n2261 9.3005
R11339 gnd.n4761 gnd.n4760 9.3005
R11340 gnd.n2259 gnd.n2258 9.3005
R11341 gnd.n4766 gnd.n4765 9.3005
R11342 gnd.n4767 gnd.n2257 9.3005
R11343 gnd.n4769 gnd.n4768 9.3005
R11344 gnd.n2250 gnd.n2249 9.3005
R11345 gnd.n4791 gnd.n4790 9.3005
R11346 gnd.n4792 gnd.n2248 9.3005
R11347 gnd.n4794 gnd.n4793 9.3005
R11348 gnd.n4825 gnd.n2247 9.3005
R11349 gnd.n4827 gnd.n4826 9.3005
R11350 gnd.n4828 gnd.n2245 9.3005
R11351 gnd.n4835 gnd.n4834 9.3005
R11352 gnd.n4833 gnd.n2246 9.3005
R11353 gnd.n4832 gnd.n4831 9.3005
R11354 gnd.n4830 gnd.n4829 9.3005
R11355 gnd.n2219 gnd.n2218 9.3005
R11356 gnd.n4890 gnd.n4889 9.3005
R11357 gnd.n4891 gnd.n2217 9.3005
R11358 gnd.n4893 gnd.n4892 9.3005
R11359 gnd.n4894 gnd.n2216 9.3005
R11360 gnd.n4898 gnd.n4897 9.3005
R11361 gnd.n4899 gnd.n2214 9.3005
R11362 gnd.n4928 gnd.n4927 9.3005
R11363 gnd.n4926 gnd.n2215 9.3005
R11364 gnd.n4925 gnd.n4924 9.3005
R11365 gnd.n4923 gnd.n4900 9.3005
R11366 gnd.n4922 gnd.n4921 9.3005
R11367 gnd.n4920 gnd.n4903 9.3005
R11368 gnd.n4919 gnd.n4918 9.3005
R11369 gnd.n4917 gnd.n4904 9.3005
R11370 gnd.n4916 gnd.n4915 9.3005
R11371 gnd.n4914 gnd.n4911 9.3005
R11372 gnd.n4913 gnd.n4912 9.3005
R11373 gnd.n2119 gnd.n2118 9.3005
R11374 gnd.n5063 gnd.n5062 9.3005
R11375 gnd.n5064 gnd.n2116 9.3005
R11376 gnd.n5087 gnd.n5086 9.3005
R11377 gnd.n5085 gnd.n2117 9.3005
R11378 gnd.n5084 gnd.n5083 9.3005
R11379 gnd.n5082 gnd.n5065 9.3005
R11380 gnd.n5081 gnd.n5080 9.3005
R11381 gnd.n5079 gnd.n5068 9.3005
R11382 gnd.n5078 gnd.n5077 9.3005
R11383 gnd.n5076 gnd.n5069 9.3005
R11384 gnd.n5075 gnd.n5074 9.3005
R11385 gnd.n5073 gnd.n5072 9.3005
R11386 gnd.n2055 gnd.n2054 9.3005
R11387 gnd.n5188 gnd.n5187 9.3005
R11388 gnd.n5189 gnd.n2052 9.3005
R11389 gnd.n5195 gnd.n5194 9.3005
R11390 gnd.n5193 gnd.n2053 9.3005
R11391 gnd.n5192 gnd.n5191 9.3005
R11392 gnd.n5190 gnd.n2030 9.3005
R11393 gnd.n2028 gnd.n2027 9.3005
R11394 gnd.n5226 gnd.n5225 9.3005
R11395 gnd.n5227 gnd.n2025 9.3005
R11396 gnd.n5258 gnd.n5257 9.3005
R11397 gnd.n5256 gnd.n2026 9.3005
R11398 gnd.n5255 gnd.n5254 9.3005
R11399 gnd.n5253 gnd.n5228 9.3005
R11400 gnd.n5252 gnd.n5251 9.3005
R11401 gnd.n5250 gnd.n5230 9.3005
R11402 gnd.n5249 gnd.n5248 9.3005
R11403 gnd.n5247 gnd.n5231 9.3005
R11404 gnd.n5246 gnd.n5245 9.3005
R11405 gnd.n5244 gnd.n5236 9.3005
R11406 gnd.n5243 gnd.n5242 9.3005
R11407 gnd.n5241 gnd.n5237 9.3005
R11408 gnd.n5240 gnd.n5239 9.3005
R11409 gnd.n1929 gnd.n1928 9.3005
R11410 gnd.n5390 gnd.n5389 9.3005
R11411 gnd.n5391 gnd.n1926 9.3005
R11412 gnd.n5394 gnd.n5393 9.3005
R11413 gnd.n5392 gnd.n1927 9.3005
R11414 gnd.n1782 gnd.n1781 9.3005
R11415 gnd.n5499 gnd.n5498 9.3005
R11416 gnd.n5500 gnd.n1780 9.3005
R11417 gnd.n5502 gnd.n5501 9.3005
R11418 gnd.n1494 gnd.n1493 9.3005
R11419 gnd.n5821 gnd.n5820 9.3005
R11420 gnd.n4758 gnd.n4757 9.3005
R11421 gnd.n5817 gnd.n1495 9.3005
R11422 gnd.n5816 gnd.n5815 9.3005
R11423 gnd.n5814 gnd.n1498 9.3005
R11424 gnd.n5813 gnd.n5812 9.3005
R11425 gnd.n5811 gnd.n1499 9.3005
R11426 gnd.n5810 gnd.n5809 9.3005
R11427 gnd.n5819 gnd.n5818 9.3005
R11428 gnd.n5762 gnd.n5761 9.3005
R11429 gnd.n1546 gnd.n1545 9.3005
R11430 gnd.n5768 gnd.n5767 9.3005
R11431 gnd.n5770 gnd.n5769 9.3005
R11432 gnd.n1538 gnd.n1537 9.3005
R11433 gnd.n5776 gnd.n5775 9.3005
R11434 gnd.n5778 gnd.n5777 9.3005
R11435 gnd.n1530 gnd.n1529 9.3005
R11436 gnd.n5784 gnd.n5783 9.3005
R11437 gnd.n5786 gnd.n5785 9.3005
R11438 gnd.n1522 gnd.n1521 9.3005
R11439 gnd.n5792 gnd.n5791 9.3005
R11440 gnd.n5794 gnd.n5793 9.3005
R11441 gnd.n1514 gnd.n1513 9.3005
R11442 gnd.n5800 gnd.n5799 9.3005
R11443 gnd.n5802 gnd.n5801 9.3005
R11444 gnd.n1510 gnd.n1505 9.3005
R11445 gnd.n5760 gnd.n1555 9.3005
R11446 gnd.n1746 gnd.n1554 9.3005
R11447 gnd.n5807 gnd.n1503 9.3005
R11448 gnd.n5806 gnd.n5805 9.3005
R11449 gnd.n5804 gnd.n5803 9.3005
R11450 gnd.n1509 gnd.n1508 9.3005
R11451 gnd.n5798 gnd.n5797 9.3005
R11452 gnd.n5796 gnd.n5795 9.3005
R11453 gnd.n1518 gnd.n1517 9.3005
R11454 gnd.n5790 gnd.n5789 9.3005
R11455 gnd.n5788 gnd.n5787 9.3005
R11456 gnd.n1526 gnd.n1525 9.3005
R11457 gnd.n5782 gnd.n5781 9.3005
R11458 gnd.n5780 gnd.n5779 9.3005
R11459 gnd.n1534 gnd.n1533 9.3005
R11460 gnd.n5774 gnd.n5773 9.3005
R11461 gnd.n5772 gnd.n5771 9.3005
R11462 gnd.n1542 gnd.n1541 9.3005
R11463 gnd.n5766 gnd.n5765 9.3005
R11464 gnd.n5764 gnd.n5763 9.3005
R11465 gnd.n1769 gnd.n1552 9.3005
R11466 gnd.n1748 gnd.n1747 9.3005
R11467 gnd.n5533 gnd.n5532 9.3005
R11468 gnd.n5570 gnd.n5569 9.3005
R11469 gnd.n5568 gnd.n1745 9.3005
R11470 gnd.n5567 gnd.n5566 9.3005
R11471 gnd.n5565 gnd.n5536 9.3005
R11472 gnd.n5564 gnd.n5563 9.3005
R11473 gnd.n5562 gnd.n5540 9.3005
R11474 gnd.n5561 gnd.n5560 9.3005
R11475 gnd.n5559 gnd.n5541 9.3005
R11476 gnd.n5558 gnd.n5557 9.3005
R11477 gnd.n5556 gnd.n5553 9.3005
R11478 gnd.n5555 gnd.n5554 9.3005
R11479 gnd.n534 gnd.n533 9.3005
R11480 gnd.n6878 gnd.n6877 9.3005
R11481 gnd.n6879 gnd.n532 9.3005
R11482 gnd.n6881 gnd.n6880 9.3005
R11483 gnd.n515 gnd.n514 9.3005
R11484 gnd.n6905 gnd.n6904 9.3005
R11485 gnd.n6906 gnd.n512 9.3005
R11486 gnd.n6908 gnd.n6907 9.3005
R11487 gnd.n513 gnd.n63 9.3005
R11488 gnd.n5535 gnd.n1744 9.3005
R11489 gnd.n7030 gnd.n64 9.3005
R11490 gnd.t323 gnd.n2633 9.24152
R11491 gnd.n2535 gnd.t171 9.24152
R11492 gnd.n3804 gnd.t158 9.24152
R11493 gnd.t36 gnd.t323 8.92286
R11494 gnd.n5960 gnd.n1276 8.92286
R11495 gnd.n4940 gnd.n2191 8.92286
R11496 gnd.n4966 gnd.n2167 8.92286
R11497 gnd.n5017 gnd.n5016 8.92286
R11498 gnd.n5127 gnd.n2084 8.92286
R11499 gnd.n5221 gnd.n2033 8.92286
R11500 gnd.n5297 gnd.n5296 8.92286
R11501 gnd.n5360 gnd.n1942 8.92286
R11502 gnd.n5496 gnd.n1784 8.92286
R11503 gnd.n3774 gnd.n3749 8.92171
R11504 gnd.n3742 gnd.n3717 8.92171
R11505 gnd.n3710 gnd.n3685 8.92171
R11506 gnd.n3679 gnd.n3654 8.92171
R11507 gnd.n3647 gnd.n3622 8.92171
R11508 gnd.n3615 gnd.n3590 8.92171
R11509 gnd.n3583 gnd.n3558 8.92171
R11510 gnd.n3552 gnd.n3527 8.92171
R11511 gnd.n1835 gnd.n1817 8.72777
R11512 gnd.n3277 gnd.t50 8.60421
R11513 gnd.n6030 gnd.n1218 8.60421
R11514 gnd.n5090 gnd.t308 8.60421
R11515 gnd.n5112 gnd.t34 8.60421
R11516 gnd.n2697 gnd.n2685 8.43656
R11517 gnd.n38 gnd.n26 8.43656
R11518 gnd.t137 gnd.n1250 8.28555
R11519 gnd.n3775 gnd.n3747 8.14595
R11520 gnd.n3743 gnd.n3715 8.14595
R11521 gnd.n3711 gnd.n3683 8.14595
R11522 gnd.n3680 gnd.n3652 8.14595
R11523 gnd.n3648 gnd.n3620 8.14595
R11524 gnd.n3616 gnd.n3588 8.14595
R11525 gnd.n3584 gnd.n3556 8.14595
R11526 gnd.n3553 gnd.n3525 8.14595
R11527 gnd.n4049 gnd.n0 8.10675
R11528 gnd.n7031 gnd.n7030 8.10675
R11529 gnd.n3780 gnd.n3779 7.97301
R11530 gnd.t184 gnd.n2792 7.9669
R11531 gnd.n4866 gnd.t2 7.9669
R11532 gnd.n5333 gnd.t4 7.9669
R11533 gnd.n7031 gnd.n62 7.78567
R11534 gnd.n5760 gnd.n1554 7.75808
R11535 gnd.n4717 gnd.n2294 7.75808
R11536 gnd.n250 gnd.n199 7.75808
R11537 gnd.n4084 gnd.n4026 7.75808
R11538 gnd.n3518 gnd.n2532 7.64824
R11539 gnd.n4788 gnd.t178 7.64824
R11540 gnd.n5933 gnd.n1392 7.64824
R11541 gnd.t6 gnd.n2223 7.64824
R11542 gnd.t33 gnd.n4908 7.64824
R11543 gnd.n4909 gnd.t33 7.64824
R11544 gnd.n5175 gnd.t12 7.64824
R11545 gnd.t12 gnd.n5174 7.64824
R11546 gnd.n1995 gnd.t45 7.64824
R11547 gnd.n5355 gnd.n1953 7.64824
R11548 gnd.n5387 gnd.t149 7.64824
R11549 gnd.n2722 gnd.n2721 7.53171
R11550 gnd.n3186 gnd.t315 7.32958
R11551 gnd.t319 gnd.t96 7.32958
R11552 gnd.n1272 gnd.n1271 7.30353
R11553 gnd.n1834 gnd.n1833 7.30353
R11554 gnd.n3146 gnd.n2865 7.01093
R11555 gnd.n2868 gnd.n2866 7.01093
R11556 gnd.n3156 gnd.n3155 7.01093
R11557 gnd.n3167 gnd.n2849 7.01093
R11558 gnd.n3166 gnd.n2852 7.01093
R11559 gnd.n3177 gnd.n2840 7.01093
R11560 gnd.n2843 gnd.n2841 7.01093
R11561 gnd.n3187 gnd.n3186 7.01093
R11562 gnd.n3197 gnd.n2821 7.01093
R11563 gnd.n3196 gnd.n2824 7.01093
R11564 gnd.n3205 gnd.n2815 7.01093
R11565 gnd.n3217 gnd.n2805 7.01093
R11566 gnd.n3227 gnd.n2790 7.01093
R11567 gnd.n3243 gnd.n3242 7.01093
R11568 gnd.n2792 gnd.n2729 7.01093
R11569 gnd.n3297 gnd.n2730 7.01093
R11570 gnd.n3291 gnd.n3290 7.01093
R11571 gnd.n2779 gnd.n2741 7.01093
R11572 gnd.n3283 gnd.n2752 7.01093
R11573 gnd.n2770 gnd.n2765 7.01093
R11574 gnd.n3277 gnd.n3276 7.01093
R11575 gnd.n3323 gnd.n2668 7.01093
R11576 gnd.n3322 gnd.n3321 7.01093
R11577 gnd.n3334 gnd.n3333 7.01093
R11578 gnd.n2661 gnd.n2653 7.01093
R11579 gnd.n3363 gnd.n2641 7.01093
R11580 gnd.n3362 gnd.n2644 7.01093
R11581 gnd.n3373 gnd.n2633 7.01093
R11582 gnd.n2634 gnd.n2622 7.01093
R11583 gnd.n3384 gnd.n2623 7.01093
R11584 gnd.n3408 gnd.n2614 7.01093
R11585 gnd.n3407 gnd.n2605 7.01093
R11586 gnd.n3430 gnd.n3429 7.01093
R11587 gnd.n3448 gnd.n2586 7.01093
R11588 gnd.n3447 gnd.n2589 7.01093
R11589 gnd.n3458 gnd.n2578 7.01093
R11590 gnd.n2579 gnd.n2566 7.01093
R11591 gnd.n3469 gnd.n2567 7.01093
R11592 gnd.n3496 gnd.n2551 7.01093
R11593 gnd.n3508 gnd.n3507 7.01093
R11594 gnd.n3490 gnd.n2544 7.01093
R11595 gnd.n3520 gnd.n3519 7.01093
R11596 gnd.n3792 gnd.n2532 7.01093
R11597 gnd.n3791 gnd.n2535 7.01093
R11598 gnd.n3804 gnd.n2524 7.01093
R11599 gnd.n2525 gnd.n2517 7.01093
R11600 gnd.n3814 gnd.n2443 7.01093
R11601 gnd.t31 gnd.n2133 7.01093
R11602 gnd.n5135 gnd.t16 7.01093
R11603 gnd.n5496 gnd.t110 7.01093
R11604 gnd.n2824 gnd.t8 6.69227
R11605 gnd.n2644 gnd.t36 6.69227
R11606 gnd.n3497 gnd.t18 6.69227
R11607 gnd.n4691 gnd.t200 6.69227
R11608 gnd.n4851 gnd.t13 6.69227
R11609 gnd.n5304 gnd.t321 6.69227
R11610 gnd.t207 gnd.n1707 6.69227
R11611 gnd.n5468 gnd.n5467 6.5566
R11612 gnd.n1302 gnd.n1301 6.5566
R11613 gnd.n5971 gnd.n5967 6.5566
R11614 gnd.n1895 gnd.n1894 6.5566
R11615 gnd.n4837 gnd.n2243 6.37362
R11616 gnd.n4879 gnd.n4877 6.37362
R11617 gnd.n4905 gnd.n2158 6.37362
R11618 gnd.n2060 gnd.n2049 6.37362
R11619 gnd.n5321 gnd.n1981 6.37362
R11620 gnd.n5234 gnd.n1957 6.37362
R11621 gnd.n5484 gnd.t65 6.37362
R11622 gnd.n4523 gnd.n4519 6.20656
R11623 gnd.n1769 gnd.n1551 6.20656
R11624 gnd.t40 gnd.n3253 6.05496
R11625 gnd.n3254 gnd.t60 6.05496
R11626 gnd.t46 gnd.n2668 6.05496
R11627 gnd.t9 gnd.n3418 6.05496
R11628 gnd.n4396 gnd.t194 6.05496
R11629 gnd.n6856 gnd.t220 6.05496
R11630 gnd.n3777 gnd.n3747 5.81868
R11631 gnd.n3745 gnd.n3715 5.81868
R11632 gnd.n3713 gnd.n3683 5.81868
R11633 gnd.n3682 gnd.n3652 5.81868
R11634 gnd.n3650 gnd.n3620 5.81868
R11635 gnd.n3618 gnd.n3588 5.81868
R11636 gnd.n3586 gnd.n3556 5.81868
R11637 gnd.n3555 gnd.n3525 5.81868
R11638 gnd.n5940 gnd.t71 5.73631
R11639 gnd.n2191 gnd.t52 5.73631
R11640 gnd.n5005 gnd.t28 5.73631
R11641 gnd.t10 gnd.n2058 5.73631
R11642 gnd.n5297 gnd.t11 5.73631
R11643 gnd.n5477 gnd.t110 5.73631
R11644 gnd.n5472 gnd.n1631 5.62001
R11645 gnd.n6033 gnd.n1214 5.62001
R11646 gnd.n6033 gnd.n1215 5.62001
R11647 gnd.n1899 gnd.n1631 5.62001
R11648 gnd.n3005 gnd.n3000 5.4308
R11649 gnd.n3822 gnd.n2510 5.4308
R11650 gnd.n3321 gnd.t61 5.41765
R11651 gnd.t51 gnd.n3344 5.41765
R11652 gnd.t25 gnd.n2598 5.41765
R11653 gnd.n4932 gnd.t324 5.41765
R11654 gnd.n2019 gnd.t55 5.41765
R11655 gnd.n4376 gnd.n1053 5.09899
R11656 gnd.n6134 gnd.n1062 5.09899
R11657 gnd.n4396 gnd.n4395 5.09899
R11658 gnd.n6128 gnd.n1073 5.09899
R11659 gnd.n4387 gnd.n1076 5.09899
R11660 gnd.n6122 gnd.n1084 5.09899
R11661 gnd.n4422 gnd.n1087 5.09899
R11662 gnd.n4430 gnd.n1096 5.09899
R11663 gnd.n6110 gnd.n1104 5.09899
R11664 gnd.n4691 gnd.n4690 5.09899
R11665 gnd.n6104 gnd.n1113 5.09899
R11666 gnd.n4437 gnd.n1116 5.09899
R11667 gnd.n6098 gnd.n1124 5.09899
R11668 gnd.n4677 gnd.n1127 5.09899
R11669 gnd.n6092 gnd.n1134 5.09899
R11670 gnd.n4714 gnd.n1137 5.09899
R11671 gnd.n4846 gnd.n4845 5.09899
R11672 gnd.n4866 gnd.n4865 5.09899
R11673 gnd.t1 gnd.n4986 5.09899
R11674 gnd.n5004 gnd.n2142 5.09899
R11675 gnd.n5011 gnd.n2144 5.09899
R11676 gnd.n5156 gnd.n2069 5.09899
R11677 gnd.n5185 gnd.n2057 5.09899
R11678 gnd.n5211 gnd.t30 5.09899
R11679 gnd.n5333 gnd.n1973 5.09899
R11680 gnd.n5340 gnd.n1967 5.09899
R11681 gnd.n5634 gnd.n1669 5.09899
R11682 gnd.n5573 gnd.n5572 5.09899
R11683 gnd.n5626 gnd.n1678 5.09899
R11684 gnd.n5537 gnd.n1691 5.09899
R11685 gnd.n5620 gnd.n1694 5.09899
R11686 gnd.n5543 gnd.n1704 5.09899
R11687 gnd.n5614 gnd.n1707 5.09899
R11688 gnd.n5550 gnd.n1716 5.09899
R11689 gnd.n5608 gnd.n1719 5.09899
R11690 gnd.n1732 gnd.n546 5.09899
R11691 gnd.n6864 gnd.n549 5.09899
R11692 gnd.n1725 gnd.n536 5.09899
R11693 gnd.n6875 gnd.n538 5.09899
R11694 gnd.n6857 gnd.n6856 5.09899
R11695 gnd.n6883 gnd.n522 5.09899
R11696 gnd.n6897 gnd.n517 5.09899
R11697 gnd.n3775 gnd.n3774 5.04292
R11698 gnd.n3743 gnd.n3742 5.04292
R11699 gnd.n3711 gnd.n3710 5.04292
R11700 gnd.n3680 gnd.n3679 5.04292
R11701 gnd.n3648 gnd.n3647 5.04292
R11702 gnd.n3616 gnd.n3615 5.04292
R11703 gnd.n3584 gnd.n3583 5.04292
R11704 gnd.n3553 gnd.n3552 5.04292
R11705 gnd.n3284 gnd.t58 4.78034
R11706 gnd.n2623 gnd.t57 4.78034
R11707 gnd.n4959 gnd.t324 4.78034
R11708 gnd.t55 gnd.n2010 4.78034
R11709 gnd.n5475 gnd.t86 4.78034
R11710 gnd.n2726 gnd.n2723 4.74817
R11711 gnd.n2776 gnd.n2674 4.74817
R11712 gnd.n2763 gnd.n2673 4.74817
R11713 gnd.n2672 gnd.n2671 4.74817
R11714 gnd.n2772 gnd.n2723 4.74817
R11715 gnd.n2773 gnd.n2674 4.74817
R11716 gnd.n2775 gnd.n2673 4.74817
R11717 gnd.n2762 gnd.n2672 4.74817
R11718 gnd.n6900 gnd.n81 4.74817
R11719 gnd.n6915 gnd.n80 4.74817
R11720 gnd.n6913 gnd.n79 4.74817
R11721 gnd.n7023 gnd.n74 4.74817
R11722 gnd.n7021 gnd.n75 4.74817
R11723 gnd.n521 gnd.n81 4.74817
R11724 gnd.n6899 gnd.n80 4.74817
R11725 gnd.n6916 gnd.n79 4.74817
R11726 gnd.n6912 gnd.n74 4.74817
R11727 gnd.n7022 gnd.n7021 4.74817
R11728 gnd.n4334 gnd.n2356 4.74817
R11729 gnd.n4338 gnd.n4336 4.74817
R11730 gnd.n4361 gnd.n2337 4.74817
R11731 gnd.n4365 gnd.n4363 4.74817
R11732 gnd.n6138 gnd.n1057 4.74817
R11733 gnd.n4317 gnd.n2356 4.74817
R11734 gnd.n4336 gnd.n4335 4.74817
R11735 gnd.n4337 gnd.n2337 4.74817
R11736 gnd.n4363 gnd.n4362 4.74817
R11737 gnd.n4364 gnd.n1057 4.74817
R11738 gnd.n2721 gnd.n2720 4.74296
R11739 gnd.n62 gnd.n61 4.74296
R11740 gnd.n2697 gnd.n2696 4.7074
R11741 gnd.n2709 gnd.n2708 4.7074
R11742 gnd.n38 gnd.n37 4.7074
R11743 gnd.n50 gnd.n49 4.7074
R11744 gnd.n2721 gnd.n2709 4.65959
R11745 gnd.n62 gnd.n50 4.65959
R11746 gnd.n5702 gnd.n1633 4.6132
R11747 gnd.n6034 gnd.n1213 4.6132
R11748 gnd.n6084 gnd.n1144 4.46168
R11749 gnd.t305 gnd.n1392 4.46168
R11750 gnd.n5355 gnd.t7 4.46168
R11751 gnd.n5755 gnd.n1599 4.46168
R11752 gnd.n1830 gnd.n1817 4.46111
R11753 gnd.n3760 gnd.n3756 4.38594
R11754 gnd.n3728 gnd.n3724 4.38594
R11755 gnd.n3696 gnd.n3692 4.38594
R11756 gnd.n3665 gnd.n3661 4.38594
R11757 gnd.n3633 gnd.n3629 4.38594
R11758 gnd.n3601 gnd.n3597 4.38594
R11759 gnd.n3569 gnd.n3565 4.38594
R11760 gnd.n3538 gnd.n3534 4.38594
R11761 gnd.n3771 gnd.n3749 4.26717
R11762 gnd.n3739 gnd.n3717 4.26717
R11763 gnd.n3707 gnd.n3685 4.26717
R11764 gnd.n3676 gnd.n3654 4.26717
R11765 gnd.n3644 gnd.n3622 4.26717
R11766 gnd.n3612 gnd.n3590 4.26717
R11767 gnd.n3580 gnd.n3558 4.26717
R11768 gnd.n3549 gnd.n3527 4.26717
R11769 gnd.n3228 gnd.t19 4.14303
R11770 gnd.n3458 gnd.t59 4.14303
R11771 gnd.n4421 gnd.t210 4.14303
R11772 gnd.n5038 gnd.t38 4.14303
R11773 gnd.n5162 gnd.t326 4.14303
R11774 gnd.t185 gnd.n5600 4.14303
R11775 gnd.n3779 gnd.n3778 4.08274
R11776 gnd.n5467 gnd.n5466 4.05904
R11777 gnd.n1303 gnd.n1302 4.05904
R11778 gnd.n5974 gnd.n5967 4.05904
R11779 gnd.n1894 gnd.n1893 4.05904
R11780 gnd.n15 gnd.n7 3.99943
R11781 gnd.n5946 gnd.t178 3.82437
R11782 gnd.n4815 gnd.n4802 3.82437
R11783 gnd.n2232 gnd.n2231 3.82437
R11784 gnd.n4994 gnd.n4993 3.82437
R11785 gnd.n5050 gnd.n2130 3.82437
R11786 gnd.n5163 gnd.n2074 3.82437
R11787 gnd.n5198 gnd.n5197 3.82437
R11788 gnd.n5314 gnd.n1978 3.82437
R11789 gnd.n5349 gnd.n5348 3.82437
R11790 gnd.n5504 gnd.t86 3.82437
R11791 gnd.n3301 gnd.n2722 3.81325
R11792 gnd.n2709 gnd.n2697 3.72967
R11793 gnd.n50 gnd.n38 3.72967
R11794 gnd.n3779 gnd.n3651 3.70378
R11795 gnd.n15 gnd.n14 3.60163
R11796 gnd.n3770 gnd.n3751 3.49141
R11797 gnd.n3738 gnd.n3719 3.49141
R11798 gnd.n3706 gnd.n3687 3.49141
R11799 gnd.n3675 gnd.n3656 3.49141
R11800 gnd.n3643 gnd.n3624 3.49141
R11801 gnd.n3611 gnd.n3592 3.49141
R11802 gnd.n3579 gnd.n3560 3.49141
R11803 gnd.n3548 gnd.n3529 3.49141
R11804 gnd.n5720 gnd.n5719 3.29747
R11805 gnd.n5719 gnd.n5718 3.29747
R11806 gnd.n392 gnd.n328 3.29747
R11807 gnd.n387 gnd.n328 3.29747
R11808 gnd.n4206 gnd.n4205 3.29747
R11809 gnd.n4205 gnd.n4204 3.29747
R11810 gnd.n6052 gnd.n6051 3.29747
R11811 gnd.n6051 gnd.n6050 3.29747
R11812 gnd.t71 gnd.n5939 3.18706
R11813 gnd.n5396 gnd.t120 3.18706
R11814 gnd.n144 gnd.n136 3.18706
R11815 gnd.n2807 gnd.t19 2.8684
R11816 gnd.n2710 gnd.t227 2.82907
R11817 gnd.n2710 gnd.t290 2.82907
R11818 gnd.n2712 gnd.t206 2.82907
R11819 gnd.n2712 gnd.t241 2.82907
R11820 gnd.n2714 gnd.t259 2.82907
R11821 gnd.n2714 gnd.t247 2.82907
R11822 gnd.n2716 gnd.t245 2.82907
R11823 gnd.n2716 gnd.t236 2.82907
R11824 gnd.n2718 gnd.t250 2.82907
R11825 gnd.n2718 gnd.t276 2.82907
R11826 gnd.n2675 gnd.t252 2.82907
R11827 gnd.n2675 gnd.t269 2.82907
R11828 gnd.n2677 gnd.t275 2.82907
R11829 gnd.n2677 gnd.t228 2.82907
R11830 gnd.n2679 gnd.t267 2.82907
R11831 gnd.n2679 gnd.t265 2.82907
R11832 gnd.n2681 gnd.t299 2.82907
R11833 gnd.n2681 gnd.t278 2.82907
R11834 gnd.n2683 gnd.t234 2.82907
R11835 gnd.n2683 gnd.t272 2.82907
R11836 gnd.n2686 gnd.t301 2.82907
R11837 gnd.n2686 gnd.t211 2.82907
R11838 gnd.n2688 gnd.t212 2.82907
R11839 gnd.n2688 gnd.t195 2.82907
R11840 gnd.n2690 gnd.t274 2.82907
R11841 gnd.n2690 gnd.t302 2.82907
R11842 gnd.n2692 gnd.t297 2.82907
R11843 gnd.n2692 gnd.t219 2.82907
R11844 gnd.n2694 gnd.t277 2.82907
R11845 gnd.n2694 gnd.t256 2.82907
R11846 gnd.n2698 gnd.t264 2.82907
R11847 gnd.n2698 gnd.t230 2.82907
R11848 gnd.n2700 gnd.t251 2.82907
R11849 gnd.n2700 gnd.t280 2.82907
R11850 gnd.n2702 gnd.t296 2.82907
R11851 gnd.n2702 gnd.t287 2.82907
R11852 gnd.n2704 gnd.t285 2.82907
R11853 gnd.n2704 gnd.t271 2.82907
R11854 gnd.n2706 gnd.t289 2.82907
R11855 gnd.n2706 gnd.t225 2.82907
R11856 gnd.n59 gnd.t254 2.82907
R11857 gnd.n59 gnd.t235 2.82907
R11858 gnd.n57 gnd.t202 2.82907
R11859 gnd.n57 gnd.t223 2.82907
R11860 gnd.n55 gnd.t217 2.82907
R11861 gnd.n55 gnd.t238 2.82907
R11862 gnd.n53 gnd.t221 2.82907
R11863 gnd.n53 gnd.t284 2.82907
R11864 gnd.n51 gnd.t263 2.82907
R11865 gnd.n51 gnd.t199 2.82907
R11866 gnd.n24 gnd.t304 2.82907
R11867 gnd.n24 gnd.t215 2.82907
R11868 gnd.n22 gnd.t209 2.82907
R11869 gnd.n22 gnd.t214 2.82907
R11870 gnd.n20 gnd.t286 2.82907
R11871 gnd.n20 gnd.t261 2.82907
R11872 gnd.n18 gnd.t249 2.82907
R11873 gnd.n18 gnd.t193 2.82907
R11874 gnd.n16 gnd.t295 2.82907
R11875 gnd.n16 gnd.t239 2.82907
R11876 gnd.n35 gnd.t266 2.82907
R11877 gnd.n35 gnd.t192 2.82907
R11878 gnd.n33 gnd.t190 2.82907
R11879 gnd.n33 gnd.t281 2.82907
R11880 gnd.n31 gnd.t288 2.82907
R11881 gnd.n31 gnd.t294 2.82907
R11882 gnd.n29 gnd.t293 2.82907
R11883 gnd.n29 gnd.t188 2.82907
R11884 gnd.n27 gnd.t186 2.82907
R11885 gnd.n27 gnd.t203 2.82907
R11886 gnd.n47 gnd.t292 2.82907
R11887 gnd.n47 gnd.t270 2.82907
R11888 gnd.n45 gnd.t248 2.82907
R11889 gnd.n45 gnd.t260 2.82907
R11890 gnd.n43 gnd.t262 2.82907
R11891 gnd.n43 gnd.t273 2.82907
R11892 gnd.n41 gnd.t255 2.82907
R11893 gnd.n41 gnd.t229 2.82907
R11894 gnd.n39 gnd.t303 2.82907
R11895 gnd.n39 gnd.t243 2.82907
R11896 gnd.n3767 gnd.n3766 2.71565
R11897 gnd.n3735 gnd.n3734 2.71565
R11898 gnd.n3703 gnd.n3702 2.71565
R11899 gnd.n3672 gnd.n3671 2.71565
R11900 gnd.n3640 gnd.n3639 2.71565
R11901 gnd.n3608 gnd.n3607 2.71565
R11902 gnd.n3576 gnd.n3575 2.71565
R11903 gnd.n3545 gnd.n3544 2.71565
R11904 gnd.n4823 gnd.n4822 2.54975
R11905 gnd.n4837 gnd.t24 2.54975
R11906 gnd.n4852 gnd.n4851 2.54975
R11907 gnd.t29 gnd.n2176 2.54975
R11908 gnd.n2168 gnd.n2162 2.54975
R11909 gnd.n4987 gnd.t1 2.54975
R11910 gnd.n5060 gnd.n2121 2.54975
R11911 gnd.n5119 gnd.n2088 2.54975
R11912 gnd.t30 gnd.n5209 2.54975
R11913 gnd.n2044 gnd.n2043 2.54975
R11914 gnd.n5275 gnd.t15 2.54975
R11915 gnd.n5304 gnd.n5303 2.54975
R11916 gnd.n5234 gnd.t17 2.54975
R11917 gnd.n5377 gnd.n1939 2.54975
R11918 gnd.n3301 gnd.n2723 2.27742
R11919 gnd.n3301 gnd.n2674 2.27742
R11920 gnd.n3301 gnd.n2673 2.27742
R11921 gnd.n3301 gnd.n2672 2.27742
R11922 gnd.n7020 gnd.n81 2.27742
R11923 gnd.n7020 gnd.n80 2.27742
R11924 gnd.n7020 gnd.n79 2.27742
R11925 gnd.n7020 gnd.n74 2.27742
R11926 gnd.n7021 gnd.n7020 2.27742
R11927 gnd.n2356 gnd.n1058 2.27742
R11928 gnd.n4336 gnd.n1058 2.27742
R11929 gnd.n2337 gnd.n1058 2.27742
R11930 gnd.n4363 gnd.n1058 2.27742
R11931 gnd.n1058 gnd.n1057 2.27742
R11932 gnd.n3155 gnd.t126 2.23109
R11933 gnd.n2778 gnd.t58 2.23109
R11934 gnd.n4909 gnd.t38 2.23109
R11935 gnd.n5175 gnd.t326 2.23109
R11936 gnd.n3763 gnd.n3753 1.93989
R11937 gnd.n3731 gnd.n3721 1.93989
R11938 gnd.n3699 gnd.n3689 1.93989
R11939 gnd.n3668 gnd.n3658 1.93989
R11940 gnd.n3636 gnd.n3626 1.93989
R11941 gnd.n3604 gnd.n3594 1.93989
R11942 gnd.n3572 gnd.n3562 1.93989
R11943 gnd.n3541 gnd.n3531 1.93989
R11944 gnd.t310 gnd.n3166 1.59378
R11945 gnd.n3345 gnd.t51 1.59378
R11946 gnd.n2607 gnd.t25 1.59378
R11947 gnd.t68 gnd.n5959 1.27512
R11948 gnd.n5959 gnd.n5958 1.27512
R11949 gnd.n1377 gnd.n1371 1.27512
R11950 gnd.n4947 gnd.n2185 1.27512
R11951 gnd.n4967 gnd.n2172 1.27512
R11952 gnd.n5090 gnd.n5089 1.27512
R11953 gnd.n5112 gnd.n2094 1.27512
R11954 gnd.n2032 gnd.n2017 1.27512
R11955 gnd.n5284 gnd.n5283 1.27512
R11956 gnd.n5387 gnd.n1931 1.27512
R11957 gnd.n5404 gnd.n5403 1.27512
R11958 gnd.n3008 gnd.n3000 1.16414
R11959 gnd.n3825 gnd.n2510 1.16414
R11960 gnd.n3762 gnd.n3755 1.16414
R11961 gnd.n3730 gnd.n3723 1.16414
R11962 gnd.n3698 gnd.n3691 1.16414
R11963 gnd.n3667 gnd.n3660 1.16414
R11964 gnd.n3635 gnd.n3628 1.16414
R11965 gnd.n3603 gnd.n3596 1.16414
R11966 gnd.n3571 gnd.n3564 1.16414
R11967 gnd.n3540 gnd.n3533 1.16414
R11968 gnd.n5702 gnd.n5701 0.970197
R11969 gnd.n6034 gnd.n1211 0.970197
R11970 gnd.n3746 gnd.n3714 0.962709
R11971 gnd.n3778 gnd.n3746 0.962709
R11972 gnd.n3619 gnd.n3587 0.962709
R11973 gnd.n3651 gnd.n3619 0.962709
R11974 gnd.n3254 gnd.t40 0.956468
R11975 gnd.n3419 gnd.t9 0.956468
R11976 gnd.n4291 gnd.t233 0.956468
R11977 gnd.n6116 gnd.t210 0.956468
R11978 gnd.n4776 gnd.t319 0.956468
R11979 gnd.n4823 gnd.t306 0.956468
R11980 gnd.n5377 gnd.t22 0.956468
R11981 gnd.t42 gnd.n1790 0.956468
R11982 gnd.n5601 gnd.t185 0.956468
R11983 gnd.n124 gnd.t191 0.956468
R11984 gnd.n2 gnd.n1 0.672012
R11985 gnd.n3 gnd.n2 0.672012
R11986 gnd.n4 gnd.n3 0.672012
R11987 gnd.n5 gnd.n4 0.672012
R11988 gnd.n6 gnd.n5 0.672012
R11989 gnd.n7 gnd.n6 0.672012
R11990 gnd.n9 gnd.n8 0.672012
R11991 gnd.n10 gnd.n9 0.672012
R11992 gnd.n11 gnd.n10 0.672012
R11993 gnd.n12 gnd.n11 0.672012
R11994 gnd.n13 gnd.n12 0.672012
R11995 gnd.n14 gnd.n13 0.672012
R11996 gnd.n5952 gnd.t102 0.637812
R11997 gnd.n4864 gnd.t0 0.637812
R11998 gnd.n5031 gnd.t31 0.637812
R11999 gnd.n5120 gnd.t16 0.637812
R12000 gnd.t21 gnd.n1979 0.637812
R12001 gnd.n5396 gnd.t92 0.637812
R12002 gnd.n2720 gnd.n2719 0.573776
R12003 gnd.n2719 gnd.n2717 0.573776
R12004 gnd.n2717 gnd.n2715 0.573776
R12005 gnd.n2715 gnd.n2713 0.573776
R12006 gnd.n2713 gnd.n2711 0.573776
R12007 gnd.n2685 gnd.n2684 0.573776
R12008 gnd.n2684 gnd.n2682 0.573776
R12009 gnd.n2682 gnd.n2680 0.573776
R12010 gnd.n2680 gnd.n2678 0.573776
R12011 gnd.n2678 gnd.n2676 0.573776
R12012 gnd.n2696 gnd.n2695 0.573776
R12013 gnd.n2695 gnd.n2693 0.573776
R12014 gnd.n2693 gnd.n2691 0.573776
R12015 gnd.n2691 gnd.n2689 0.573776
R12016 gnd.n2689 gnd.n2687 0.573776
R12017 gnd.n2708 gnd.n2707 0.573776
R12018 gnd.n2707 gnd.n2705 0.573776
R12019 gnd.n2705 gnd.n2703 0.573776
R12020 gnd.n2703 gnd.n2701 0.573776
R12021 gnd.n2701 gnd.n2699 0.573776
R12022 gnd.n54 gnd.n52 0.573776
R12023 gnd.n56 gnd.n54 0.573776
R12024 gnd.n58 gnd.n56 0.573776
R12025 gnd.n60 gnd.n58 0.573776
R12026 gnd.n61 gnd.n60 0.573776
R12027 gnd.n19 gnd.n17 0.573776
R12028 gnd.n21 gnd.n19 0.573776
R12029 gnd.n23 gnd.n21 0.573776
R12030 gnd.n25 gnd.n23 0.573776
R12031 gnd.n26 gnd.n25 0.573776
R12032 gnd.n30 gnd.n28 0.573776
R12033 gnd.n32 gnd.n30 0.573776
R12034 gnd.n34 gnd.n32 0.573776
R12035 gnd.n36 gnd.n34 0.573776
R12036 gnd.n37 gnd.n36 0.573776
R12037 gnd.n42 gnd.n40 0.573776
R12038 gnd.n44 gnd.n42 0.573776
R12039 gnd.n46 gnd.n44 0.573776
R12040 gnd.n48 gnd.n46 0.573776
R12041 gnd.n49 gnd.n48 0.573776
R12042 gnd gnd.n0 0.551497
R12043 gnd.n248 gnd.n247 0.532512
R12044 gnd.n4085 gnd.n4083 0.532512
R12045 gnd.n344 gnd.n160 0.497451
R12046 gnd.n6088 gnd.n6087 0.497451
R12047 gnd.n1684 gnd.n1603 0.497451
R12048 gnd.n3945 gnd.n2427 0.497451
R12049 gnd.n5826 gnd.n1485 0.489829
R12050 gnd.n4735 gnd.n4734 0.489829
R12051 gnd.n4758 gnd.n2262 0.489829
R12052 gnd.n5820 gnd.n5819 0.489829
R12053 gnd.n3481 gnd.n2514 0.486781
R12054 gnd.n3057 gnd.n3056 0.48678
R12055 gnd.n3799 gnd.n2468 0.480683
R12056 gnd.n3141 gnd.n3140 0.480683
R12057 gnd.n7032 gnd.n7031 0.470187
R12058 gnd.n7020 gnd.n78 0.420375
R12059 gnd.n4399 gnd.n1058 0.420375
R12060 gnd.n6313 gnd.n6312 0.416659
R12061 gnd.n6635 gnd.n6634 0.416659
R12062 gnd.n4519 gnd.n4510 0.388379
R12063 gnd.n3759 gnd.n3758 0.388379
R12064 gnd.n3727 gnd.n3726 0.388379
R12065 gnd.n3695 gnd.n3694 0.388379
R12066 gnd.n3664 gnd.n3663 0.388379
R12067 gnd.n3632 gnd.n3631 0.388379
R12068 gnd.n3600 gnd.n3599 0.388379
R12069 gnd.n3568 gnd.n3567 0.388379
R12070 gnd.n3537 gnd.n3536 0.388379
R12071 gnd.n5764 gnd.n1551 0.388379
R12072 gnd.n7032 gnd.n15 0.374463
R12073 gnd.n2569 gnd.t18 0.319156
R12074 gnd.n4332 gnd.t218 0.319156
R12075 gnd.t205 gnd.n6140 0.319156
R12076 gnd.n4984 gnd.t53 0.319156
R12077 gnd.t20 gnd.t308 0.319156
R12078 gnd.t34 gnd.t27 0.319156
R12079 gnd.t312 gnd.n2040 0.319156
R12080 gnd.n6902 gnd.t187 0.319156
R12081 gnd.n85 gnd.t189 0.319156
R12082 gnd.n2975 gnd.n2953 0.311721
R12083 gnd.n4720 gnd.n2290 0.302329
R12084 gnd.n5535 gnd.n5534 0.302329
R12085 gnd gnd.n7032 0.295112
R12086 gnd.n493 gnd.n280 0.293183
R12087 gnd.n4123 gnd.n4122 0.293183
R12088 gnd.n6846 gnd.n78 0.280988
R12089 gnd.n4399 gnd.n1048 0.280988
R12090 gnd.n3870 gnd.n3869 0.268793
R12091 gnd.n493 gnd.n492 0.258122
R12092 gnd.n5640 gnd.n1504 0.258122
R12093 gnd.n4671 gnd.n4670 0.258122
R12094 gnd.n4124 gnd.n4123 0.258122
R12095 gnd.n3869 gnd.n3868 0.241354
R12096 gnd.n1633 gnd.n1630 0.229039
R12097 gnd.n1634 gnd.n1633 0.229039
R12098 gnd.n1213 gnd.n1210 0.229039
R12099 gnd.n4595 gnd.n1213 0.229039
R12100 gnd.n3129 gnd.n2928 0.206293
R12101 gnd.n3776 gnd.n3748 0.155672
R12102 gnd.n3769 gnd.n3748 0.155672
R12103 gnd.n3769 gnd.n3768 0.155672
R12104 gnd.n3768 gnd.n3752 0.155672
R12105 gnd.n3761 gnd.n3752 0.155672
R12106 gnd.n3761 gnd.n3760 0.155672
R12107 gnd.n3744 gnd.n3716 0.155672
R12108 gnd.n3737 gnd.n3716 0.155672
R12109 gnd.n3737 gnd.n3736 0.155672
R12110 gnd.n3736 gnd.n3720 0.155672
R12111 gnd.n3729 gnd.n3720 0.155672
R12112 gnd.n3729 gnd.n3728 0.155672
R12113 gnd.n3712 gnd.n3684 0.155672
R12114 gnd.n3705 gnd.n3684 0.155672
R12115 gnd.n3705 gnd.n3704 0.155672
R12116 gnd.n3704 gnd.n3688 0.155672
R12117 gnd.n3697 gnd.n3688 0.155672
R12118 gnd.n3697 gnd.n3696 0.155672
R12119 gnd.n3681 gnd.n3653 0.155672
R12120 gnd.n3674 gnd.n3653 0.155672
R12121 gnd.n3674 gnd.n3673 0.155672
R12122 gnd.n3673 gnd.n3657 0.155672
R12123 gnd.n3666 gnd.n3657 0.155672
R12124 gnd.n3666 gnd.n3665 0.155672
R12125 gnd.n3649 gnd.n3621 0.155672
R12126 gnd.n3642 gnd.n3621 0.155672
R12127 gnd.n3642 gnd.n3641 0.155672
R12128 gnd.n3641 gnd.n3625 0.155672
R12129 gnd.n3634 gnd.n3625 0.155672
R12130 gnd.n3634 gnd.n3633 0.155672
R12131 gnd.n3617 gnd.n3589 0.155672
R12132 gnd.n3610 gnd.n3589 0.155672
R12133 gnd.n3610 gnd.n3609 0.155672
R12134 gnd.n3609 gnd.n3593 0.155672
R12135 gnd.n3602 gnd.n3593 0.155672
R12136 gnd.n3602 gnd.n3601 0.155672
R12137 gnd.n3585 gnd.n3557 0.155672
R12138 gnd.n3578 gnd.n3557 0.155672
R12139 gnd.n3578 gnd.n3577 0.155672
R12140 gnd.n3577 gnd.n3561 0.155672
R12141 gnd.n3570 gnd.n3561 0.155672
R12142 gnd.n3570 gnd.n3569 0.155672
R12143 gnd.n3554 gnd.n3526 0.155672
R12144 gnd.n3547 gnd.n3526 0.155672
R12145 gnd.n3547 gnd.n3546 0.155672
R12146 gnd.n3546 gnd.n3530 0.155672
R12147 gnd.n3539 gnd.n3530 0.155672
R12148 gnd.n3539 gnd.n3538 0.155672
R12149 gnd.n3901 gnd.n2468 0.152939
R12150 gnd.n3901 gnd.n3900 0.152939
R12151 gnd.n3900 gnd.n3899 0.152939
R12152 gnd.n3899 gnd.n2470 0.152939
R12153 gnd.n2471 gnd.n2470 0.152939
R12154 gnd.n2472 gnd.n2471 0.152939
R12155 gnd.n2473 gnd.n2472 0.152939
R12156 gnd.n2474 gnd.n2473 0.152939
R12157 gnd.n2475 gnd.n2474 0.152939
R12158 gnd.n2476 gnd.n2475 0.152939
R12159 gnd.n2477 gnd.n2476 0.152939
R12160 gnd.n2478 gnd.n2477 0.152939
R12161 gnd.n2479 gnd.n2478 0.152939
R12162 gnd.n2480 gnd.n2479 0.152939
R12163 gnd.n3871 gnd.n2480 0.152939
R12164 gnd.n3871 gnd.n3870 0.152939
R12165 gnd.n3142 gnd.n3141 0.152939
R12166 gnd.n3142 gnd.n2846 0.152939
R12167 gnd.n3170 gnd.n2846 0.152939
R12168 gnd.n3171 gnd.n3170 0.152939
R12169 gnd.n3172 gnd.n3171 0.152939
R12170 gnd.n3173 gnd.n3172 0.152939
R12171 gnd.n3173 gnd.n2818 0.152939
R12172 gnd.n3200 gnd.n2818 0.152939
R12173 gnd.n3201 gnd.n3200 0.152939
R12174 gnd.n3202 gnd.n3201 0.152939
R12175 gnd.n3202 gnd.n2796 0.152939
R12176 gnd.n3231 gnd.n2796 0.152939
R12177 gnd.n3232 gnd.n3231 0.152939
R12178 gnd.n3233 gnd.n3232 0.152939
R12179 gnd.n3234 gnd.n3233 0.152939
R12180 gnd.n3236 gnd.n3234 0.152939
R12181 gnd.n3236 gnd.n3235 0.152939
R12182 gnd.n3235 gnd.n2745 0.152939
R12183 gnd.n2746 gnd.n2745 0.152939
R12184 gnd.n2747 gnd.n2746 0.152939
R12185 gnd.n2766 gnd.n2747 0.152939
R12186 gnd.n2767 gnd.n2766 0.152939
R12187 gnd.n2767 gnd.n2665 0.152939
R12188 gnd.n3326 gnd.n2665 0.152939
R12189 gnd.n3327 gnd.n3326 0.152939
R12190 gnd.n3328 gnd.n3327 0.152939
R12191 gnd.n3329 gnd.n3328 0.152939
R12192 gnd.n3329 gnd.n2638 0.152939
R12193 gnd.n3366 gnd.n2638 0.152939
R12194 gnd.n3367 gnd.n3366 0.152939
R12195 gnd.n3368 gnd.n3367 0.152939
R12196 gnd.n3369 gnd.n3368 0.152939
R12197 gnd.n3369 gnd.n2611 0.152939
R12198 gnd.n3411 gnd.n2611 0.152939
R12199 gnd.n3412 gnd.n3411 0.152939
R12200 gnd.n3413 gnd.n3412 0.152939
R12201 gnd.n3414 gnd.n3413 0.152939
R12202 gnd.n3414 gnd.n2583 0.152939
R12203 gnd.n3451 gnd.n2583 0.152939
R12204 gnd.n3452 gnd.n3451 0.152939
R12205 gnd.n3453 gnd.n3452 0.152939
R12206 gnd.n3454 gnd.n3453 0.152939
R12207 gnd.n3454 gnd.n2556 0.152939
R12208 gnd.n3500 gnd.n2556 0.152939
R12209 gnd.n3501 gnd.n3500 0.152939
R12210 gnd.n3502 gnd.n3501 0.152939
R12211 gnd.n3503 gnd.n3502 0.152939
R12212 gnd.n3503 gnd.n2529 0.152939
R12213 gnd.n3795 gnd.n2529 0.152939
R12214 gnd.n3796 gnd.n3795 0.152939
R12215 gnd.n3797 gnd.n3796 0.152939
R12216 gnd.n3798 gnd.n3797 0.152939
R12217 gnd.n3799 gnd.n3798 0.152939
R12218 gnd.n3140 gnd.n2870 0.152939
R12219 gnd.n2891 gnd.n2870 0.152939
R12220 gnd.n2892 gnd.n2891 0.152939
R12221 gnd.n2898 gnd.n2892 0.152939
R12222 gnd.n2899 gnd.n2898 0.152939
R12223 gnd.n2900 gnd.n2899 0.152939
R12224 gnd.n2900 gnd.n2889 0.152939
R12225 gnd.n2908 gnd.n2889 0.152939
R12226 gnd.n2909 gnd.n2908 0.152939
R12227 gnd.n2910 gnd.n2909 0.152939
R12228 gnd.n2910 gnd.n2887 0.152939
R12229 gnd.n2918 gnd.n2887 0.152939
R12230 gnd.n2919 gnd.n2918 0.152939
R12231 gnd.n2920 gnd.n2919 0.152939
R12232 gnd.n2920 gnd.n2885 0.152939
R12233 gnd.n2928 gnd.n2885 0.152939
R12234 gnd.n3868 gnd.n2485 0.152939
R12235 gnd.n2487 gnd.n2485 0.152939
R12236 gnd.n2488 gnd.n2487 0.152939
R12237 gnd.n2489 gnd.n2488 0.152939
R12238 gnd.n2490 gnd.n2489 0.152939
R12239 gnd.n2491 gnd.n2490 0.152939
R12240 gnd.n2492 gnd.n2491 0.152939
R12241 gnd.n2493 gnd.n2492 0.152939
R12242 gnd.n2494 gnd.n2493 0.152939
R12243 gnd.n2495 gnd.n2494 0.152939
R12244 gnd.n2496 gnd.n2495 0.152939
R12245 gnd.n2497 gnd.n2496 0.152939
R12246 gnd.n2498 gnd.n2497 0.152939
R12247 gnd.n2499 gnd.n2498 0.152939
R12248 gnd.n2500 gnd.n2499 0.152939
R12249 gnd.n2501 gnd.n2500 0.152939
R12250 gnd.n2502 gnd.n2501 0.152939
R12251 gnd.n2503 gnd.n2502 0.152939
R12252 gnd.n2504 gnd.n2503 0.152939
R12253 gnd.n2505 gnd.n2504 0.152939
R12254 gnd.n2506 gnd.n2505 0.152939
R12255 gnd.n2507 gnd.n2506 0.152939
R12256 gnd.n2511 gnd.n2507 0.152939
R12257 gnd.n2512 gnd.n2511 0.152939
R12258 gnd.n2513 gnd.n2512 0.152939
R12259 gnd.n2514 gnd.n2513 0.152939
R12260 gnd.n3303 gnd.n3302 0.152939
R12261 gnd.n3304 gnd.n3303 0.152939
R12262 gnd.n3305 gnd.n3304 0.152939
R12263 gnd.n3306 gnd.n3305 0.152939
R12264 gnd.n3307 gnd.n3306 0.152939
R12265 gnd.n3308 gnd.n3307 0.152939
R12266 gnd.n3308 gnd.n2619 0.152939
R12267 gnd.n3387 gnd.n2619 0.152939
R12268 gnd.n3388 gnd.n3387 0.152939
R12269 gnd.n3389 gnd.n3388 0.152939
R12270 gnd.n3390 gnd.n3389 0.152939
R12271 gnd.n3391 gnd.n3390 0.152939
R12272 gnd.n3392 gnd.n3391 0.152939
R12273 gnd.n3393 gnd.n3392 0.152939
R12274 gnd.n3394 gnd.n3393 0.152939
R12275 gnd.n3395 gnd.n3394 0.152939
R12276 gnd.n3395 gnd.n2563 0.152939
R12277 gnd.n3472 gnd.n2563 0.152939
R12278 gnd.n3473 gnd.n3472 0.152939
R12279 gnd.n3474 gnd.n3473 0.152939
R12280 gnd.n3475 gnd.n3474 0.152939
R12281 gnd.n3476 gnd.n3475 0.152939
R12282 gnd.n3477 gnd.n3476 0.152939
R12283 gnd.n3478 gnd.n3477 0.152939
R12284 gnd.n3479 gnd.n3478 0.152939
R12285 gnd.n3480 gnd.n3479 0.152939
R12286 gnd.n3482 gnd.n3480 0.152939
R12287 gnd.n3482 gnd.n3481 0.152939
R12288 gnd.n3058 gnd.n3057 0.152939
R12289 gnd.n3058 gnd.n2948 0.152939
R12290 gnd.n3073 gnd.n2948 0.152939
R12291 gnd.n3074 gnd.n3073 0.152939
R12292 gnd.n3075 gnd.n3074 0.152939
R12293 gnd.n3075 gnd.n2936 0.152939
R12294 gnd.n3089 gnd.n2936 0.152939
R12295 gnd.n3090 gnd.n3089 0.152939
R12296 gnd.n3091 gnd.n3090 0.152939
R12297 gnd.n3092 gnd.n3091 0.152939
R12298 gnd.n3093 gnd.n3092 0.152939
R12299 gnd.n3094 gnd.n3093 0.152939
R12300 gnd.n3095 gnd.n3094 0.152939
R12301 gnd.n3096 gnd.n3095 0.152939
R12302 gnd.n3097 gnd.n3096 0.152939
R12303 gnd.n3098 gnd.n3097 0.152939
R12304 gnd.n3099 gnd.n3098 0.152939
R12305 gnd.n3100 gnd.n3099 0.152939
R12306 gnd.n3101 gnd.n3100 0.152939
R12307 gnd.n3102 gnd.n3101 0.152939
R12308 gnd.n3103 gnd.n3102 0.152939
R12309 gnd.n3103 gnd.n2802 0.152939
R12310 gnd.n3220 gnd.n2802 0.152939
R12311 gnd.n3221 gnd.n3220 0.152939
R12312 gnd.n3222 gnd.n3221 0.152939
R12313 gnd.n3223 gnd.n3222 0.152939
R12314 gnd.n3223 gnd.n2724 0.152939
R12315 gnd.n3300 gnd.n2724 0.152939
R12316 gnd.n2976 gnd.n2975 0.152939
R12317 gnd.n2977 gnd.n2976 0.152939
R12318 gnd.n2978 gnd.n2977 0.152939
R12319 gnd.n2979 gnd.n2978 0.152939
R12320 gnd.n2980 gnd.n2979 0.152939
R12321 gnd.n2981 gnd.n2980 0.152939
R12322 gnd.n2982 gnd.n2981 0.152939
R12323 gnd.n2983 gnd.n2982 0.152939
R12324 gnd.n2984 gnd.n2983 0.152939
R12325 gnd.n2985 gnd.n2984 0.152939
R12326 gnd.n2986 gnd.n2985 0.152939
R12327 gnd.n2987 gnd.n2986 0.152939
R12328 gnd.n2988 gnd.n2987 0.152939
R12329 gnd.n2989 gnd.n2988 0.152939
R12330 gnd.n2990 gnd.n2989 0.152939
R12331 gnd.n2991 gnd.n2990 0.152939
R12332 gnd.n2992 gnd.n2991 0.152939
R12333 gnd.n2993 gnd.n2992 0.152939
R12334 gnd.n2994 gnd.n2993 0.152939
R12335 gnd.n2995 gnd.n2994 0.152939
R12336 gnd.n2996 gnd.n2995 0.152939
R12337 gnd.n2997 gnd.n2996 0.152939
R12338 gnd.n3001 gnd.n2997 0.152939
R12339 gnd.n3002 gnd.n3001 0.152939
R12340 gnd.n3002 gnd.n2959 0.152939
R12341 gnd.n3056 gnd.n2959 0.152939
R12342 gnd.n6314 gnd.n6313 0.152939
R12343 gnd.n6314 gnd.n875 0.152939
R12344 gnd.n6322 gnd.n875 0.152939
R12345 gnd.n6323 gnd.n6322 0.152939
R12346 gnd.n6324 gnd.n6323 0.152939
R12347 gnd.n6324 gnd.n869 0.152939
R12348 gnd.n6332 gnd.n869 0.152939
R12349 gnd.n6333 gnd.n6332 0.152939
R12350 gnd.n6334 gnd.n6333 0.152939
R12351 gnd.n6334 gnd.n863 0.152939
R12352 gnd.n6342 gnd.n863 0.152939
R12353 gnd.n6343 gnd.n6342 0.152939
R12354 gnd.n6344 gnd.n6343 0.152939
R12355 gnd.n6344 gnd.n857 0.152939
R12356 gnd.n6352 gnd.n857 0.152939
R12357 gnd.n6353 gnd.n6352 0.152939
R12358 gnd.n6354 gnd.n6353 0.152939
R12359 gnd.n6354 gnd.n851 0.152939
R12360 gnd.n6362 gnd.n851 0.152939
R12361 gnd.n6363 gnd.n6362 0.152939
R12362 gnd.n6364 gnd.n6363 0.152939
R12363 gnd.n6364 gnd.n845 0.152939
R12364 gnd.n6372 gnd.n845 0.152939
R12365 gnd.n6373 gnd.n6372 0.152939
R12366 gnd.n6374 gnd.n6373 0.152939
R12367 gnd.n6374 gnd.n839 0.152939
R12368 gnd.n6382 gnd.n839 0.152939
R12369 gnd.n6383 gnd.n6382 0.152939
R12370 gnd.n6384 gnd.n6383 0.152939
R12371 gnd.n6384 gnd.n833 0.152939
R12372 gnd.n6392 gnd.n833 0.152939
R12373 gnd.n6393 gnd.n6392 0.152939
R12374 gnd.n6394 gnd.n6393 0.152939
R12375 gnd.n6394 gnd.n827 0.152939
R12376 gnd.n6402 gnd.n827 0.152939
R12377 gnd.n6403 gnd.n6402 0.152939
R12378 gnd.n6404 gnd.n6403 0.152939
R12379 gnd.n6404 gnd.n821 0.152939
R12380 gnd.n6412 gnd.n821 0.152939
R12381 gnd.n6413 gnd.n6412 0.152939
R12382 gnd.n6414 gnd.n6413 0.152939
R12383 gnd.n6414 gnd.n815 0.152939
R12384 gnd.n6422 gnd.n815 0.152939
R12385 gnd.n6423 gnd.n6422 0.152939
R12386 gnd.n6424 gnd.n6423 0.152939
R12387 gnd.n6424 gnd.n809 0.152939
R12388 gnd.n6432 gnd.n809 0.152939
R12389 gnd.n6433 gnd.n6432 0.152939
R12390 gnd.n6434 gnd.n6433 0.152939
R12391 gnd.n6434 gnd.n803 0.152939
R12392 gnd.n6442 gnd.n803 0.152939
R12393 gnd.n6443 gnd.n6442 0.152939
R12394 gnd.n6444 gnd.n6443 0.152939
R12395 gnd.n6444 gnd.n797 0.152939
R12396 gnd.n6452 gnd.n797 0.152939
R12397 gnd.n6453 gnd.n6452 0.152939
R12398 gnd.n6454 gnd.n6453 0.152939
R12399 gnd.n6454 gnd.n791 0.152939
R12400 gnd.n6462 gnd.n791 0.152939
R12401 gnd.n6463 gnd.n6462 0.152939
R12402 gnd.n6464 gnd.n6463 0.152939
R12403 gnd.n6464 gnd.n785 0.152939
R12404 gnd.n6472 gnd.n785 0.152939
R12405 gnd.n6473 gnd.n6472 0.152939
R12406 gnd.n6474 gnd.n6473 0.152939
R12407 gnd.n6474 gnd.n779 0.152939
R12408 gnd.n6482 gnd.n779 0.152939
R12409 gnd.n6483 gnd.n6482 0.152939
R12410 gnd.n6484 gnd.n6483 0.152939
R12411 gnd.n6484 gnd.n773 0.152939
R12412 gnd.n6492 gnd.n773 0.152939
R12413 gnd.n6493 gnd.n6492 0.152939
R12414 gnd.n6494 gnd.n6493 0.152939
R12415 gnd.n6494 gnd.n767 0.152939
R12416 gnd.n6502 gnd.n767 0.152939
R12417 gnd.n6503 gnd.n6502 0.152939
R12418 gnd.n6504 gnd.n6503 0.152939
R12419 gnd.n6504 gnd.n761 0.152939
R12420 gnd.n6512 gnd.n761 0.152939
R12421 gnd.n6513 gnd.n6512 0.152939
R12422 gnd.n6514 gnd.n6513 0.152939
R12423 gnd.n6514 gnd.n755 0.152939
R12424 gnd.n6522 gnd.n755 0.152939
R12425 gnd.n6523 gnd.n6522 0.152939
R12426 gnd.n6524 gnd.n6523 0.152939
R12427 gnd.n6524 gnd.n749 0.152939
R12428 gnd.n6532 gnd.n749 0.152939
R12429 gnd.n6533 gnd.n6532 0.152939
R12430 gnd.n6534 gnd.n6533 0.152939
R12431 gnd.n6534 gnd.n743 0.152939
R12432 gnd.n6542 gnd.n743 0.152939
R12433 gnd.n6543 gnd.n6542 0.152939
R12434 gnd.n6544 gnd.n6543 0.152939
R12435 gnd.n6544 gnd.n737 0.152939
R12436 gnd.n6552 gnd.n737 0.152939
R12437 gnd.n6553 gnd.n6552 0.152939
R12438 gnd.n6554 gnd.n6553 0.152939
R12439 gnd.n6554 gnd.n731 0.152939
R12440 gnd.n6562 gnd.n731 0.152939
R12441 gnd.n6563 gnd.n6562 0.152939
R12442 gnd.n6564 gnd.n6563 0.152939
R12443 gnd.n6564 gnd.n725 0.152939
R12444 gnd.n6572 gnd.n725 0.152939
R12445 gnd.n6573 gnd.n6572 0.152939
R12446 gnd.n6574 gnd.n6573 0.152939
R12447 gnd.n6574 gnd.n719 0.152939
R12448 gnd.n6582 gnd.n719 0.152939
R12449 gnd.n6583 gnd.n6582 0.152939
R12450 gnd.n6584 gnd.n6583 0.152939
R12451 gnd.n6584 gnd.n713 0.152939
R12452 gnd.n6592 gnd.n713 0.152939
R12453 gnd.n6593 gnd.n6592 0.152939
R12454 gnd.n6594 gnd.n6593 0.152939
R12455 gnd.n6594 gnd.n707 0.152939
R12456 gnd.n6602 gnd.n707 0.152939
R12457 gnd.n6603 gnd.n6602 0.152939
R12458 gnd.n6604 gnd.n6603 0.152939
R12459 gnd.n6604 gnd.n701 0.152939
R12460 gnd.n6612 gnd.n701 0.152939
R12461 gnd.n6613 gnd.n6612 0.152939
R12462 gnd.n6614 gnd.n6613 0.152939
R12463 gnd.n6614 gnd.n695 0.152939
R12464 gnd.n6622 gnd.n695 0.152939
R12465 gnd.n6623 gnd.n6622 0.152939
R12466 gnd.n6625 gnd.n6623 0.152939
R12467 gnd.n6625 gnd.n6624 0.152939
R12468 gnd.n6624 gnd.n689 0.152939
R12469 gnd.n6634 gnd.n689 0.152939
R12470 gnd.n6635 gnd.n684 0.152939
R12471 gnd.n6643 gnd.n684 0.152939
R12472 gnd.n6644 gnd.n6643 0.152939
R12473 gnd.n6645 gnd.n6644 0.152939
R12474 gnd.n6645 gnd.n678 0.152939
R12475 gnd.n6653 gnd.n678 0.152939
R12476 gnd.n6654 gnd.n6653 0.152939
R12477 gnd.n6655 gnd.n6654 0.152939
R12478 gnd.n6655 gnd.n672 0.152939
R12479 gnd.n6663 gnd.n672 0.152939
R12480 gnd.n6664 gnd.n6663 0.152939
R12481 gnd.n6665 gnd.n6664 0.152939
R12482 gnd.n6665 gnd.n666 0.152939
R12483 gnd.n6673 gnd.n666 0.152939
R12484 gnd.n6674 gnd.n6673 0.152939
R12485 gnd.n6675 gnd.n6674 0.152939
R12486 gnd.n6675 gnd.n660 0.152939
R12487 gnd.n6683 gnd.n660 0.152939
R12488 gnd.n6684 gnd.n6683 0.152939
R12489 gnd.n6685 gnd.n6684 0.152939
R12490 gnd.n6685 gnd.n654 0.152939
R12491 gnd.n6693 gnd.n654 0.152939
R12492 gnd.n6694 gnd.n6693 0.152939
R12493 gnd.n6695 gnd.n6694 0.152939
R12494 gnd.n6695 gnd.n648 0.152939
R12495 gnd.n6703 gnd.n648 0.152939
R12496 gnd.n6704 gnd.n6703 0.152939
R12497 gnd.n6705 gnd.n6704 0.152939
R12498 gnd.n6705 gnd.n642 0.152939
R12499 gnd.n6713 gnd.n642 0.152939
R12500 gnd.n6714 gnd.n6713 0.152939
R12501 gnd.n6715 gnd.n6714 0.152939
R12502 gnd.n6715 gnd.n636 0.152939
R12503 gnd.n6723 gnd.n636 0.152939
R12504 gnd.n6724 gnd.n6723 0.152939
R12505 gnd.n6725 gnd.n6724 0.152939
R12506 gnd.n6725 gnd.n630 0.152939
R12507 gnd.n6733 gnd.n630 0.152939
R12508 gnd.n6734 gnd.n6733 0.152939
R12509 gnd.n6735 gnd.n6734 0.152939
R12510 gnd.n6735 gnd.n624 0.152939
R12511 gnd.n6743 gnd.n624 0.152939
R12512 gnd.n6744 gnd.n6743 0.152939
R12513 gnd.n6745 gnd.n6744 0.152939
R12514 gnd.n6745 gnd.n618 0.152939
R12515 gnd.n6753 gnd.n618 0.152939
R12516 gnd.n6754 gnd.n6753 0.152939
R12517 gnd.n6755 gnd.n6754 0.152939
R12518 gnd.n6755 gnd.n612 0.152939
R12519 gnd.n6763 gnd.n612 0.152939
R12520 gnd.n6764 gnd.n6763 0.152939
R12521 gnd.n6765 gnd.n6764 0.152939
R12522 gnd.n6765 gnd.n606 0.152939
R12523 gnd.n6773 gnd.n606 0.152939
R12524 gnd.n6774 gnd.n6773 0.152939
R12525 gnd.n6775 gnd.n6774 0.152939
R12526 gnd.n6775 gnd.n600 0.152939
R12527 gnd.n6783 gnd.n600 0.152939
R12528 gnd.n6784 gnd.n6783 0.152939
R12529 gnd.n6785 gnd.n6784 0.152939
R12530 gnd.n6785 gnd.n594 0.152939
R12531 gnd.n6793 gnd.n594 0.152939
R12532 gnd.n6794 gnd.n6793 0.152939
R12533 gnd.n6795 gnd.n6794 0.152939
R12534 gnd.n6795 gnd.n588 0.152939
R12535 gnd.n6803 gnd.n588 0.152939
R12536 gnd.n6804 gnd.n6803 0.152939
R12537 gnd.n6805 gnd.n6804 0.152939
R12538 gnd.n6805 gnd.n582 0.152939
R12539 gnd.n6813 gnd.n582 0.152939
R12540 gnd.n6814 gnd.n6813 0.152939
R12541 gnd.n6815 gnd.n6814 0.152939
R12542 gnd.n6815 gnd.n576 0.152939
R12543 gnd.n6823 gnd.n576 0.152939
R12544 gnd.n6824 gnd.n6823 0.152939
R12545 gnd.n6825 gnd.n6824 0.152939
R12546 gnd.n6825 gnd.n570 0.152939
R12547 gnd.n6833 gnd.n570 0.152939
R12548 gnd.n6834 gnd.n6833 0.152939
R12549 gnd.n6835 gnd.n6834 0.152939
R12550 gnd.n6835 gnd.n564 0.152939
R12551 gnd.n6844 gnd.n564 0.152939
R12552 gnd.n6845 gnd.n6844 0.152939
R12553 gnd.n6846 gnd.n6845 0.152939
R12554 gnd.n7020 gnd.n76 0.152939
R12555 gnd.n101 gnd.n76 0.152939
R12556 gnd.n102 gnd.n101 0.152939
R12557 gnd.n103 gnd.n102 0.152939
R12558 gnd.n118 gnd.n103 0.152939
R12559 gnd.n119 gnd.n118 0.152939
R12560 gnd.n120 gnd.n119 0.152939
R12561 gnd.n121 gnd.n120 0.152939
R12562 gnd.n138 gnd.n121 0.152939
R12563 gnd.n139 gnd.n138 0.152939
R12564 gnd.n140 gnd.n139 0.152939
R12565 gnd.n141 gnd.n140 0.152939
R12566 gnd.n157 gnd.n141 0.152939
R12567 gnd.n158 gnd.n157 0.152939
R12568 gnd.n159 gnd.n158 0.152939
R12569 gnd.n160 gnd.n159 0.152939
R12570 gnd.n7029 gnd.n65 0.152939
R12571 gnd.n214 gnd.n65 0.152939
R12572 gnd.n215 gnd.n214 0.152939
R12573 gnd.n219 gnd.n215 0.152939
R12574 gnd.n220 gnd.n219 0.152939
R12575 gnd.n221 gnd.n220 0.152939
R12576 gnd.n221 gnd.n211 0.152939
R12577 gnd.n226 gnd.n211 0.152939
R12578 gnd.n227 gnd.n226 0.152939
R12579 gnd.n228 gnd.n227 0.152939
R12580 gnd.n228 gnd.n208 0.152939
R12581 gnd.n233 gnd.n208 0.152939
R12582 gnd.n234 gnd.n233 0.152939
R12583 gnd.n235 gnd.n234 0.152939
R12584 gnd.n235 gnd.n205 0.152939
R12585 gnd.n240 gnd.n205 0.152939
R12586 gnd.n241 gnd.n240 0.152939
R12587 gnd.n242 gnd.n241 0.152939
R12588 gnd.n242 gnd.n202 0.152939
R12589 gnd.n247 gnd.n202 0.152939
R12590 gnd.n280 gnd.n168 0.152939
R12591 gnd.n170 gnd.n168 0.152939
R12592 gnd.n174 gnd.n170 0.152939
R12593 gnd.n175 gnd.n174 0.152939
R12594 gnd.n176 gnd.n175 0.152939
R12595 gnd.n177 gnd.n176 0.152939
R12596 gnd.n181 gnd.n177 0.152939
R12597 gnd.n182 gnd.n181 0.152939
R12598 gnd.n183 gnd.n182 0.152939
R12599 gnd.n184 gnd.n183 0.152939
R12600 gnd.n188 gnd.n184 0.152939
R12601 gnd.n189 gnd.n188 0.152939
R12602 gnd.n190 gnd.n189 0.152939
R12603 gnd.n191 gnd.n190 0.152939
R12604 gnd.n195 gnd.n191 0.152939
R12605 gnd.n196 gnd.n195 0.152939
R12606 gnd.n249 gnd.n196 0.152939
R12607 gnd.n249 gnd.n248 0.152939
R12608 gnd.n344 gnd.n343 0.152939
R12609 gnd.n352 gnd.n343 0.152939
R12610 gnd.n353 gnd.n352 0.152939
R12611 gnd.n354 gnd.n353 0.152939
R12612 gnd.n354 gnd.n339 0.152939
R12613 gnd.n362 gnd.n339 0.152939
R12614 gnd.n363 gnd.n362 0.152939
R12615 gnd.n364 gnd.n363 0.152939
R12616 gnd.n364 gnd.n335 0.152939
R12617 gnd.n372 gnd.n335 0.152939
R12618 gnd.n373 gnd.n372 0.152939
R12619 gnd.n374 gnd.n373 0.152939
R12620 gnd.n374 gnd.n331 0.152939
R12621 gnd.n383 gnd.n331 0.152939
R12622 gnd.n384 gnd.n383 0.152939
R12623 gnd.n385 gnd.n384 0.152939
R12624 gnd.n385 gnd.n325 0.152939
R12625 gnd.n393 gnd.n325 0.152939
R12626 gnd.n394 gnd.n393 0.152939
R12627 gnd.n395 gnd.n394 0.152939
R12628 gnd.n395 gnd.n321 0.152939
R12629 gnd.n403 gnd.n321 0.152939
R12630 gnd.n404 gnd.n403 0.152939
R12631 gnd.n405 gnd.n404 0.152939
R12632 gnd.n405 gnd.n317 0.152939
R12633 gnd.n413 gnd.n317 0.152939
R12634 gnd.n414 gnd.n413 0.152939
R12635 gnd.n415 gnd.n414 0.152939
R12636 gnd.n415 gnd.n313 0.152939
R12637 gnd.n423 gnd.n313 0.152939
R12638 gnd.n424 gnd.n423 0.152939
R12639 gnd.n425 gnd.n424 0.152939
R12640 gnd.n425 gnd.n309 0.152939
R12641 gnd.n433 gnd.n309 0.152939
R12642 gnd.n434 gnd.n433 0.152939
R12643 gnd.n435 gnd.n434 0.152939
R12644 gnd.n435 gnd.n303 0.152939
R12645 gnd.n443 gnd.n303 0.152939
R12646 gnd.n444 gnd.n443 0.152939
R12647 gnd.n445 gnd.n444 0.152939
R12648 gnd.n445 gnd.n299 0.152939
R12649 gnd.n453 gnd.n299 0.152939
R12650 gnd.n454 gnd.n453 0.152939
R12651 gnd.n455 gnd.n454 0.152939
R12652 gnd.n455 gnd.n295 0.152939
R12653 gnd.n463 gnd.n295 0.152939
R12654 gnd.n464 gnd.n463 0.152939
R12655 gnd.n465 gnd.n464 0.152939
R12656 gnd.n465 gnd.n291 0.152939
R12657 gnd.n473 gnd.n291 0.152939
R12658 gnd.n474 gnd.n473 0.152939
R12659 gnd.n475 gnd.n474 0.152939
R12660 gnd.n475 gnd.n287 0.152939
R12661 gnd.n483 gnd.n287 0.152939
R12662 gnd.n484 gnd.n483 0.152939
R12663 gnd.n485 gnd.n484 0.152939
R12664 gnd.n485 gnd.n281 0.152939
R12665 gnd.n492 gnd.n281 0.152939
R12666 gnd.n1604 gnd.n1603 0.152939
R12667 gnd.n1605 gnd.n1604 0.152939
R12668 gnd.n1606 gnd.n1605 0.152939
R12669 gnd.n1607 gnd.n1606 0.152939
R12670 gnd.n1608 gnd.n1607 0.152939
R12671 gnd.n1609 gnd.n1608 0.152939
R12672 gnd.n1610 gnd.n1609 0.152939
R12673 gnd.n1611 gnd.n1610 0.152939
R12674 gnd.n1612 gnd.n1611 0.152939
R12675 gnd.n1613 gnd.n1612 0.152939
R12676 gnd.n1614 gnd.n1613 0.152939
R12677 gnd.n1615 gnd.n1614 0.152939
R12678 gnd.n1616 gnd.n1615 0.152939
R12679 gnd.n1617 gnd.n1616 0.152939
R12680 gnd.n1618 gnd.n1617 0.152939
R12681 gnd.n1619 gnd.n1618 0.152939
R12682 gnd.n1620 gnd.n1619 0.152939
R12683 gnd.n1623 gnd.n1620 0.152939
R12684 gnd.n1624 gnd.n1623 0.152939
R12685 gnd.n1625 gnd.n1624 0.152939
R12686 gnd.n1626 gnd.n1625 0.152939
R12687 gnd.n1627 gnd.n1626 0.152939
R12688 gnd.n1628 gnd.n1627 0.152939
R12689 gnd.n1629 gnd.n1628 0.152939
R12690 gnd.n1630 gnd.n1629 0.152939
R12691 gnd.n1635 gnd.n1634 0.152939
R12692 gnd.n1636 gnd.n1635 0.152939
R12693 gnd.n1637 gnd.n1636 0.152939
R12694 gnd.n1638 gnd.n1637 0.152939
R12695 gnd.n1639 gnd.n1638 0.152939
R12696 gnd.n1640 gnd.n1639 0.152939
R12697 gnd.n1641 gnd.n1640 0.152939
R12698 gnd.n1642 gnd.n1641 0.152939
R12699 gnd.n1643 gnd.n1642 0.152939
R12700 gnd.n1646 gnd.n1643 0.152939
R12701 gnd.n1647 gnd.n1646 0.152939
R12702 gnd.n1648 gnd.n1647 0.152939
R12703 gnd.n1649 gnd.n1648 0.152939
R12704 gnd.n1650 gnd.n1649 0.152939
R12705 gnd.n1651 gnd.n1650 0.152939
R12706 gnd.n1652 gnd.n1651 0.152939
R12707 gnd.n1653 gnd.n1652 0.152939
R12708 gnd.n1654 gnd.n1653 0.152939
R12709 gnd.n1655 gnd.n1654 0.152939
R12710 gnd.n1656 gnd.n1655 0.152939
R12711 gnd.n1657 gnd.n1656 0.152939
R12712 gnd.n1658 gnd.n1657 0.152939
R12713 gnd.n1659 gnd.n1658 0.152939
R12714 gnd.n1660 gnd.n1659 0.152939
R12715 gnd.n1661 gnd.n1660 0.152939
R12716 gnd.n1662 gnd.n1661 0.152939
R12717 gnd.n1663 gnd.n1662 0.152939
R12718 gnd.n1664 gnd.n1663 0.152939
R12719 gnd.n5641 gnd.n1664 0.152939
R12720 gnd.n5641 gnd.n5640 0.152939
R12721 gnd.n1685 gnd.n1684 0.152939
R12722 gnd.n1686 gnd.n1685 0.152939
R12723 gnd.n1687 gnd.n1686 0.152939
R12724 gnd.n1688 gnd.n1687 0.152939
R12725 gnd.n1709 gnd.n1688 0.152939
R12726 gnd.n1710 gnd.n1709 0.152939
R12727 gnd.n1711 gnd.n1710 0.152939
R12728 gnd.n1712 gnd.n1711 0.152939
R12729 gnd.n1713 gnd.n1712 0.152939
R12730 gnd.n1713 gnd.n543 0.152939
R12731 gnd.n6867 gnd.n543 0.152939
R12732 gnd.n6868 gnd.n6867 0.152939
R12733 gnd.n6869 gnd.n6868 0.152939
R12734 gnd.n6870 gnd.n6869 0.152939
R12735 gnd.n6870 gnd.n77 0.152939
R12736 gnd.n7020 gnd.n77 0.152939
R12737 gnd.n6851 gnd.n561 0.152939
R12738 gnd.n4404 gnd.n4400 0.152939
R12739 gnd.n4405 gnd.n4404 0.152939
R12740 gnd.n4406 gnd.n4405 0.152939
R12741 gnd.n4406 gnd.n2322 0.152939
R12742 gnd.n4412 gnd.n2322 0.152939
R12743 gnd.n4413 gnd.n4412 0.152939
R12744 gnd.n4414 gnd.n4413 0.152939
R12745 gnd.n4415 gnd.n4414 0.152939
R12746 gnd.n4416 gnd.n4415 0.152939
R12747 gnd.n4416 gnd.n2304 0.152939
R12748 gnd.n4695 gnd.n2304 0.152939
R12749 gnd.n4696 gnd.n4695 0.152939
R12750 gnd.n4697 gnd.n4696 0.152939
R12751 gnd.n4697 gnd.n2300 0.152939
R12752 gnd.n4703 gnd.n2300 0.152939
R12753 gnd.n4704 gnd.n4703 0.152939
R12754 gnd.n4705 gnd.n4704 0.152939
R12755 gnd.n4706 gnd.n4705 0.152939
R12756 gnd.n4707 gnd.n4706 0.152939
R12757 gnd.n4707 gnd.n2270 0.152939
R12758 gnd.n4741 gnd.n2270 0.152939
R12759 gnd.n4742 gnd.n4741 0.152939
R12760 gnd.n4743 gnd.n4742 0.152939
R12761 gnd.n4744 gnd.n4743 0.152939
R12762 gnd.n4745 gnd.n4744 0.152939
R12763 gnd.n4747 gnd.n4745 0.152939
R12764 gnd.n4747 gnd.n4746 0.152939
R12765 gnd.n4746 gnd.n1285 0.152939
R12766 gnd.n1286 gnd.n1285 0.152939
R12767 gnd.n1287 gnd.n1286 0.152939
R12768 gnd.n1385 gnd.n1287 0.152939
R12769 gnd.n1386 gnd.n1385 0.152939
R12770 gnd.n1387 gnd.n1386 0.152939
R12771 gnd.n1388 gnd.n1387 0.152939
R12772 gnd.n1389 gnd.n1388 0.152939
R12773 gnd.n4840 gnd.n1389 0.152939
R12774 gnd.n4841 gnd.n4840 0.152939
R12775 gnd.n4842 gnd.n4841 0.152939
R12776 gnd.n4842 gnd.n2226 0.152939
R12777 gnd.n4882 gnd.n2226 0.152939
R12778 gnd.n4883 gnd.n4882 0.152939
R12779 gnd.n4885 gnd.n4883 0.152939
R12780 gnd.n4885 gnd.n4884 0.152939
R12781 gnd.n4884 gnd.n2196 0.152939
R12782 gnd.n2197 gnd.n2196 0.152939
R12783 gnd.n2198 gnd.n2197 0.152939
R12784 gnd.n2201 gnd.n2198 0.152939
R12785 gnd.n2202 gnd.n2201 0.152939
R12786 gnd.n2203 gnd.n2202 0.152939
R12787 gnd.n2204 gnd.n2203 0.152939
R12788 gnd.n2205 gnd.n2204 0.152939
R12789 gnd.n2205 gnd.n2153 0.152939
R12790 gnd.n4997 gnd.n2153 0.152939
R12791 gnd.n4998 gnd.n4997 0.152939
R12792 gnd.n4999 gnd.n4998 0.152939
R12793 gnd.n5000 gnd.n4999 0.152939
R12794 gnd.n5000 gnd.n2127 0.152939
R12795 gnd.n5053 gnd.n2127 0.152939
R12796 gnd.n5054 gnd.n5053 0.152939
R12797 gnd.n5055 gnd.n5054 0.152939
R12798 gnd.n5056 gnd.n5055 0.152939
R12799 gnd.n5056 gnd.n2105 0.152939
R12800 gnd.n5100 gnd.n2105 0.152939
R12801 gnd.n5101 gnd.n5100 0.152939
R12802 gnd.n5102 gnd.n5101 0.152939
R12803 gnd.n5102 gnd.n2081 0.152939
R12804 gnd.n5130 gnd.n2081 0.152939
R12805 gnd.n5131 gnd.n5130 0.152939
R12806 gnd.n5132 gnd.n5131 0.152939
R12807 gnd.n5132 gnd.n2063 0.152939
R12808 gnd.n5178 gnd.n2063 0.152939
R12809 gnd.n5179 gnd.n5178 0.152939
R12810 gnd.n5180 gnd.n5179 0.152939
R12811 gnd.n5181 gnd.n5180 0.152939
R12812 gnd.n5181 gnd.n2037 0.152939
R12813 gnd.n5214 gnd.n2037 0.152939
R12814 gnd.n5215 gnd.n5214 0.152939
R12815 gnd.n5216 gnd.n5215 0.152939
R12816 gnd.n5217 gnd.n5216 0.152939
R12817 gnd.n5217 gnd.n2007 0.152939
R12818 gnd.n5278 gnd.n2007 0.152939
R12819 gnd.n5279 gnd.n5278 0.152939
R12820 gnd.n5280 gnd.n5279 0.152939
R12821 gnd.n5280 gnd.n1990 0.152939
R12822 gnd.n5307 gnd.n1990 0.152939
R12823 gnd.n5308 gnd.n5307 0.152939
R12824 gnd.n5309 gnd.n5308 0.152939
R12825 gnd.n5310 gnd.n5309 0.152939
R12826 gnd.n5310 gnd.n1964 0.152939
R12827 gnd.n5343 gnd.n1964 0.152939
R12828 gnd.n5344 gnd.n5343 0.152939
R12829 gnd.n5345 gnd.n5344 0.152939
R12830 gnd.n5345 gnd.n1936 0.152939
R12831 gnd.n5380 gnd.n1936 0.152939
R12832 gnd.n5381 gnd.n5380 0.152939
R12833 gnd.n5382 gnd.n5381 0.152939
R12834 gnd.n5383 gnd.n5382 0.152939
R12835 gnd.n5383 gnd.n1787 0.152939
R12836 gnd.n5488 gnd.n1787 0.152939
R12837 gnd.n5489 gnd.n5488 0.152939
R12838 gnd.n5490 gnd.n5489 0.152939
R12839 gnd.n5492 gnd.n5490 0.152939
R12840 gnd.n5492 gnd.n5491 0.152939
R12841 gnd.n5491 gnd.n1776 0.152939
R12842 gnd.n5509 gnd.n1776 0.152939
R12843 gnd.n5510 gnd.n5509 0.152939
R12844 gnd.n5511 gnd.n5510 0.152939
R12845 gnd.n5512 gnd.n5511 0.152939
R12846 gnd.n5513 gnd.n5512 0.152939
R12847 gnd.n5515 gnd.n5513 0.152939
R12848 gnd.n5516 gnd.n5515 0.152939
R12849 gnd.n5518 gnd.n5516 0.152939
R12850 gnd.n5518 gnd.n5517 0.152939
R12851 gnd.n5517 gnd.n1740 0.152939
R12852 gnd.n5578 gnd.n1740 0.152939
R12853 gnd.n5579 gnd.n5578 0.152939
R12854 gnd.n5580 gnd.n5579 0.152939
R12855 gnd.n5580 gnd.n1736 0.152939
R12856 gnd.n5586 gnd.n1736 0.152939
R12857 gnd.n5587 gnd.n5586 0.152939
R12858 gnd.n5588 gnd.n5587 0.152939
R12859 gnd.n5589 gnd.n5588 0.152939
R12860 gnd.n5590 gnd.n5589 0.152939
R12861 gnd.n5592 gnd.n5590 0.152939
R12862 gnd.n5592 gnd.n5591 0.152939
R12863 gnd.n5591 gnd.n560 0.152939
R12864 gnd.n561 gnd.n560 0.152939
R12865 gnd.n4083 gnd.n4027 0.152939
R12866 gnd.n4028 gnd.n4027 0.152939
R12867 gnd.n4029 gnd.n4028 0.152939
R12868 gnd.n4030 gnd.n4029 0.152939
R12869 gnd.n4031 gnd.n4030 0.152939
R12870 gnd.n4032 gnd.n4031 0.152939
R12871 gnd.n4033 gnd.n4032 0.152939
R12872 gnd.n4034 gnd.n4033 0.152939
R12873 gnd.n4035 gnd.n4034 0.152939
R12874 gnd.n4036 gnd.n4035 0.152939
R12875 gnd.n4037 gnd.n4036 0.152939
R12876 gnd.n4038 gnd.n4037 0.152939
R12877 gnd.n4039 gnd.n4038 0.152939
R12878 gnd.n4040 gnd.n4039 0.152939
R12879 gnd.n4041 gnd.n4040 0.152939
R12880 gnd.n4042 gnd.n4041 0.152939
R12881 gnd.n4043 gnd.n4042 0.152939
R12882 gnd.n4044 gnd.n4043 0.152939
R12883 gnd.n4045 gnd.n4044 0.152939
R12884 gnd.n4046 gnd.n4045 0.152939
R12885 gnd.n4122 gnd.n4008 0.152939
R12886 gnd.n4009 gnd.n4008 0.152939
R12887 gnd.n4010 gnd.n4009 0.152939
R12888 gnd.n4011 gnd.n4010 0.152939
R12889 gnd.n4012 gnd.n4011 0.152939
R12890 gnd.n4013 gnd.n4012 0.152939
R12891 gnd.n4014 gnd.n4013 0.152939
R12892 gnd.n4015 gnd.n4014 0.152939
R12893 gnd.n4016 gnd.n4015 0.152939
R12894 gnd.n4017 gnd.n4016 0.152939
R12895 gnd.n4018 gnd.n4017 0.152939
R12896 gnd.n4019 gnd.n4018 0.152939
R12897 gnd.n4020 gnd.n4019 0.152939
R12898 gnd.n4021 gnd.n4020 0.152939
R12899 gnd.n4022 gnd.n4021 0.152939
R12900 gnd.n4087 gnd.n4022 0.152939
R12901 gnd.n4087 gnd.n4086 0.152939
R12902 gnd.n4086 gnd.n4085 0.152939
R12903 gnd.n1059 gnd.n1058 0.152939
R12904 gnd.n1078 gnd.n1059 0.152939
R12905 gnd.n1079 gnd.n1078 0.152939
R12906 gnd.n1080 gnd.n1079 0.152939
R12907 gnd.n1081 gnd.n1080 0.152939
R12908 gnd.n1098 gnd.n1081 0.152939
R12909 gnd.n1099 gnd.n1098 0.152939
R12910 gnd.n1100 gnd.n1099 0.152939
R12911 gnd.n1101 gnd.n1100 0.152939
R12912 gnd.n1118 gnd.n1101 0.152939
R12913 gnd.n1119 gnd.n1118 0.152939
R12914 gnd.n1120 gnd.n1119 0.152939
R12915 gnd.n1121 gnd.n1120 0.152939
R12916 gnd.n1139 gnd.n1121 0.152939
R12917 gnd.n1140 gnd.n1139 0.152939
R12918 gnd.n6088 gnd.n1140 0.152939
R12919 gnd.n6087 gnd.n1141 0.152939
R12920 gnd.n1185 gnd.n1141 0.152939
R12921 gnd.n1186 gnd.n1185 0.152939
R12922 gnd.n1187 gnd.n1186 0.152939
R12923 gnd.n1188 gnd.n1187 0.152939
R12924 gnd.n1189 gnd.n1188 0.152939
R12925 gnd.n1190 gnd.n1189 0.152939
R12926 gnd.n1191 gnd.n1190 0.152939
R12927 gnd.n1192 gnd.n1191 0.152939
R12928 gnd.n1193 gnd.n1192 0.152939
R12929 gnd.n1194 gnd.n1193 0.152939
R12930 gnd.n1195 gnd.n1194 0.152939
R12931 gnd.n1196 gnd.n1195 0.152939
R12932 gnd.n1197 gnd.n1196 0.152939
R12933 gnd.n1198 gnd.n1197 0.152939
R12934 gnd.n1199 gnd.n1198 0.152939
R12935 gnd.n1200 gnd.n1199 0.152939
R12936 gnd.n1203 gnd.n1200 0.152939
R12937 gnd.n1204 gnd.n1203 0.152939
R12938 gnd.n1205 gnd.n1204 0.152939
R12939 gnd.n1206 gnd.n1205 0.152939
R12940 gnd.n1207 gnd.n1206 0.152939
R12941 gnd.n1208 gnd.n1207 0.152939
R12942 gnd.n1209 gnd.n1208 0.152939
R12943 gnd.n1210 gnd.n1209 0.152939
R12944 gnd.n4596 gnd.n4595 0.152939
R12945 gnd.n4603 gnd.n4596 0.152939
R12946 gnd.n4604 gnd.n4603 0.152939
R12947 gnd.n4605 gnd.n4604 0.152939
R12948 gnd.n4605 gnd.n4593 0.152939
R12949 gnd.n4613 gnd.n4593 0.152939
R12950 gnd.n4614 gnd.n4613 0.152939
R12951 gnd.n4615 gnd.n4614 0.152939
R12952 gnd.n4615 gnd.n4588 0.152939
R12953 gnd.n4622 gnd.n4588 0.152939
R12954 gnd.n4623 gnd.n4622 0.152939
R12955 gnd.n4624 gnd.n4623 0.152939
R12956 gnd.n4624 gnd.n4586 0.152939
R12957 gnd.n4632 gnd.n4586 0.152939
R12958 gnd.n4633 gnd.n4632 0.152939
R12959 gnd.n4634 gnd.n4633 0.152939
R12960 gnd.n4634 gnd.n4584 0.152939
R12961 gnd.n4642 gnd.n4584 0.152939
R12962 gnd.n4643 gnd.n4642 0.152939
R12963 gnd.n4644 gnd.n4643 0.152939
R12964 gnd.n4644 gnd.n4582 0.152939
R12965 gnd.n4652 gnd.n4582 0.152939
R12966 gnd.n4653 gnd.n4652 0.152939
R12967 gnd.n4654 gnd.n4653 0.152939
R12968 gnd.n4654 gnd.n4580 0.152939
R12969 gnd.n4662 gnd.n4580 0.152939
R12970 gnd.n4663 gnd.n4662 0.152939
R12971 gnd.n4664 gnd.n4663 0.152939
R12972 gnd.n4664 gnd.n4575 0.152939
R12973 gnd.n4670 gnd.n4575 0.152939
R12974 gnd.n3946 gnd.n3945 0.152939
R12975 gnd.n3947 gnd.n3946 0.152939
R12976 gnd.n3948 gnd.n3947 0.152939
R12977 gnd.n3949 gnd.n3948 0.152939
R12978 gnd.n3950 gnd.n3949 0.152939
R12979 gnd.n3951 gnd.n3950 0.152939
R12980 gnd.n3952 gnd.n3951 0.152939
R12981 gnd.n3953 gnd.n3952 0.152939
R12982 gnd.n3954 gnd.n3953 0.152939
R12983 gnd.n3955 gnd.n3954 0.152939
R12984 gnd.n3956 gnd.n3955 0.152939
R12985 gnd.n3957 gnd.n3956 0.152939
R12986 gnd.n3958 gnd.n3957 0.152939
R12987 gnd.n3959 gnd.n3958 0.152939
R12988 gnd.n3960 gnd.n3959 0.152939
R12989 gnd.n3961 gnd.n3960 0.152939
R12990 gnd.n3962 gnd.n3961 0.152939
R12991 gnd.n3965 gnd.n3962 0.152939
R12992 gnd.n3966 gnd.n3965 0.152939
R12993 gnd.n3967 gnd.n3966 0.152939
R12994 gnd.n3968 gnd.n3967 0.152939
R12995 gnd.n3969 gnd.n3968 0.152939
R12996 gnd.n3970 gnd.n3969 0.152939
R12997 gnd.n3971 gnd.n3970 0.152939
R12998 gnd.n3972 gnd.n3971 0.152939
R12999 gnd.n3973 gnd.n3972 0.152939
R13000 gnd.n3974 gnd.n3973 0.152939
R13001 gnd.n3975 gnd.n3974 0.152939
R13002 gnd.n3976 gnd.n3975 0.152939
R13003 gnd.n3977 gnd.n3976 0.152939
R13004 gnd.n3978 gnd.n3977 0.152939
R13005 gnd.n3979 gnd.n3978 0.152939
R13006 gnd.n3980 gnd.n3979 0.152939
R13007 gnd.n3981 gnd.n3980 0.152939
R13008 gnd.n3982 gnd.n3981 0.152939
R13009 gnd.n3983 gnd.n3982 0.152939
R13010 gnd.n3984 gnd.n3983 0.152939
R13011 gnd.n3987 gnd.n3984 0.152939
R13012 gnd.n3988 gnd.n3987 0.152939
R13013 gnd.n3989 gnd.n3988 0.152939
R13014 gnd.n3990 gnd.n3989 0.152939
R13015 gnd.n3991 gnd.n3990 0.152939
R13016 gnd.n3992 gnd.n3991 0.152939
R13017 gnd.n3993 gnd.n3992 0.152939
R13018 gnd.n3994 gnd.n3993 0.152939
R13019 gnd.n3995 gnd.n3994 0.152939
R13020 gnd.n3996 gnd.n3995 0.152939
R13021 gnd.n3997 gnd.n3996 0.152939
R13022 gnd.n3998 gnd.n3997 0.152939
R13023 gnd.n3999 gnd.n3998 0.152939
R13024 gnd.n4000 gnd.n3999 0.152939
R13025 gnd.n4001 gnd.n4000 0.152939
R13026 gnd.n4002 gnd.n4001 0.152939
R13027 gnd.n4003 gnd.n4002 0.152939
R13028 gnd.n4004 gnd.n4003 0.152939
R13029 gnd.n4005 gnd.n4004 0.152939
R13030 gnd.n4125 gnd.n4005 0.152939
R13031 gnd.n4125 gnd.n4124 0.152939
R13032 gnd.n4254 gnd.n2427 0.152939
R13033 gnd.n4255 gnd.n4254 0.152939
R13034 gnd.n4256 gnd.n4255 0.152939
R13035 gnd.n4256 gnd.n2408 0.152939
R13036 gnd.n4274 gnd.n2408 0.152939
R13037 gnd.n4275 gnd.n4274 0.152939
R13038 gnd.n4276 gnd.n4275 0.152939
R13039 gnd.n4276 gnd.n2391 0.152939
R13040 gnd.n4294 gnd.n2391 0.152939
R13041 gnd.n4295 gnd.n4294 0.152939
R13042 gnd.n4296 gnd.n4295 0.152939
R13043 gnd.n4296 gnd.n2372 0.152939
R13044 gnd.n4314 gnd.n2372 0.152939
R13045 gnd.n4315 gnd.n4314 0.152939
R13046 gnd.n4316 gnd.n4315 0.152939
R13047 gnd.n4316 gnd.n1058 0.152939
R13048 gnd.n6312 gnd.n881 0.152939
R13049 gnd.n886 gnd.n881 0.152939
R13050 gnd.n887 gnd.n886 0.152939
R13051 gnd.n888 gnd.n887 0.152939
R13052 gnd.n893 gnd.n888 0.152939
R13053 gnd.n894 gnd.n893 0.152939
R13054 gnd.n895 gnd.n894 0.152939
R13055 gnd.n896 gnd.n895 0.152939
R13056 gnd.n901 gnd.n896 0.152939
R13057 gnd.n902 gnd.n901 0.152939
R13058 gnd.n903 gnd.n902 0.152939
R13059 gnd.n904 gnd.n903 0.152939
R13060 gnd.n909 gnd.n904 0.152939
R13061 gnd.n910 gnd.n909 0.152939
R13062 gnd.n911 gnd.n910 0.152939
R13063 gnd.n912 gnd.n911 0.152939
R13064 gnd.n917 gnd.n912 0.152939
R13065 gnd.n918 gnd.n917 0.152939
R13066 gnd.n919 gnd.n918 0.152939
R13067 gnd.n920 gnd.n919 0.152939
R13068 gnd.n925 gnd.n920 0.152939
R13069 gnd.n926 gnd.n925 0.152939
R13070 gnd.n927 gnd.n926 0.152939
R13071 gnd.n928 gnd.n927 0.152939
R13072 gnd.n933 gnd.n928 0.152939
R13073 gnd.n934 gnd.n933 0.152939
R13074 gnd.n935 gnd.n934 0.152939
R13075 gnd.n936 gnd.n935 0.152939
R13076 gnd.n941 gnd.n936 0.152939
R13077 gnd.n942 gnd.n941 0.152939
R13078 gnd.n943 gnd.n942 0.152939
R13079 gnd.n944 gnd.n943 0.152939
R13080 gnd.n949 gnd.n944 0.152939
R13081 gnd.n950 gnd.n949 0.152939
R13082 gnd.n951 gnd.n950 0.152939
R13083 gnd.n952 gnd.n951 0.152939
R13084 gnd.n957 gnd.n952 0.152939
R13085 gnd.n958 gnd.n957 0.152939
R13086 gnd.n959 gnd.n958 0.152939
R13087 gnd.n960 gnd.n959 0.152939
R13088 gnd.n965 gnd.n960 0.152939
R13089 gnd.n966 gnd.n965 0.152939
R13090 gnd.n967 gnd.n966 0.152939
R13091 gnd.n968 gnd.n967 0.152939
R13092 gnd.n973 gnd.n968 0.152939
R13093 gnd.n974 gnd.n973 0.152939
R13094 gnd.n975 gnd.n974 0.152939
R13095 gnd.n976 gnd.n975 0.152939
R13096 gnd.n981 gnd.n976 0.152939
R13097 gnd.n982 gnd.n981 0.152939
R13098 gnd.n983 gnd.n982 0.152939
R13099 gnd.n984 gnd.n983 0.152939
R13100 gnd.n989 gnd.n984 0.152939
R13101 gnd.n990 gnd.n989 0.152939
R13102 gnd.n991 gnd.n990 0.152939
R13103 gnd.n992 gnd.n991 0.152939
R13104 gnd.n997 gnd.n992 0.152939
R13105 gnd.n998 gnd.n997 0.152939
R13106 gnd.n999 gnd.n998 0.152939
R13107 gnd.n1000 gnd.n999 0.152939
R13108 gnd.n1005 gnd.n1000 0.152939
R13109 gnd.n1006 gnd.n1005 0.152939
R13110 gnd.n1007 gnd.n1006 0.152939
R13111 gnd.n1008 gnd.n1007 0.152939
R13112 gnd.n1013 gnd.n1008 0.152939
R13113 gnd.n1014 gnd.n1013 0.152939
R13114 gnd.n1015 gnd.n1014 0.152939
R13115 gnd.n1016 gnd.n1015 0.152939
R13116 gnd.n1021 gnd.n1016 0.152939
R13117 gnd.n1022 gnd.n1021 0.152939
R13118 gnd.n1023 gnd.n1022 0.152939
R13119 gnd.n1024 gnd.n1023 0.152939
R13120 gnd.n1029 gnd.n1024 0.152939
R13121 gnd.n1030 gnd.n1029 0.152939
R13122 gnd.n1031 gnd.n1030 0.152939
R13123 gnd.n1032 gnd.n1031 0.152939
R13124 gnd.n1037 gnd.n1032 0.152939
R13125 gnd.n1038 gnd.n1037 0.152939
R13126 gnd.n1039 gnd.n1038 0.152939
R13127 gnd.n1040 gnd.n1039 0.152939
R13128 gnd.n1045 gnd.n1040 0.152939
R13129 gnd.n1046 gnd.n1045 0.152939
R13130 gnd.n1047 gnd.n1046 0.152939
R13131 gnd.n1048 gnd.n1047 0.152939
R13132 gnd.n4734 gnd.n4721 0.152939
R13133 gnd.n4730 gnd.n4721 0.152939
R13134 gnd.n4730 gnd.n4729 0.152939
R13135 gnd.n4729 gnd.n4728 0.152939
R13136 gnd.n4728 gnd.n2255 0.152939
R13137 gnd.n4780 gnd.n2255 0.152939
R13138 gnd.n4781 gnd.n4780 0.152939
R13139 gnd.n4785 gnd.n4781 0.152939
R13140 gnd.n4785 gnd.n4784 0.152939
R13141 gnd.n4784 gnd.n4783 0.152939
R13142 gnd.n4783 gnd.n1399 0.152939
R13143 gnd.n5930 gnd.n1399 0.152939
R13144 gnd.n5930 gnd.n5929 0.152939
R13145 gnd.n5929 gnd.n5928 0.152939
R13146 gnd.n5928 gnd.n1400 0.152939
R13147 gnd.n5924 gnd.n1400 0.152939
R13148 gnd.n5924 gnd.n5923 0.152939
R13149 gnd.n5923 gnd.n5922 0.152939
R13150 gnd.n5922 gnd.n1405 0.152939
R13151 gnd.n5918 gnd.n1405 0.152939
R13152 gnd.n5918 gnd.n5917 0.152939
R13153 gnd.n5917 gnd.n5916 0.152939
R13154 gnd.n5916 gnd.n1410 0.152939
R13155 gnd.n5912 gnd.n1410 0.152939
R13156 gnd.n5912 gnd.n5911 0.152939
R13157 gnd.n5911 gnd.n5910 0.152939
R13158 gnd.n5910 gnd.n1415 0.152939
R13159 gnd.n5906 gnd.n1415 0.152939
R13160 gnd.n5906 gnd.n5905 0.152939
R13161 gnd.n5905 gnd.n5904 0.152939
R13162 gnd.n5904 gnd.n1420 0.152939
R13163 gnd.n5900 gnd.n1420 0.152939
R13164 gnd.n5900 gnd.n5899 0.152939
R13165 gnd.n5899 gnd.n5898 0.152939
R13166 gnd.n5898 gnd.n1425 0.152939
R13167 gnd.n5894 gnd.n1425 0.152939
R13168 gnd.n5894 gnd.n5893 0.152939
R13169 gnd.n5893 gnd.n5892 0.152939
R13170 gnd.n5892 gnd.n1430 0.152939
R13171 gnd.n5888 gnd.n1430 0.152939
R13172 gnd.n5888 gnd.n5887 0.152939
R13173 gnd.n5887 gnd.n5886 0.152939
R13174 gnd.n5886 gnd.n1435 0.152939
R13175 gnd.n5882 gnd.n1435 0.152939
R13176 gnd.n5882 gnd.n5881 0.152939
R13177 gnd.n5881 gnd.n5880 0.152939
R13178 gnd.n5880 gnd.n1440 0.152939
R13179 gnd.n5876 gnd.n1440 0.152939
R13180 gnd.n5876 gnd.n5875 0.152939
R13181 gnd.n5875 gnd.n5874 0.152939
R13182 gnd.n5874 gnd.n1445 0.152939
R13183 gnd.n5870 gnd.n1445 0.152939
R13184 gnd.n5870 gnd.n5869 0.152939
R13185 gnd.n5869 gnd.n5868 0.152939
R13186 gnd.n5868 gnd.n1450 0.152939
R13187 gnd.n5864 gnd.n1450 0.152939
R13188 gnd.n5864 gnd.n5863 0.152939
R13189 gnd.n5863 gnd.n5862 0.152939
R13190 gnd.n5862 gnd.n1455 0.152939
R13191 gnd.n5858 gnd.n1455 0.152939
R13192 gnd.n5858 gnd.n5857 0.152939
R13193 gnd.n5857 gnd.n5856 0.152939
R13194 gnd.n5856 gnd.n1460 0.152939
R13195 gnd.n5852 gnd.n1460 0.152939
R13196 gnd.n5852 gnd.n5851 0.152939
R13197 gnd.n5851 gnd.n5850 0.152939
R13198 gnd.n5850 gnd.n1465 0.152939
R13199 gnd.n5846 gnd.n1465 0.152939
R13200 gnd.n5846 gnd.n5845 0.152939
R13201 gnd.n5845 gnd.n5844 0.152939
R13202 gnd.n5844 gnd.n1470 0.152939
R13203 gnd.n5840 gnd.n1470 0.152939
R13204 gnd.n5840 gnd.n5839 0.152939
R13205 gnd.n5839 gnd.n5838 0.152939
R13206 gnd.n5838 gnd.n1475 0.152939
R13207 gnd.n5834 gnd.n1475 0.152939
R13208 gnd.n5834 gnd.n5833 0.152939
R13209 gnd.n5833 gnd.n5832 0.152939
R13210 gnd.n5832 gnd.n1480 0.152939
R13211 gnd.n5828 gnd.n1480 0.152939
R13212 gnd.n5828 gnd.n5827 0.152939
R13213 gnd.n5827 gnd.n5826 0.152939
R13214 gnd.n4048 gnd.n2331 0.152939
R13215 gnd.n4371 gnd.n2331 0.152939
R13216 gnd.n4372 gnd.n4371 0.152939
R13217 gnd.n4373 gnd.n4372 0.152939
R13218 gnd.n4373 gnd.n2327 0.152939
R13219 gnd.n4392 gnd.n2327 0.152939
R13220 gnd.n4392 gnd.n4391 0.152939
R13221 gnd.n4391 gnd.n4390 0.152939
R13222 gnd.n4390 gnd.n2316 0.152939
R13223 gnd.n4425 gnd.n2316 0.152939
R13224 gnd.n4426 gnd.n4425 0.152939
R13225 gnd.n4427 gnd.n4426 0.152939
R13226 gnd.n4427 gnd.n2310 0.152939
R13227 gnd.n4687 gnd.n2310 0.152939
R13228 gnd.n4687 gnd.n4686 0.152939
R13229 gnd.n4686 gnd.n4685 0.152939
R13230 gnd.n4685 gnd.n2311 0.152939
R13231 gnd.n4681 gnd.n2311 0.152939
R13232 gnd.n4681 gnd.n4680 0.152939
R13233 gnd.n4680 gnd.n2290 0.152939
R13234 gnd.n4446 gnd.n2262 0.152939
R13235 gnd.n4452 gnd.n4446 0.152939
R13236 gnd.n4453 gnd.n4452 0.152939
R13237 gnd.n4454 gnd.n4453 0.152939
R13238 gnd.n4454 gnd.n4442 0.152939
R13239 gnd.n4573 gnd.n4442 0.152939
R13240 gnd.n4759 gnd.n4758 0.152939
R13241 gnd.n4760 gnd.n4759 0.152939
R13242 gnd.n4760 gnd.n2258 0.152939
R13243 gnd.n4766 gnd.n2258 0.152939
R13244 gnd.n4767 gnd.n4766 0.152939
R13245 gnd.n4768 gnd.n4767 0.152939
R13246 gnd.n4768 gnd.n2249 0.152939
R13247 gnd.n4791 gnd.n2249 0.152939
R13248 gnd.n4792 gnd.n4791 0.152939
R13249 gnd.n4793 gnd.n4792 0.152939
R13250 gnd.n4793 gnd.n2247 0.152939
R13251 gnd.n4827 gnd.n2247 0.152939
R13252 gnd.n4828 gnd.n4827 0.152939
R13253 gnd.n4834 gnd.n4828 0.152939
R13254 gnd.n4834 gnd.n4833 0.152939
R13255 gnd.n4833 gnd.n4832 0.152939
R13256 gnd.n4832 gnd.n4829 0.152939
R13257 gnd.n4829 gnd.n2218 0.152939
R13258 gnd.n4890 gnd.n2218 0.152939
R13259 gnd.n4891 gnd.n4890 0.152939
R13260 gnd.n4892 gnd.n4891 0.152939
R13261 gnd.n4892 gnd.n2216 0.152939
R13262 gnd.n4898 gnd.n2216 0.152939
R13263 gnd.n4899 gnd.n4898 0.152939
R13264 gnd.n4927 gnd.n4899 0.152939
R13265 gnd.n4927 gnd.n4926 0.152939
R13266 gnd.n4926 gnd.n4925 0.152939
R13267 gnd.n4925 gnd.n4900 0.152939
R13268 gnd.n4921 gnd.n4900 0.152939
R13269 gnd.n4921 gnd.n4920 0.152939
R13270 gnd.n4920 gnd.n4919 0.152939
R13271 gnd.n4919 gnd.n4904 0.152939
R13272 gnd.n4915 gnd.n4904 0.152939
R13273 gnd.n4915 gnd.n4914 0.152939
R13274 gnd.n4914 gnd.n4913 0.152939
R13275 gnd.n4913 gnd.n2118 0.152939
R13276 gnd.n5063 gnd.n2118 0.152939
R13277 gnd.n5064 gnd.n5063 0.152939
R13278 gnd.n5086 gnd.n5064 0.152939
R13279 gnd.n5086 gnd.n5085 0.152939
R13280 gnd.n5085 gnd.n5084 0.152939
R13281 gnd.n5084 gnd.n5065 0.152939
R13282 gnd.n5080 gnd.n5065 0.152939
R13283 gnd.n5080 gnd.n5079 0.152939
R13284 gnd.n5079 gnd.n5078 0.152939
R13285 gnd.n5078 gnd.n5069 0.152939
R13286 gnd.n5074 gnd.n5069 0.152939
R13287 gnd.n5074 gnd.n5073 0.152939
R13288 gnd.n5073 gnd.n2054 0.152939
R13289 gnd.n5188 gnd.n2054 0.152939
R13290 gnd.n5189 gnd.n5188 0.152939
R13291 gnd.n5194 gnd.n5189 0.152939
R13292 gnd.n5194 gnd.n5193 0.152939
R13293 gnd.n5193 gnd.n5192 0.152939
R13294 gnd.n5192 gnd.n5190 0.152939
R13295 gnd.n5190 gnd.n2027 0.152939
R13296 gnd.n5226 gnd.n2027 0.152939
R13297 gnd.n5227 gnd.n5226 0.152939
R13298 gnd.n5257 gnd.n5227 0.152939
R13299 gnd.n5257 gnd.n5256 0.152939
R13300 gnd.n5256 gnd.n5255 0.152939
R13301 gnd.n5255 gnd.n5228 0.152939
R13302 gnd.n5251 gnd.n5228 0.152939
R13303 gnd.n5251 gnd.n5250 0.152939
R13304 gnd.n5250 gnd.n5249 0.152939
R13305 gnd.n5249 gnd.n5231 0.152939
R13306 gnd.n5245 gnd.n5231 0.152939
R13307 gnd.n5245 gnd.n5244 0.152939
R13308 gnd.n5244 gnd.n5243 0.152939
R13309 gnd.n5243 gnd.n5237 0.152939
R13310 gnd.n5239 gnd.n5237 0.152939
R13311 gnd.n5239 gnd.n1928 0.152939
R13312 gnd.n5390 gnd.n1928 0.152939
R13313 gnd.n5391 gnd.n5390 0.152939
R13314 gnd.n5393 gnd.n5391 0.152939
R13315 gnd.n5393 gnd.n5392 0.152939
R13316 gnd.n5392 gnd.n1781 0.152939
R13317 gnd.n5499 gnd.n1781 0.152939
R13318 gnd.n5500 gnd.n5499 0.152939
R13319 gnd.n5501 gnd.n5500 0.152939
R13320 gnd.n5501 gnd.n1494 0.152939
R13321 gnd.n5820 gnd.n1494 0.152939
R13322 gnd.n5819 gnd.n1495 0.152939
R13323 gnd.n5815 gnd.n1495 0.152939
R13324 gnd.n5815 gnd.n5814 0.152939
R13325 gnd.n5814 gnd.n5813 0.152939
R13326 gnd.n5813 gnd.n1499 0.152939
R13327 gnd.n5809 gnd.n1499 0.152939
R13328 gnd.n5569 gnd.n5535 0.152939
R13329 gnd.n5569 gnd.n5568 0.152939
R13330 gnd.n5568 gnd.n5567 0.152939
R13331 gnd.n5567 gnd.n5536 0.152939
R13332 gnd.n5563 gnd.n5536 0.152939
R13333 gnd.n5563 gnd.n5562 0.152939
R13334 gnd.n5562 gnd.n5561 0.152939
R13335 gnd.n5561 gnd.n5541 0.152939
R13336 gnd.n5557 gnd.n5541 0.152939
R13337 gnd.n5557 gnd.n5556 0.152939
R13338 gnd.n5556 gnd.n5555 0.152939
R13339 gnd.n5555 gnd.n533 0.152939
R13340 gnd.n6878 gnd.n533 0.152939
R13341 gnd.n6879 gnd.n6878 0.152939
R13342 gnd.n6880 gnd.n6879 0.152939
R13343 gnd.n6880 gnd.n514 0.152939
R13344 gnd.n6905 gnd.n514 0.152939
R13345 gnd.n6906 gnd.n6905 0.152939
R13346 gnd.n6907 gnd.n6906 0.152939
R13347 gnd.n6907 gnd.n63 0.152939
R13348 gnd.n7030 gnd.n7029 0.145814
R13349 gnd.n4049 gnd.n4046 0.145814
R13350 gnd.n4049 gnd.n4048 0.145814
R13351 gnd.n7030 gnd.n63 0.145814
R13352 gnd.n6851 gnd.n78 0.136171
R13353 gnd.n4400 gnd.n4399 0.136171
R13354 gnd.n4574 gnd.n4573 0.128549
R13355 gnd.n5809 gnd.n5808 0.128549
R13356 gnd.n2722 gnd.n0 0.127478
R13357 gnd.n3302 gnd.n3301 0.0767195
R13358 gnd.n3301 gnd.n3300 0.0767195
R13359 gnd.n4671 gnd.n4574 0.063
R13360 gnd.n5808 gnd.n1504 0.063
R13361 gnd.n1672 gnd.n1504 0.0538288
R13362 gnd.n6966 gnd.n493 0.0538288
R13363 gnd.n4123 gnd.n2437 0.0538288
R13364 gnd.n4672 gnd.n4671 0.0538288
R13365 gnd.n3869 gnd.n2484 0.0477147
R13366 gnd.n3065 gnd.n2953 0.0442063
R13367 gnd.n3066 gnd.n3065 0.0442063
R13368 gnd.n3067 gnd.n3066 0.0442063
R13369 gnd.n3067 gnd.n2942 0.0442063
R13370 gnd.n3081 gnd.n2942 0.0442063
R13371 gnd.n3082 gnd.n3081 0.0442063
R13372 gnd.n3083 gnd.n3082 0.0442063
R13373 gnd.n3083 gnd.n2929 0.0442063
R13374 gnd.n3127 gnd.n2929 0.0442063
R13375 gnd.n3128 gnd.n3127 0.0442063
R13376 gnd.n3130 gnd.n2863 0.0344674
R13377 gnd.n5630 gnd.n1672 0.0344674
R13378 gnd.n5630 gnd.n1674 0.0344674
R13379 gnd.n1698 gnd.n1674 0.0344674
R13380 gnd.n1699 gnd.n1698 0.0344674
R13381 gnd.n1700 gnd.n1699 0.0344674
R13382 gnd.n1701 gnd.n1700 0.0344674
R13383 gnd.n5547 gnd.n1701 0.0344674
R13384 gnd.n5547 gnd.n1721 0.0344674
R13385 gnd.n5604 gnd.n1721 0.0344674
R13386 gnd.n5604 gnd.n1722 0.0344674
R13387 gnd.n1722 gnd.n553 0.0344674
R13388 gnd.n554 gnd.n553 0.0344674
R13389 gnd.n555 gnd.n554 0.0344674
R13390 gnd.n556 gnd.n555 0.0344674
R13391 gnd.n556 gnd.n529 0.0344674
R13392 gnd.n529 gnd.n526 0.0344674
R13393 gnd.n527 gnd.n526 0.0344674
R13394 gnd.n6891 gnd.n527 0.0344674
R13395 gnd.n6891 gnd.n502 0.0344674
R13396 gnd.n6921 gnd.n502 0.0344674
R13397 gnd.n6922 gnd.n6921 0.0344674
R13398 gnd.n6922 gnd.n497 0.0344674
R13399 gnd.n497 gnd.n495 0.0344674
R13400 gnd.n6933 gnd.n495 0.0344674
R13401 gnd.n6934 gnd.n6933 0.0344674
R13402 gnd.n6934 gnd.n92 0.0344674
R13403 gnd.n93 gnd.n92 0.0344674
R13404 gnd.n94 gnd.n93 0.0344674
R13405 gnd.n6942 gnd.n94 0.0344674
R13406 gnd.n6942 gnd.n109 0.0344674
R13407 gnd.n110 gnd.n109 0.0344674
R13408 gnd.n111 gnd.n110 0.0344674
R13409 gnd.n6949 gnd.n111 0.0344674
R13410 gnd.n6949 gnd.n129 0.0344674
R13411 gnd.n130 gnd.n129 0.0344674
R13412 gnd.n131 gnd.n130 0.0344674
R13413 gnd.n6956 gnd.n131 0.0344674
R13414 gnd.n6956 gnd.n149 0.0344674
R13415 gnd.n150 gnd.n149 0.0344674
R13416 gnd.n151 gnd.n150 0.0344674
R13417 gnd.n167 gnd.n151 0.0344674
R13418 gnd.n6966 gnd.n167 0.0344674
R13419 gnd.n4248 gnd.n2437 0.0344674
R13420 gnd.n4248 gnd.n2440 0.0344674
R13421 gnd.n2440 gnd.n2439 0.0344674
R13422 gnd.n2439 gnd.n2420 0.0344674
R13423 gnd.n2420 gnd.n2418 0.0344674
R13424 gnd.n4265 gnd.n2418 0.0344674
R13425 gnd.n4266 gnd.n4265 0.0344674
R13426 gnd.n4266 gnd.n2402 0.0344674
R13427 gnd.n2402 gnd.n2400 0.0344674
R13428 gnd.n4285 gnd.n2400 0.0344674
R13429 gnd.n4286 gnd.n4285 0.0344674
R13430 gnd.n4286 gnd.n2384 0.0344674
R13431 gnd.n2384 gnd.n2382 0.0344674
R13432 gnd.n4305 gnd.n2382 0.0344674
R13433 gnd.n4306 gnd.n4305 0.0344674
R13434 gnd.n4306 gnd.n2366 0.0344674
R13435 gnd.n2366 gnd.n2364 0.0344674
R13436 gnd.n4326 gnd.n2364 0.0344674
R13437 gnd.n4327 gnd.n4326 0.0344674
R13438 gnd.n4327 gnd.n2350 0.0344674
R13439 gnd.n2350 gnd.n2346 0.0344674
R13440 gnd.n2347 gnd.n2346 0.0344674
R13441 gnd.n2348 gnd.n2347 0.0344674
R13442 gnd.n4350 gnd.n2348 0.0344674
R13443 gnd.n4351 gnd.n4350 0.0344674
R13444 gnd.n4351 gnd.n2329 0.0344674
R13445 gnd.n2329 gnd.n1068 0.0344674
R13446 gnd.n1069 gnd.n1068 0.0344674
R13447 gnd.n1070 gnd.n1069 0.0344674
R13448 gnd.n4382 gnd.n1070 0.0344674
R13449 gnd.n4382 gnd.n1089 0.0344674
R13450 gnd.n1090 gnd.n1089 0.0344674
R13451 gnd.n1091 gnd.n1090 0.0344674
R13452 gnd.n2314 gnd.n1091 0.0344674
R13453 gnd.n2314 gnd.n1108 0.0344674
R13454 gnd.n1109 gnd.n1108 0.0344674
R13455 gnd.n1110 gnd.n1109 0.0344674
R13456 gnd.n4436 gnd.n1110 0.0344674
R13457 gnd.n4436 gnd.n1129 0.0344674
R13458 gnd.n1130 gnd.n1129 0.0344674
R13459 gnd.n1131 gnd.n1130 0.0344674
R13460 gnd.n4672 gnd.n1131 0.0344674
R13461 gnd.n4569 gnd.n4441 0.0344674
R13462 gnd.n5807 gnd.n5806 0.0344674
R13463 gnd.n4720 gnd.n4719 0.029712
R13464 gnd.n5534 gnd.n5533 0.029712
R13465 gnd.n3150 gnd.n3149 0.0269946
R13466 gnd.n3152 gnd.n3151 0.0269946
R13467 gnd.n2858 gnd.n2856 0.0269946
R13468 gnd.n3162 gnd.n3160 0.0269946
R13469 gnd.n3161 gnd.n2837 0.0269946
R13470 gnd.n3181 gnd.n3180 0.0269946
R13471 gnd.n3183 gnd.n3182 0.0269946
R13472 gnd.n2832 gnd.n2831 0.0269946
R13473 gnd.n3193 gnd.n2827 0.0269946
R13474 gnd.n3192 gnd.n2829 0.0269946
R13475 gnd.n2828 gnd.n2810 0.0269946
R13476 gnd.n3213 gnd.n2811 0.0269946
R13477 gnd.n3212 gnd.n2812 0.0269946
R13478 gnd.n3246 gnd.n2787 0.0269946
R13479 gnd.n3248 gnd.n3247 0.0269946
R13480 gnd.n3249 gnd.n2734 0.0269946
R13481 gnd.n2782 gnd.n2735 0.0269946
R13482 gnd.n2784 gnd.n2736 0.0269946
R13483 gnd.n3259 gnd.n3258 0.0269946
R13484 gnd.n3261 gnd.n3260 0.0269946
R13485 gnd.n3262 gnd.n2756 0.0269946
R13486 gnd.n3264 gnd.n2757 0.0269946
R13487 gnd.n3267 gnd.n2758 0.0269946
R13488 gnd.n3270 gnd.n3269 0.0269946
R13489 gnd.n3272 gnd.n3271 0.0269946
R13490 gnd.n3337 gnd.n2657 0.0269946
R13491 gnd.n3339 gnd.n3338 0.0269946
R13492 gnd.n3348 gnd.n2650 0.0269946
R13493 gnd.n3350 gnd.n3349 0.0269946
R13494 gnd.n3351 gnd.n2648 0.0269946
R13495 gnd.n3358 gnd.n3354 0.0269946
R13496 gnd.n3357 gnd.n3356 0.0269946
R13497 gnd.n3355 gnd.n2627 0.0269946
R13498 gnd.n3380 gnd.n2628 0.0269946
R13499 gnd.n3379 gnd.n2629 0.0269946
R13500 gnd.n3422 gnd.n2602 0.0269946
R13501 gnd.n3424 gnd.n3423 0.0269946
R13502 gnd.n3433 gnd.n2595 0.0269946
R13503 gnd.n3435 gnd.n3434 0.0269946
R13504 gnd.n3436 gnd.n2593 0.0269946
R13505 gnd.n3443 gnd.n3439 0.0269946
R13506 gnd.n3442 gnd.n3441 0.0269946
R13507 gnd.n3440 gnd.n2572 0.0269946
R13508 gnd.n3465 gnd.n2573 0.0269946
R13509 gnd.n3464 gnd.n2574 0.0269946
R13510 gnd.n3511 gnd.n2548 0.0269946
R13511 gnd.n3513 gnd.n3512 0.0269946
R13512 gnd.n3523 gnd.n2541 0.0269946
R13513 gnd.n3782 gnd.n2539 0.0269946
R13514 gnd.n3787 gnd.n3785 0.0269946
R13515 gnd.n3786 gnd.n2520 0.0269946
R13516 gnd.n3811 gnd.n3810 0.0269946
R13517 gnd.n4568 gnd.n4462 0.0225788
R13518 gnd.n4565 gnd.n4564 0.0225788
R13519 gnd.n4561 gnd.n4465 0.0225788
R13520 gnd.n4560 gnd.n4471 0.0225788
R13521 gnd.n4557 gnd.n4556 0.0225788
R13522 gnd.n4553 gnd.n4477 0.0225788
R13523 gnd.n4552 gnd.n4481 0.0225788
R13524 gnd.n4549 gnd.n4548 0.0225788
R13525 gnd.n4545 gnd.n4485 0.0225788
R13526 gnd.n4544 gnd.n4491 0.0225788
R13527 gnd.n4541 gnd.n4540 0.0225788
R13528 gnd.n4537 gnd.n4497 0.0225788
R13529 gnd.n4536 gnd.n4501 0.0225788
R13530 gnd.n4533 gnd.n4532 0.0225788
R13531 gnd.n4529 gnd.n4505 0.0225788
R13532 gnd.n4528 gnd.n4511 0.0225788
R13533 gnd.n4525 gnd.n4524 0.0225788
R13534 gnd.n4516 gnd.n2291 0.0225788
R13535 gnd.n4719 gnd.n4718 0.0225788
R13536 gnd.n5803 gnd.n1505 0.0225788
R13537 gnd.n5802 gnd.n1509 0.0225788
R13538 gnd.n5799 gnd.n5798 0.0225788
R13539 gnd.n5795 gnd.n1514 0.0225788
R13540 gnd.n5794 gnd.n1518 0.0225788
R13541 gnd.n5791 gnd.n5790 0.0225788
R13542 gnd.n5787 gnd.n1522 0.0225788
R13543 gnd.n5786 gnd.n1526 0.0225788
R13544 gnd.n5783 gnd.n5782 0.0225788
R13545 gnd.n5779 gnd.n1530 0.0225788
R13546 gnd.n5778 gnd.n1534 0.0225788
R13547 gnd.n5775 gnd.n5774 0.0225788
R13548 gnd.n5771 gnd.n1538 0.0225788
R13549 gnd.n5770 gnd.n1542 0.0225788
R13550 gnd.n5767 gnd.n5766 0.0225788
R13551 gnd.n5763 gnd.n1546 0.0225788
R13552 gnd.n5762 gnd.n1552 0.0225788
R13553 gnd.n1747 gnd.n1555 0.0225788
R13554 gnd.n5533 gnd.n1746 0.0225788
R13555 gnd.n5534 gnd.n1485 0.0218415
R13556 gnd.n4735 gnd.n4720 0.0218415
R13557 gnd.n3130 gnd.n3129 0.0202011
R13558 gnd.n3129 gnd.n3128 0.0148637
R13559 gnd.n3780 gnd.n3524 0.0144266
R13560 gnd.n3781 gnd.n3780 0.0130679
R13561 gnd.n4569 gnd.n4568 0.0123886
R13562 gnd.n4565 gnd.n4462 0.0123886
R13563 gnd.n4564 gnd.n4465 0.0123886
R13564 gnd.n4561 gnd.n4560 0.0123886
R13565 gnd.n4557 gnd.n4471 0.0123886
R13566 gnd.n4556 gnd.n4477 0.0123886
R13567 gnd.n4553 gnd.n4552 0.0123886
R13568 gnd.n4549 gnd.n4481 0.0123886
R13569 gnd.n4548 gnd.n4485 0.0123886
R13570 gnd.n4545 gnd.n4544 0.0123886
R13571 gnd.n4541 gnd.n4491 0.0123886
R13572 gnd.n4540 gnd.n4497 0.0123886
R13573 gnd.n4537 gnd.n4536 0.0123886
R13574 gnd.n4533 gnd.n4501 0.0123886
R13575 gnd.n4532 gnd.n4505 0.0123886
R13576 gnd.n4529 gnd.n4528 0.0123886
R13577 gnd.n4525 gnd.n4511 0.0123886
R13578 gnd.n4524 gnd.n4516 0.0123886
R13579 gnd.n4718 gnd.n2291 0.0123886
R13580 gnd.n5806 gnd.n1505 0.0123886
R13581 gnd.n5803 gnd.n5802 0.0123886
R13582 gnd.n5799 gnd.n1509 0.0123886
R13583 gnd.n5798 gnd.n1514 0.0123886
R13584 gnd.n5795 gnd.n5794 0.0123886
R13585 gnd.n5791 gnd.n1518 0.0123886
R13586 gnd.n5790 gnd.n1522 0.0123886
R13587 gnd.n5787 gnd.n5786 0.0123886
R13588 gnd.n5783 gnd.n1526 0.0123886
R13589 gnd.n5782 gnd.n1530 0.0123886
R13590 gnd.n5779 gnd.n5778 0.0123886
R13591 gnd.n5775 gnd.n1534 0.0123886
R13592 gnd.n5774 gnd.n1538 0.0123886
R13593 gnd.n5771 gnd.n5770 0.0123886
R13594 gnd.n5767 gnd.n1542 0.0123886
R13595 gnd.n5766 gnd.n1546 0.0123886
R13596 gnd.n5763 gnd.n5762 0.0123886
R13597 gnd.n1555 gnd.n1552 0.0123886
R13598 gnd.n1747 gnd.n1746 0.0123886
R13599 gnd.n3149 gnd.n2863 0.00797283
R13600 gnd.n3151 gnd.n3150 0.00797283
R13601 gnd.n3152 gnd.n2858 0.00797283
R13602 gnd.n3160 gnd.n2856 0.00797283
R13603 gnd.n3162 gnd.n3161 0.00797283
R13604 gnd.n3180 gnd.n2837 0.00797283
R13605 gnd.n3182 gnd.n3181 0.00797283
R13606 gnd.n3183 gnd.n2832 0.00797283
R13607 gnd.n2831 gnd.n2827 0.00797283
R13608 gnd.n3193 gnd.n3192 0.00797283
R13609 gnd.n2829 gnd.n2828 0.00797283
R13610 gnd.n2811 gnd.n2810 0.00797283
R13611 gnd.n3213 gnd.n3212 0.00797283
R13612 gnd.n2812 gnd.n2787 0.00797283
R13613 gnd.n3247 gnd.n3246 0.00797283
R13614 gnd.n3249 gnd.n3248 0.00797283
R13615 gnd.n2782 gnd.n2734 0.00797283
R13616 gnd.n2784 gnd.n2735 0.00797283
R13617 gnd.n3258 gnd.n2736 0.00797283
R13618 gnd.n3260 gnd.n3259 0.00797283
R13619 gnd.n3262 gnd.n3261 0.00797283
R13620 gnd.n3264 gnd.n2756 0.00797283
R13621 gnd.n3267 gnd.n2757 0.00797283
R13622 gnd.n3269 gnd.n2758 0.00797283
R13623 gnd.n3272 gnd.n3270 0.00797283
R13624 gnd.n3271 gnd.n2657 0.00797283
R13625 gnd.n3339 gnd.n3337 0.00797283
R13626 gnd.n3338 gnd.n2650 0.00797283
R13627 gnd.n3349 gnd.n3348 0.00797283
R13628 gnd.n3351 gnd.n3350 0.00797283
R13629 gnd.n3354 gnd.n2648 0.00797283
R13630 gnd.n3358 gnd.n3357 0.00797283
R13631 gnd.n3356 gnd.n3355 0.00797283
R13632 gnd.n2628 gnd.n2627 0.00797283
R13633 gnd.n3380 gnd.n3379 0.00797283
R13634 gnd.n2629 gnd.n2602 0.00797283
R13635 gnd.n3424 gnd.n3422 0.00797283
R13636 gnd.n3423 gnd.n2595 0.00797283
R13637 gnd.n3434 gnd.n3433 0.00797283
R13638 gnd.n3436 gnd.n3435 0.00797283
R13639 gnd.n3439 gnd.n2593 0.00797283
R13640 gnd.n3443 gnd.n3442 0.00797283
R13641 gnd.n3441 gnd.n3440 0.00797283
R13642 gnd.n2573 gnd.n2572 0.00797283
R13643 gnd.n3465 gnd.n3464 0.00797283
R13644 gnd.n2574 gnd.n2548 0.00797283
R13645 gnd.n3513 gnd.n3511 0.00797283
R13646 gnd.n3512 gnd.n2541 0.00797283
R13647 gnd.n3524 gnd.n3523 0.00797283
R13648 gnd.n3782 gnd.n3781 0.00797283
R13649 gnd.n3785 gnd.n2539 0.00797283
R13650 gnd.n3787 gnd.n3786 0.00797283
R13651 gnd.n3810 gnd.n2520 0.00797283
R13652 gnd.n3811 gnd.n2484 0.00797283
R13653 gnd.n4574 gnd.n4441 0.00593478
R13654 gnd.n5808 gnd.n5807 0.00593478
R13655 CSoutput.n19 CSoutput.t133 184.661
R13656 CSoutput.n78 CSoutput.n77 165.8
R13657 CSoutput.n76 CSoutput.n0 165.8
R13658 CSoutput.n75 CSoutput.n74 165.8
R13659 CSoutput.n73 CSoutput.n72 165.8
R13660 CSoutput.n71 CSoutput.n2 165.8
R13661 CSoutput.n69 CSoutput.n68 165.8
R13662 CSoutput.n67 CSoutput.n3 165.8
R13663 CSoutput.n66 CSoutput.n65 165.8
R13664 CSoutput.n63 CSoutput.n4 165.8
R13665 CSoutput.n61 CSoutput.n60 165.8
R13666 CSoutput.n59 CSoutput.n5 165.8
R13667 CSoutput.n58 CSoutput.n57 165.8
R13668 CSoutput.n55 CSoutput.n6 165.8
R13669 CSoutput.n54 CSoutput.n53 165.8
R13670 CSoutput.n52 CSoutput.n51 165.8
R13671 CSoutput.n50 CSoutput.n8 165.8
R13672 CSoutput.n48 CSoutput.n47 165.8
R13673 CSoutput.n46 CSoutput.n9 165.8
R13674 CSoutput.n45 CSoutput.n44 165.8
R13675 CSoutput.n42 CSoutput.n10 165.8
R13676 CSoutput.n41 CSoutput.n40 165.8
R13677 CSoutput.n39 CSoutput.n38 165.8
R13678 CSoutput.n37 CSoutput.n12 165.8
R13679 CSoutput.n35 CSoutput.n34 165.8
R13680 CSoutput.n33 CSoutput.n13 165.8
R13681 CSoutput.n32 CSoutput.n31 165.8
R13682 CSoutput.n29 CSoutput.n14 165.8
R13683 CSoutput.n28 CSoutput.n27 165.8
R13684 CSoutput.n26 CSoutput.n25 165.8
R13685 CSoutput.n24 CSoutput.n16 165.8
R13686 CSoutput.n22 CSoutput.n21 165.8
R13687 CSoutput.n20 CSoutput.n17 165.8
R13688 CSoutput.n77 CSoutput.t134 162.194
R13689 CSoutput.n18 CSoutput.t135 120.501
R13690 CSoutput.n23 CSoutput.t122 120.501
R13691 CSoutput.n15 CSoutput.t141 120.501
R13692 CSoutput.n30 CSoutput.t138 120.501
R13693 CSoutput.n36 CSoutput.t124 120.501
R13694 CSoutput.n11 CSoutput.t126 120.501
R13695 CSoutput.n43 CSoutput.t139 120.501
R13696 CSoutput.n49 CSoutput.t128 120.501
R13697 CSoutput.n7 CSoutput.t129 120.501
R13698 CSoutput.n56 CSoutput.t123 120.501
R13699 CSoutput.n62 CSoutput.t137 120.501
R13700 CSoutput.n64 CSoutput.t132 120.501
R13701 CSoutput.n70 CSoutput.t125 120.501
R13702 CSoutput.n1 CSoutput.t121 120.501
R13703 CSoutput.n270 CSoutput.n268 103.469
R13704 CSoutput.n262 CSoutput.n260 103.469
R13705 CSoutput.n255 CSoutput.n253 103.469
R13706 CSoutput.n96 CSoutput.n94 103.469
R13707 CSoutput.n88 CSoutput.n86 103.469
R13708 CSoutput.n81 CSoutput.n79 103.469
R13709 CSoutput.n272 CSoutput.n271 103.111
R13710 CSoutput.n270 CSoutput.n269 103.111
R13711 CSoutput.n266 CSoutput.n265 103.111
R13712 CSoutput.n264 CSoutput.n263 103.111
R13713 CSoutput.n262 CSoutput.n261 103.111
R13714 CSoutput.n259 CSoutput.n258 103.111
R13715 CSoutput.n257 CSoutput.n256 103.111
R13716 CSoutput.n255 CSoutput.n254 103.111
R13717 CSoutput.n96 CSoutput.n95 103.111
R13718 CSoutput.n98 CSoutput.n97 103.111
R13719 CSoutput.n100 CSoutput.n99 103.111
R13720 CSoutput.n88 CSoutput.n87 103.111
R13721 CSoutput.n90 CSoutput.n89 103.111
R13722 CSoutput.n92 CSoutput.n91 103.111
R13723 CSoutput.n81 CSoutput.n80 103.111
R13724 CSoutput.n83 CSoutput.n82 103.111
R13725 CSoutput.n85 CSoutput.n84 103.111
R13726 CSoutput.n274 CSoutput.n273 103.111
R13727 CSoutput.n302 CSoutput.n300 81.5057
R13728 CSoutput.n290 CSoutput.n288 81.5057
R13729 CSoutput.n279 CSoutput.n277 81.5057
R13730 CSoutput.n338 CSoutput.n336 81.5057
R13731 CSoutput.n326 CSoutput.n324 81.5057
R13732 CSoutput.n315 CSoutput.n313 81.5057
R13733 CSoutput.n310 CSoutput.n309 80.9324
R13734 CSoutput.n308 CSoutput.n307 80.9324
R13735 CSoutput.n306 CSoutput.n305 80.9324
R13736 CSoutput.n304 CSoutput.n303 80.9324
R13737 CSoutput.n302 CSoutput.n301 80.9324
R13738 CSoutput.n298 CSoutput.n297 80.9324
R13739 CSoutput.n296 CSoutput.n295 80.9324
R13740 CSoutput.n294 CSoutput.n293 80.9324
R13741 CSoutput.n292 CSoutput.n291 80.9324
R13742 CSoutput.n290 CSoutput.n289 80.9324
R13743 CSoutput.n287 CSoutput.n286 80.9324
R13744 CSoutput.n285 CSoutput.n284 80.9324
R13745 CSoutput.n283 CSoutput.n282 80.9324
R13746 CSoutput.n281 CSoutput.n280 80.9324
R13747 CSoutput.n279 CSoutput.n278 80.9324
R13748 CSoutput.n338 CSoutput.n337 80.9324
R13749 CSoutput.n340 CSoutput.n339 80.9324
R13750 CSoutput.n342 CSoutput.n341 80.9324
R13751 CSoutput.n344 CSoutput.n343 80.9324
R13752 CSoutput.n346 CSoutput.n345 80.9324
R13753 CSoutput.n326 CSoutput.n325 80.9324
R13754 CSoutput.n328 CSoutput.n327 80.9324
R13755 CSoutput.n330 CSoutput.n329 80.9324
R13756 CSoutput.n332 CSoutput.n331 80.9324
R13757 CSoutput.n334 CSoutput.n333 80.9324
R13758 CSoutput.n315 CSoutput.n314 80.9324
R13759 CSoutput.n317 CSoutput.n316 80.9324
R13760 CSoutput.n319 CSoutput.n318 80.9324
R13761 CSoutput.n321 CSoutput.n320 80.9324
R13762 CSoutput.n323 CSoutput.n322 80.9324
R13763 CSoutput.n25 CSoutput.n24 48.1486
R13764 CSoutput.n69 CSoutput.n3 48.1486
R13765 CSoutput.n38 CSoutput.n37 48.1486
R13766 CSoutput.n42 CSoutput.n41 48.1486
R13767 CSoutput.n51 CSoutput.n50 48.1486
R13768 CSoutput.n55 CSoutput.n54 48.1486
R13769 CSoutput.n22 CSoutput.n17 46.462
R13770 CSoutput.n72 CSoutput.n71 46.462
R13771 CSoutput.n20 CSoutput.n19 44.9055
R13772 CSoutput.n29 CSoutput.n28 43.7635
R13773 CSoutput.n65 CSoutput.n63 43.7635
R13774 CSoutput.n35 CSoutput.n13 41.7396
R13775 CSoutput.n57 CSoutput.n5 41.7396
R13776 CSoutput.n44 CSoutput.n9 37.0171
R13777 CSoutput.n48 CSoutput.n9 37.0171
R13778 CSoutput.n76 CSoutput.n75 34.9932
R13779 CSoutput.n31 CSoutput.n13 32.2947
R13780 CSoutput.n61 CSoutput.n5 32.2947
R13781 CSoutput.n30 CSoutput.n29 29.6014
R13782 CSoutput.n63 CSoutput.n62 29.6014
R13783 CSoutput.n19 CSoutput.n18 28.4085
R13784 CSoutput.n18 CSoutput.n17 25.1176
R13785 CSoutput.n72 CSoutput.n1 25.1176
R13786 CSoutput.n43 CSoutput.n42 22.0922
R13787 CSoutput.n50 CSoutput.n49 22.0922
R13788 CSoutput.n77 CSoutput.n76 21.8586
R13789 CSoutput.n37 CSoutput.n36 18.9681
R13790 CSoutput.n56 CSoutput.n55 18.9681
R13791 CSoutput.n25 CSoutput.n15 17.6292
R13792 CSoutput.n64 CSoutput.n3 17.6292
R13793 CSoutput.n24 CSoutput.n23 15.844
R13794 CSoutput.n70 CSoutput.n69 15.844
R13795 CSoutput.n38 CSoutput.n11 14.5051
R13796 CSoutput.n54 CSoutput.n7 14.5051
R13797 CSoutput.n349 CSoutput.n78 11.4982
R13798 CSoutput.n41 CSoutput.n11 11.3811
R13799 CSoutput.n51 CSoutput.n7 11.3811
R13800 CSoutput.n23 CSoutput.n22 10.0422
R13801 CSoutput.n71 CSoutput.n70 10.0422
R13802 CSoutput.n267 CSoutput.n259 9.25285
R13803 CSoutput.n93 CSoutput.n85 9.25285
R13804 CSoutput.n299 CSoutput.n287 8.98182
R13805 CSoutput.n335 CSoutput.n323 8.98182
R13806 CSoutput.n312 CSoutput.n276 8.92829
R13807 CSoutput.n28 CSoutput.n15 8.25698
R13808 CSoutput.n65 CSoutput.n64 8.25698
R13809 CSoutput.n276 CSoutput.n275 7.12641
R13810 CSoutput.n102 CSoutput.n101 7.12641
R13811 CSoutput.n36 CSoutput.n35 6.91809
R13812 CSoutput.n57 CSoutput.n56 6.91809
R13813 CSoutput.n312 CSoutput.n311 6.02792
R13814 CSoutput.n348 CSoutput.n347 6.02792
R13815 CSoutput.n349 CSoutput.n102 5.33585
R13816 CSoutput.n311 CSoutput.n310 5.25266
R13817 CSoutput.n299 CSoutput.n298 5.25266
R13818 CSoutput.n347 CSoutput.n346 5.25266
R13819 CSoutput.n335 CSoutput.n334 5.25266
R13820 CSoutput.n275 CSoutput.n274 5.1449
R13821 CSoutput.n267 CSoutput.n266 5.1449
R13822 CSoutput.n101 CSoutput.n100 5.1449
R13823 CSoutput.n93 CSoutput.n92 5.1449
R13824 CSoutput.n193 CSoutput.n146 4.5005
R13825 CSoutput.n162 CSoutput.n146 4.5005
R13826 CSoutput.n157 CSoutput.n141 4.5005
R13827 CSoutput.n157 CSoutput.n143 4.5005
R13828 CSoutput.n157 CSoutput.n140 4.5005
R13829 CSoutput.n157 CSoutput.n144 4.5005
R13830 CSoutput.n157 CSoutput.n139 4.5005
R13831 CSoutput.n157 CSoutput.t127 4.5005
R13832 CSoutput.n157 CSoutput.n138 4.5005
R13833 CSoutput.n157 CSoutput.n145 4.5005
R13834 CSoutput.n157 CSoutput.n146 4.5005
R13835 CSoutput.n155 CSoutput.n141 4.5005
R13836 CSoutput.n155 CSoutput.n143 4.5005
R13837 CSoutput.n155 CSoutput.n140 4.5005
R13838 CSoutput.n155 CSoutput.n144 4.5005
R13839 CSoutput.n155 CSoutput.n139 4.5005
R13840 CSoutput.n155 CSoutput.t127 4.5005
R13841 CSoutput.n155 CSoutput.n138 4.5005
R13842 CSoutput.n155 CSoutput.n145 4.5005
R13843 CSoutput.n155 CSoutput.n146 4.5005
R13844 CSoutput.n154 CSoutput.n141 4.5005
R13845 CSoutput.n154 CSoutput.n143 4.5005
R13846 CSoutput.n154 CSoutput.n140 4.5005
R13847 CSoutput.n154 CSoutput.n144 4.5005
R13848 CSoutput.n154 CSoutput.n139 4.5005
R13849 CSoutput.n154 CSoutput.t127 4.5005
R13850 CSoutput.n154 CSoutput.n138 4.5005
R13851 CSoutput.n154 CSoutput.n145 4.5005
R13852 CSoutput.n154 CSoutput.n146 4.5005
R13853 CSoutput.n239 CSoutput.n141 4.5005
R13854 CSoutput.n239 CSoutput.n143 4.5005
R13855 CSoutput.n239 CSoutput.n140 4.5005
R13856 CSoutput.n239 CSoutput.n144 4.5005
R13857 CSoutput.n239 CSoutput.n139 4.5005
R13858 CSoutput.n239 CSoutput.t127 4.5005
R13859 CSoutput.n239 CSoutput.n138 4.5005
R13860 CSoutput.n239 CSoutput.n145 4.5005
R13861 CSoutput.n239 CSoutput.n146 4.5005
R13862 CSoutput.n237 CSoutput.n141 4.5005
R13863 CSoutput.n237 CSoutput.n143 4.5005
R13864 CSoutput.n237 CSoutput.n140 4.5005
R13865 CSoutput.n237 CSoutput.n144 4.5005
R13866 CSoutput.n237 CSoutput.n139 4.5005
R13867 CSoutput.n237 CSoutput.t127 4.5005
R13868 CSoutput.n237 CSoutput.n138 4.5005
R13869 CSoutput.n237 CSoutput.n145 4.5005
R13870 CSoutput.n235 CSoutput.n141 4.5005
R13871 CSoutput.n235 CSoutput.n143 4.5005
R13872 CSoutput.n235 CSoutput.n140 4.5005
R13873 CSoutput.n235 CSoutput.n144 4.5005
R13874 CSoutput.n235 CSoutput.n139 4.5005
R13875 CSoutput.n235 CSoutput.t127 4.5005
R13876 CSoutput.n235 CSoutput.n138 4.5005
R13877 CSoutput.n235 CSoutput.n145 4.5005
R13878 CSoutput.n165 CSoutput.n141 4.5005
R13879 CSoutput.n165 CSoutput.n143 4.5005
R13880 CSoutput.n165 CSoutput.n140 4.5005
R13881 CSoutput.n165 CSoutput.n144 4.5005
R13882 CSoutput.n165 CSoutput.n139 4.5005
R13883 CSoutput.n165 CSoutput.t127 4.5005
R13884 CSoutput.n165 CSoutput.n138 4.5005
R13885 CSoutput.n165 CSoutput.n145 4.5005
R13886 CSoutput.n165 CSoutput.n146 4.5005
R13887 CSoutput.n164 CSoutput.n141 4.5005
R13888 CSoutput.n164 CSoutput.n143 4.5005
R13889 CSoutput.n164 CSoutput.n140 4.5005
R13890 CSoutput.n164 CSoutput.n144 4.5005
R13891 CSoutput.n164 CSoutput.n139 4.5005
R13892 CSoutput.n164 CSoutput.t127 4.5005
R13893 CSoutput.n164 CSoutput.n138 4.5005
R13894 CSoutput.n164 CSoutput.n145 4.5005
R13895 CSoutput.n164 CSoutput.n146 4.5005
R13896 CSoutput.n168 CSoutput.n141 4.5005
R13897 CSoutput.n168 CSoutput.n143 4.5005
R13898 CSoutput.n168 CSoutput.n140 4.5005
R13899 CSoutput.n168 CSoutput.n144 4.5005
R13900 CSoutput.n168 CSoutput.n139 4.5005
R13901 CSoutput.n168 CSoutput.t127 4.5005
R13902 CSoutput.n168 CSoutput.n138 4.5005
R13903 CSoutput.n168 CSoutput.n145 4.5005
R13904 CSoutput.n168 CSoutput.n146 4.5005
R13905 CSoutput.n167 CSoutput.n141 4.5005
R13906 CSoutput.n167 CSoutput.n143 4.5005
R13907 CSoutput.n167 CSoutput.n140 4.5005
R13908 CSoutput.n167 CSoutput.n144 4.5005
R13909 CSoutput.n167 CSoutput.n139 4.5005
R13910 CSoutput.n167 CSoutput.t127 4.5005
R13911 CSoutput.n167 CSoutput.n138 4.5005
R13912 CSoutput.n167 CSoutput.n145 4.5005
R13913 CSoutput.n167 CSoutput.n146 4.5005
R13914 CSoutput.n150 CSoutput.n141 4.5005
R13915 CSoutput.n150 CSoutput.n143 4.5005
R13916 CSoutput.n150 CSoutput.n140 4.5005
R13917 CSoutput.n150 CSoutput.n144 4.5005
R13918 CSoutput.n150 CSoutput.n139 4.5005
R13919 CSoutput.n150 CSoutput.t127 4.5005
R13920 CSoutput.n150 CSoutput.n138 4.5005
R13921 CSoutput.n150 CSoutput.n145 4.5005
R13922 CSoutput.n150 CSoutput.n146 4.5005
R13923 CSoutput.n242 CSoutput.n141 4.5005
R13924 CSoutput.n242 CSoutput.n143 4.5005
R13925 CSoutput.n242 CSoutput.n140 4.5005
R13926 CSoutput.n242 CSoutput.n144 4.5005
R13927 CSoutput.n242 CSoutput.n139 4.5005
R13928 CSoutput.n242 CSoutput.t127 4.5005
R13929 CSoutput.n242 CSoutput.n138 4.5005
R13930 CSoutput.n242 CSoutput.n145 4.5005
R13931 CSoutput.n242 CSoutput.n146 4.5005
R13932 CSoutput.n229 CSoutput.n200 4.5005
R13933 CSoutput.n229 CSoutput.n206 4.5005
R13934 CSoutput.n187 CSoutput.n176 4.5005
R13935 CSoutput.n187 CSoutput.n178 4.5005
R13936 CSoutput.n187 CSoutput.n175 4.5005
R13937 CSoutput.n187 CSoutput.n179 4.5005
R13938 CSoutput.n187 CSoutput.n174 4.5005
R13939 CSoutput.n187 CSoutput.t120 4.5005
R13940 CSoutput.n187 CSoutput.n173 4.5005
R13941 CSoutput.n187 CSoutput.n180 4.5005
R13942 CSoutput.n229 CSoutput.n187 4.5005
R13943 CSoutput.n208 CSoutput.n176 4.5005
R13944 CSoutput.n208 CSoutput.n178 4.5005
R13945 CSoutput.n208 CSoutput.n175 4.5005
R13946 CSoutput.n208 CSoutput.n179 4.5005
R13947 CSoutput.n208 CSoutput.n174 4.5005
R13948 CSoutput.n208 CSoutput.t120 4.5005
R13949 CSoutput.n208 CSoutput.n173 4.5005
R13950 CSoutput.n208 CSoutput.n180 4.5005
R13951 CSoutput.n229 CSoutput.n208 4.5005
R13952 CSoutput.n186 CSoutput.n176 4.5005
R13953 CSoutput.n186 CSoutput.n178 4.5005
R13954 CSoutput.n186 CSoutput.n175 4.5005
R13955 CSoutput.n186 CSoutput.n179 4.5005
R13956 CSoutput.n186 CSoutput.n174 4.5005
R13957 CSoutput.n186 CSoutput.t120 4.5005
R13958 CSoutput.n186 CSoutput.n173 4.5005
R13959 CSoutput.n186 CSoutput.n180 4.5005
R13960 CSoutput.n229 CSoutput.n186 4.5005
R13961 CSoutput.n210 CSoutput.n176 4.5005
R13962 CSoutput.n210 CSoutput.n178 4.5005
R13963 CSoutput.n210 CSoutput.n175 4.5005
R13964 CSoutput.n210 CSoutput.n179 4.5005
R13965 CSoutput.n210 CSoutput.n174 4.5005
R13966 CSoutput.n210 CSoutput.t120 4.5005
R13967 CSoutput.n210 CSoutput.n173 4.5005
R13968 CSoutput.n210 CSoutput.n180 4.5005
R13969 CSoutput.n229 CSoutput.n210 4.5005
R13970 CSoutput.n176 CSoutput.n171 4.5005
R13971 CSoutput.n178 CSoutput.n171 4.5005
R13972 CSoutput.n175 CSoutput.n171 4.5005
R13973 CSoutput.n179 CSoutput.n171 4.5005
R13974 CSoutput.n174 CSoutput.n171 4.5005
R13975 CSoutput.t120 CSoutput.n171 4.5005
R13976 CSoutput.n173 CSoutput.n171 4.5005
R13977 CSoutput.n180 CSoutput.n171 4.5005
R13978 CSoutput.n232 CSoutput.n176 4.5005
R13979 CSoutput.n232 CSoutput.n178 4.5005
R13980 CSoutput.n232 CSoutput.n175 4.5005
R13981 CSoutput.n232 CSoutput.n179 4.5005
R13982 CSoutput.n232 CSoutput.n174 4.5005
R13983 CSoutput.n232 CSoutput.t120 4.5005
R13984 CSoutput.n232 CSoutput.n173 4.5005
R13985 CSoutput.n232 CSoutput.n180 4.5005
R13986 CSoutput.n230 CSoutput.n176 4.5005
R13987 CSoutput.n230 CSoutput.n178 4.5005
R13988 CSoutput.n230 CSoutput.n175 4.5005
R13989 CSoutput.n230 CSoutput.n179 4.5005
R13990 CSoutput.n230 CSoutput.n174 4.5005
R13991 CSoutput.n230 CSoutput.t120 4.5005
R13992 CSoutput.n230 CSoutput.n173 4.5005
R13993 CSoutput.n230 CSoutput.n180 4.5005
R13994 CSoutput.n230 CSoutput.n229 4.5005
R13995 CSoutput.n212 CSoutput.n176 4.5005
R13996 CSoutput.n212 CSoutput.n178 4.5005
R13997 CSoutput.n212 CSoutput.n175 4.5005
R13998 CSoutput.n212 CSoutput.n179 4.5005
R13999 CSoutput.n212 CSoutput.n174 4.5005
R14000 CSoutput.n212 CSoutput.t120 4.5005
R14001 CSoutput.n212 CSoutput.n173 4.5005
R14002 CSoutput.n212 CSoutput.n180 4.5005
R14003 CSoutput.n229 CSoutput.n212 4.5005
R14004 CSoutput.n184 CSoutput.n176 4.5005
R14005 CSoutput.n184 CSoutput.n178 4.5005
R14006 CSoutput.n184 CSoutput.n175 4.5005
R14007 CSoutput.n184 CSoutput.n179 4.5005
R14008 CSoutput.n184 CSoutput.n174 4.5005
R14009 CSoutput.n184 CSoutput.t120 4.5005
R14010 CSoutput.n184 CSoutput.n173 4.5005
R14011 CSoutput.n184 CSoutput.n180 4.5005
R14012 CSoutput.n229 CSoutput.n184 4.5005
R14013 CSoutput.n214 CSoutput.n176 4.5005
R14014 CSoutput.n214 CSoutput.n178 4.5005
R14015 CSoutput.n214 CSoutput.n175 4.5005
R14016 CSoutput.n214 CSoutput.n179 4.5005
R14017 CSoutput.n214 CSoutput.n174 4.5005
R14018 CSoutput.n214 CSoutput.t120 4.5005
R14019 CSoutput.n214 CSoutput.n173 4.5005
R14020 CSoutput.n214 CSoutput.n180 4.5005
R14021 CSoutput.n229 CSoutput.n214 4.5005
R14022 CSoutput.n183 CSoutput.n176 4.5005
R14023 CSoutput.n183 CSoutput.n178 4.5005
R14024 CSoutput.n183 CSoutput.n175 4.5005
R14025 CSoutput.n183 CSoutput.n179 4.5005
R14026 CSoutput.n183 CSoutput.n174 4.5005
R14027 CSoutput.n183 CSoutput.t120 4.5005
R14028 CSoutput.n183 CSoutput.n173 4.5005
R14029 CSoutput.n183 CSoutput.n180 4.5005
R14030 CSoutput.n229 CSoutput.n183 4.5005
R14031 CSoutput.n228 CSoutput.n176 4.5005
R14032 CSoutput.n228 CSoutput.n178 4.5005
R14033 CSoutput.n228 CSoutput.n175 4.5005
R14034 CSoutput.n228 CSoutput.n179 4.5005
R14035 CSoutput.n228 CSoutput.n174 4.5005
R14036 CSoutput.n228 CSoutput.t120 4.5005
R14037 CSoutput.n228 CSoutput.n173 4.5005
R14038 CSoutput.n228 CSoutput.n180 4.5005
R14039 CSoutput.n229 CSoutput.n228 4.5005
R14040 CSoutput.n227 CSoutput.n112 4.5005
R14041 CSoutput.n128 CSoutput.n112 4.5005
R14042 CSoutput.n123 CSoutput.n107 4.5005
R14043 CSoutput.n123 CSoutput.n109 4.5005
R14044 CSoutput.n123 CSoutput.n106 4.5005
R14045 CSoutput.n123 CSoutput.n110 4.5005
R14046 CSoutput.n123 CSoutput.n105 4.5005
R14047 CSoutput.n123 CSoutput.t140 4.5005
R14048 CSoutput.n123 CSoutput.n104 4.5005
R14049 CSoutput.n123 CSoutput.n111 4.5005
R14050 CSoutput.n123 CSoutput.n112 4.5005
R14051 CSoutput.n121 CSoutput.n107 4.5005
R14052 CSoutput.n121 CSoutput.n109 4.5005
R14053 CSoutput.n121 CSoutput.n106 4.5005
R14054 CSoutput.n121 CSoutput.n110 4.5005
R14055 CSoutput.n121 CSoutput.n105 4.5005
R14056 CSoutput.n121 CSoutput.t140 4.5005
R14057 CSoutput.n121 CSoutput.n104 4.5005
R14058 CSoutput.n121 CSoutput.n111 4.5005
R14059 CSoutput.n121 CSoutput.n112 4.5005
R14060 CSoutput.n120 CSoutput.n107 4.5005
R14061 CSoutput.n120 CSoutput.n109 4.5005
R14062 CSoutput.n120 CSoutput.n106 4.5005
R14063 CSoutput.n120 CSoutput.n110 4.5005
R14064 CSoutput.n120 CSoutput.n105 4.5005
R14065 CSoutput.n120 CSoutput.t140 4.5005
R14066 CSoutput.n120 CSoutput.n104 4.5005
R14067 CSoutput.n120 CSoutput.n111 4.5005
R14068 CSoutput.n120 CSoutput.n112 4.5005
R14069 CSoutput.n249 CSoutput.n107 4.5005
R14070 CSoutput.n249 CSoutput.n109 4.5005
R14071 CSoutput.n249 CSoutput.n106 4.5005
R14072 CSoutput.n249 CSoutput.n110 4.5005
R14073 CSoutput.n249 CSoutput.n105 4.5005
R14074 CSoutput.n249 CSoutput.t140 4.5005
R14075 CSoutput.n249 CSoutput.n104 4.5005
R14076 CSoutput.n249 CSoutput.n111 4.5005
R14077 CSoutput.n249 CSoutput.n112 4.5005
R14078 CSoutput.n247 CSoutput.n107 4.5005
R14079 CSoutput.n247 CSoutput.n109 4.5005
R14080 CSoutput.n247 CSoutput.n106 4.5005
R14081 CSoutput.n247 CSoutput.n110 4.5005
R14082 CSoutput.n247 CSoutput.n105 4.5005
R14083 CSoutput.n247 CSoutput.t140 4.5005
R14084 CSoutput.n247 CSoutput.n104 4.5005
R14085 CSoutput.n247 CSoutput.n111 4.5005
R14086 CSoutput.n245 CSoutput.n107 4.5005
R14087 CSoutput.n245 CSoutput.n109 4.5005
R14088 CSoutput.n245 CSoutput.n106 4.5005
R14089 CSoutput.n245 CSoutput.n110 4.5005
R14090 CSoutput.n245 CSoutput.n105 4.5005
R14091 CSoutput.n245 CSoutput.t140 4.5005
R14092 CSoutput.n245 CSoutput.n104 4.5005
R14093 CSoutput.n245 CSoutput.n111 4.5005
R14094 CSoutput.n131 CSoutput.n107 4.5005
R14095 CSoutput.n131 CSoutput.n109 4.5005
R14096 CSoutput.n131 CSoutput.n106 4.5005
R14097 CSoutput.n131 CSoutput.n110 4.5005
R14098 CSoutput.n131 CSoutput.n105 4.5005
R14099 CSoutput.n131 CSoutput.t140 4.5005
R14100 CSoutput.n131 CSoutput.n104 4.5005
R14101 CSoutput.n131 CSoutput.n111 4.5005
R14102 CSoutput.n131 CSoutput.n112 4.5005
R14103 CSoutput.n130 CSoutput.n107 4.5005
R14104 CSoutput.n130 CSoutput.n109 4.5005
R14105 CSoutput.n130 CSoutput.n106 4.5005
R14106 CSoutput.n130 CSoutput.n110 4.5005
R14107 CSoutput.n130 CSoutput.n105 4.5005
R14108 CSoutput.n130 CSoutput.t140 4.5005
R14109 CSoutput.n130 CSoutput.n104 4.5005
R14110 CSoutput.n130 CSoutput.n111 4.5005
R14111 CSoutput.n130 CSoutput.n112 4.5005
R14112 CSoutput.n134 CSoutput.n107 4.5005
R14113 CSoutput.n134 CSoutput.n109 4.5005
R14114 CSoutput.n134 CSoutput.n106 4.5005
R14115 CSoutput.n134 CSoutput.n110 4.5005
R14116 CSoutput.n134 CSoutput.n105 4.5005
R14117 CSoutput.n134 CSoutput.t140 4.5005
R14118 CSoutput.n134 CSoutput.n104 4.5005
R14119 CSoutput.n134 CSoutput.n111 4.5005
R14120 CSoutput.n134 CSoutput.n112 4.5005
R14121 CSoutput.n133 CSoutput.n107 4.5005
R14122 CSoutput.n133 CSoutput.n109 4.5005
R14123 CSoutput.n133 CSoutput.n106 4.5005
R14124 CSoutput.n133 CSoutput.n110 4.5005
R14125 CSoutput.n133 CSoutput.n105 4.5005
R14126 CSoutput.n133 CSoutput.t140 4.5005
R14127 CSoutput.n133 CSoutput.n104 4.5005
R14128 CSoutput.n133 CSoutput.n111 4.5005
R14129 CSoutput.n133 CSoutput.n112 4.5005
R14130 CSoutput.n116 CSoutput.n107 4.5005
R14131 CSoutput.n116 CSoutput.n109 4.5005
R14132 CSoutput.n116 CSoutput.n106 4.5005
R14133 CSoutput.n116 CSoutput.n110 4.5005
R14134 CSoutput.n116 CSoutput.n105 4.5005
R14135 CSoutput.n116 CSoutput.t140 4.5005
R14136 CSoutput.n116 CSoutput.n104 4.5005
R14137 CSoutput.n116 CSoutput.n111 4.5005
R14138 CSoutput.n116 CSoutput.n112 4.5005
R14139 CSoutput.n252 CSoutput.n107 4.5005
R14140 CSoutput.n252 CSoutput.n109 4.5005
R14141 CSoutput.n252 CSoutput.n106 4.5005
R14142 CSoutput.n252 CSoutput.n110 4.5005
R14143 CSoutput.n252 CSoutput.n105 4.5005
R14144 CSoutput.n252 CSoutput.t140 4.5005
R14145 CSoutput.n252 CSoutput.n104 4.5005
R14146 CSoutput.n252 CSoutput.n111 4.5005
R14147 CSoutput.n252 CSoutput.n112 4.5005
R14148 CSoutput.n275 CSoutput.n267 4.10845
R14149 CSoutput.n101 CSoutput.n93 4.10845
R14150 CSoutput.n273 CSoutput.t2 4.06363
R14151 CSoutput.n273 CSoutput.t35 4.06363
R14152 CSoutput.n271 CSoutput.t32 4.06363
R14153 CSoutput.n271 CSoutput.t28 4.06363
R14154 CSoutput.n269 CSoutput.t119 4.06363
R14155 CSoutput.n269 CSoutput.t34 4.06363
R14156 CSoutput.n268 CSoutput.t114 4.06363
R14157 CSoutput.n268 CSoutput.t6 4.06363
R14158 CSoutput.n265 CSoutput.t113 4.06363
R14159 CSoutput.n265 CSoutput.t17 4.06363
R14160 CSoutput.n263 CSoutput.t11 4.06363
R14161 CSoutput.n263 CSoutput.t36 4.06363
R14162 CSoutput.n261 CSoutput.t20 4.06363
R14163 CSoutput.n261 CSoutput.t24 4.06363
R14164 CSoutput.n260 CSoutput.t15 4.06363
R14165 CSoutput.n260 CSoutput.t23 4.06363
R14166 CSoutput.n258 CSoutput.t25 4.06363
R14167 CSoutput.n258 CSoutput.t16 4.06363
R14168 CSoutput.n256 CSoutput.t12 4.06363
R14169 CSoutput.n256 CSoutput.t1 4.06363
R14170 CSoutput.n254 CSoutput.t29 4.06363
R14171 CSoutput.n254 CSoutput.t31 4.06363
R14172 CSoutput.n253 CSoutput.t22 4.06363
R14173 CSoutput.n253 CSoutput.t14 4.06363
R14174 CSoutput.n94 CSoutput.t4 4.06363
R14175 CSoutput.n94 CSoutput.t33 4.06363
R14176 CSoutput.n95 CSoutput.t18 4.06363
R14177 CSoutput.n95 CSoutput.t115 4.06363
R14178 CSoutput.n97 CSoutput.t27 4.06363
R14179 CSoutput.n97 CSoutput.t10 4.06363
R14180 CSoutput.n99 CSoutput.t26 4.06363
R14181 CSoutput.n99 CSoutput.t8 4.06363
R14182 CSoutput.n86 CSoutput.t0 4.06363
R14183 CSoutput.n86 CSoutput.t5 4.06363
R14184 CSoutput.n87 CSoutput.t111 4.06363
R14185 CSoutput.n87 CSoutput.t21 4.06363
R14186 CSoutput.n89 CSoutput.t118 4.06363
R14187 CSoutput.n89 CSoutput.t13 4.06363
R14188 CSoutput.n91 CSoutput.t112 4.06363
R14189 CSoutput.n91 CSoutput.t3 4.06363
R14190 CSoutput.n79 CSoutput.t9 4.06363
R14191 CSoutput.n79 CSoutput.t110 4.06363
R14192 CSoutput.n80 CSoutput.t116 4.06363
R14193 CSoutput.n80 CSoutput.t117 4.06363
R14194 CSoutput.n82 CSoutput.t7 4.06363
R14195 CSoutput.n82 CSoutput.t19 4.06363
R14196 CSoutput.n84 CSoutput.t37 4.06363
R14197 CSoutput.n84 CSoutput.t30 4.06363
R14198 CSoutput.n44 CSoutput.n43 3.79402
R14199 CSoutput.n49 CSoutput.n48 3.79402
R14200 CSoutput.n311 CSoutput.n299 3.72967
R14201 CSoutput.n347 CSoutput.n335 3.72967
R14202 CSoutput.n349 CSoutput.n348 3.57343
R14203 CSoutput.n309 CSoutput.t55 2.82907
R14204 CSoutput.n309 CSoutput.t59 2.82907
R14205 CSoutput.n307 CSoutput.t54 2.82907
R14206 CSoutput.n307 CSoutput.t109 2.82907
R14207 CSoutput.n305 CSoutput.t70 2.82907
R14208 CSoutput.n305 CSoutput.t49 2.82907
R14209 CSoutput.n303 CSoutput.t42 2.82907
R14210 CSoutput.n303 CSoutput.t90 2.82907
R14211 CSoutput.n301 CSoutput.t61 2.82907
R14212 CSoutput.n301 CSoutput.t64 2.82907
R14213 CSoutput.n300 CSoutput.t48 2.82907
R14214 CSoutput.n300 CSoutput.t100 2.82907
R14215 CSoutput.n297 CSoutput.t41 2.82907
R14216 CSoutput.n297 CSoutput.t88 2.82907
R14217 CSoutput.n295 CSoutput.t86 2.82907
R14218 CSoutput.n295 CSoutput.t74 2.82907
R14219 CSoutput.n293 CSoutput.t99 2.82907
R14220 CSoutput.n293 CSoutput.t40 2.82907
R14221 CSoutput.n291 CSoutput.t39 2.82907
R14222 CSoutput.n291 CSoutput.t92 2.82907
R14223 CSoutput.n289 CSoutput.t47 2.82907
R14224 CSoutput.n289 CSoutput.t98 2.82907
R14225 CSoutput.n288 CSoutput.t105 2.82907
R14226 CSoutput.n288 CSoutput.t38 2.82907
R14227 CSoutput.n286 CSoutput.t77 2.82907
R14228 CSoutput.n286 CSoutput.t84 2.82907
R14229 CSoutput.n284 CSoutput.t69 2.82907
R14230 CSoutput.n284 CSoutput.t97 2.82907
R14231 CSoutput.n282 CSoutput.t80 2.82907
R14232 CSoutput.n282 CSoutput.t63 2.82907
R14233 CSoutput.n280 CSoutput.t57 2.82907
R14234 CSoutput.n280 CSoutput.t71 2.82907
R14235 CSoutput.n278 CSoutput.t62 2.82907
R14236 CSoutput.n278 CSoutput.t67 2.82907
R14237 CSoutput.n277 CSoutput.t68 2.82907
R14238 CSoutput.n277 CSoutput.t108 2.82907
R14239 CSoutput.n336 CSoutput.t76 2.82907
R14240 CSoutput.n336 CSoutput.t94 2.82907
R14241 CSoutput.n337 CSoutput.t56 2.82907
R14242 CSoutput.n337 CSoutput.t66 2.82907
R14243 CSoutput.n339 CSoutput.t72 2.82907
R14244 CSoutput.n339 CSoutput.t83 2.82907
R14245 CSoutput.n341 CSoutput.t95 2.82907
R14246 CSoutput.n341 CSoutput.t75 2.82907
R14247 CSoutput.n343 CSoutput.t79 2.82907
R14248 CSoutput.n343 CSoutput.t104 2.82907
R14249 CSoutput.n345 CSoutput.t44 2.82907
R14250 CSoutput.n345 CSoutput.t60 2.82907
R14251 CSoutput.n324 CSoutput.t50 2.82907
R14252 CSoutput.n324 CSoutput.t45 2.82907
R14253 CSoutput.n325 CSoutput.t43 2.82907
R14254 CSoutput.n325 CSoutput.t106 2.82907
R14255 CSoutput.n327 CSoutput.t107 2.82907
R14256 CSoutput.n327 CSoutput.t51 2.82907
R14257 CSoutput.n329 CSoutput.t52 2.82907
R14258 CSoutput.n329 CSoutput.t81 2.82907
R14259 CSoutput.n331 CSoutput.t82 2.82907
R14260 CSoutput.n331 CSoutput.t102 2.82907
R14261 CSoutput.n333 CSoutput.t103 2.82907
R14262 CSoutput.n333 CSoutput.t96 2.82907
R14263 CSoutput.n313 CSoutput.t58 2.82907
R14264 CSoutput.n313 CSoutput.t87 2.82907
R14265 CSoutput.n314 CSoutput.t85 2.82907
R14266 CSoutput.n314 CSoutput.t73 2.82907
R14267 CSoutput.n316 CSoutput.t91 2.82907
R14268 CSoutput.n316 CSoutput.t65 2.82907
R14269 CSoutput.n318 CSoutput.t78 2.82907
R14270 CSoutput.n318 CSoutput.t101 2.82907
R14271 CSoutput.n320 CSoutput.t53 2.82907
R14272 CSoutput.n320 CSoutput.t89 2.82907
R14273 CSoutput.n322 CSoutput.t46 2.82907
R14274 CSoutput.n322 CSoutput.t93 2.82907
R14275 CSoutput.n348 CSoutput.n312 2.75627
R14276 CSoutput.n75 CSoutput.n1 2.45513
R14277 CSoutput.n193 CSoutput.n191 2.251
R14278 CSoutput.n193 CSoutput.n190 2.251
R14279 CSoutput.n193 CSoutput.n189 2.251
R14280 CSoutput.n193 CSoutput.n188 2.251
R14281 CSoutput.n162 CSoutput.n161 2.251
R14282 CSoutput.n162 CSoutput.n160 2.251
R14283 CSoutput.n162 CSoutput.n159 2.251
R14284 CSoutput.n162 CSoutput.n158 2.251
R14285 CSoutput.n235 CSoutput.n234 2.251
R14286 CSoutput.n200 CSoutput.n198 2.251
R14287 CSoutput.n200 CSoutput.n197 2.251
R14288 CSoutput.n200 CSoutput.n196 2.251
R14289 CSoutput.n218 CSoutput.n200 2.251
R14290 CSoutput.n206 CSoutput.n205 2.251
R14291 CSoutput.n206 CSoutput.n204 2.251
R14292 CSoutput.n206 CSoutput.n203 2.251
R14293 CSoutput.n206 CSoutput.n202 2.251
R14294 CSoutput.n232 CSoutput.n172 2.251
R14295 CSoutput.n227 CSoutput.n225 2.251
R14296 CSoutput.n227 CSoutput.n224 2.251
R14297 CSoutput.n227 CSoutput.n223 2.251
R14298 CSoutput.n227 CSoutput.n222 2.251
R14299 CSoutput.n128 CSoutput.n127 2.251
R14300 CSoutput.n128 CSoutput.n126 2.251
R14301 CSoutput.n128 CSoutput.n125 2.251
R14302 CSoutput.n128 CSoutput.n124 2.251
R14303 CSoutput.n245 CSoutput.n244 2.251
R14304 CSoutput.n162 CSoutput.n142 2.2505
R14305 CSoutput.n157 CSoutput.n142 2.2505
R14306 CSoutput.n155 CSoutput.n142 2.2505
R14307 CSoutput.n154 CSoutput.n142 2.2505
R14308 CSoutput.n239 CSoutput.n142 2.2505
R14309 CSoutput.n237 CSoutput.n142 2.2505
R14310 CSoutput.n235 CSoutput.n142 2.2505
R14311 CSoutput.n165 CSoutput.n142 2.2505
R14312 CSoutput.n164 CSoutput.n142 2.2505
R14313 CSoutput.n168 CSoutput.n142 2.2505
R14314 CSoutput.n167 CSoutput.n142 2.2505
R14315 CSoutput.n150 CSoutput.n142 2.2505
R14316 CSoutput.n242 CSoutput.n142 2.2505
R14317 CSoutput.n242 CSoutput.n241 2.2505
R14318 CSoutput.n206 CSoutput.n177 2.2505
R14319 CSoutput.n187 CSoutput.n177 2.2505
R14320 CSoutput.n208 CSoutput.n177 2.2505
R14321 CSoutput.n186 CSoutput.n177 2.2505
R14322 CSoutput.n210 CSoutput.n177 2.2505
R14323 CSoutput.n177 CSoutput.n171 2.2505
R14324 CSoutput.n232 CSoutput.n177 2.2505
R14325 CSoutput.n230 CSoutput.n177 2.2505
R14326 CSoutput.n212 CSoutput.n177 2.2505
R14327 CSoutput.n184 CSoutput.n177 2.2505
R14328 CSoutput.n214 CSoutput.n177 2.2505
R14329 CSoutput.n183 CSoutput.n177 2.2505
R14330 CSoutput.n228 CSoutput.n177 2.2505
R14331 CSoutput.n228 CSoutput.n181 2.2505
R14332 CSoutput.n128 CSoutput.n108 2.2505
R14333 CSoutput.n123 CSoutput.n108 2.2505
R14334 CSoutput.n121 CSoutput.n108 2.2505
R14335 CSoutput.n120 CSoutput.n108 2.2505
R14336 CSoutput.n249 CSoutput.n108 2.2505
R14337 CSoutput.n247 CSoutput.n108 2.2505
R14338 CSoutput.n245 CSoutput.n108 2.2505
R14339 CSoutput.n131 CSoutput.n108 2.2505
R14340 CSoutput.n130 CSoutput.n108 2.2505
R14341 CSoutput.n134 CSoutput.n108 2.2505
R14342 CSoutput.n133 CSoutput.n108 2.2505
R14343 CSoutput.n116 CSoutput.n108 2.2505
R14344 CSoutput.n252 CSoutput.n108 2.2505
R14345 CSoutput.n252 CSoutput.n251 2.2505
R14346 CSoutput.n170 CSoutput.n163 2.25024
R14347 CSoutput.n170 CSoutput.n156 2.25024
R14348 CSoutput.n238 CSoutput.n170 2.25024
R14349 CSoutput.n170 CSoutput.n166 2.25024
R14350 CSoutput.n170 CSoutput.n169 2.25024
R14351 CSoutput.n170 CSoutput.n137 2.25024
R14352 CSoutput.n220 CSoutput.n217 2.25024
R14353 CSoutput.n220 CSoutput.n216 2.25024
R14354 CSoutput.n220 CSoutput.n215 2.25024
R14355 CSoutput.n220 CSoutput.n182 2.25024
R14356 CSoutput.n220 CSoutput.n219 2.25024
R14357 CSoutput.n221 CSoutput.n220 2.25024
R14358 CSoutput.n136 CSoutput.n129 2.25024
R14359 CSoutput.n136 CSoutput.n122 2.25024
R14360 CSoutput.n248 CSoutput.n136 2.25024
R14361 CSoutput.n136 CSoutput.n132 2.25024
R14362 CSoutput.n136 CSoutput.n135 2.25024
R14363 CSoutput.n136 CSoutput.n103 2.25024
R14364 CSoutput.n276 CSoutput.n102 1.95131
R14365 CSoutput.n237 CSoutput.n147 1.50111
R14366 CSoutput.n185 CSoutput.n171 1.50111
R14367 CSoutput.n247 CSoutput.n113 1.50111
R14368 CSoutput.n193 CSoutput.n192 1.501
R14369 CSoutput.n200 CSoutput.n199 1.501
R14370 CSoutput.n227 CSoutput.n226 1.501
R14371 CSoutput.n241 CSoutput.n152 1.12536
R14372 CSoutput.n241 CSoutput.n153 1.12536
R14373 CSoutput.n241 CSoutput.n240 1.12536
R14374 CSoutput.n201 CSoutput.n181 1.12536
R14375 CSoutput.n207 CSoutput.n181 1.12536
R14376 CSoutput.n209 CSoutput.n181 1.12536
R14377 CSoutput.n251 CSoutput.n118 1.12536
R14378 CSoutput.n251 CSoutput.n119 1.12536
R14379 CSoutput.n251 CSoutput.n250 1.12536
R14380 CSoutput.n241 CSoutput.n148 1.12536
R14381 CSoutput.n241 CSoutput.n149 1.12536
R14382 CSoutput.n241 CSoutput.n151 1.12536
R14383 CSoutput.n231 CSoutput.n181 1.12536
R14384 CSoutput.n211 CSoutput.n181 1.12536
R14385 CSoutput.n213 CSoutput.n181 1.12536
R14386 CSoutput.n251 CSoutput.n114 1.12536
R14387 CSoutput.n251 CSoutput.n115 1.12536
R14388 CSoutput.n251 CSoutput.n117 1.12536
R14389 CSoutput.n31 CSoutput.n30 0.669944
R14390 CSoutput.n62 CSoutput.n61 0.669944
R14391 CSoutput.n304 CSoutput.n302 0.573776
R14392 CSoutput.n306 CSoutput.n304 0.573776
R14393 CSoutput.n308 CSoutput.n306 0.573776
R14394 CSoutput.n310 CSoutput.n308 0.573776
R14395 CSoutput.n292 CSoutput.n290 0.573776
R14396 CSoutput.n294 CSoutput.n292 0.573776
R14397 CSoutput.n296 CSoutput.n294 0.573776
R14398 CSoutput.n298 CSoutput.n296 0.573776
R14399 CSoutput.n281 CSoutput.n279 0.573776
R14400 CSoutput.n283 CSoutput.n281 0.573776
R14401 CSoutput.n285 CSoutput.n283 0.573776
R14402 CSoutput.n287 CSoutput.n285 0.573776
R14403 CSoutput.n346 CSoutput.n344 0.573776
R14404 CSoutput.n344 CSoutput.n342 0.573776
R14405 CSoutput.n342 CSoutput.n340 0.573776
R14406 CSoutput.n340 CSoutput.n338 0.573776
R14407 CSoutput.n334 CSoutput.n332 0.573776
R14408 CSoutput.n332 CSoutput.n330 0.573776
R14409 CSoutput.n330 CSoutput.n328 0.573776
R14410 CSoutput.n328 CSoutput.n326 0.573776
R14411 CSoutput.n323 CSoutput.n321 0.573776
R14412 CSoutput.n321 CSoutput.n319 0.573776
R14413 CSoutput.n319 CSoutput.n317 0.573776
R14414 CSoutput.n317 CSoutput.n315 0.573776
R14415 CSoutput.n349 CSoutput.n252 0.53442
R14416 CSoutput.n272 CSoutput.n270 0.358259
R14417 CSoutput.n274 CSoutput.n272 0.358259
R14418 CSoutput.n264 CSoutput.n262 0.358259
R14419 CSoutput.n266 CSoutput.n264 0.358259
R14420 CSoutput.n257 CSoutput.n255 0.358259
R14421 CSoutput.n259 CSoutput.n257 0.358259
R14422 CSoutput.n100 CSoutput.n98 0.358259
R14423 CSoutput.n98 CSoutput.n96 0.358259
R14424 CSoutput.n92 CSoutput.n90 0.358259
R14425 CSoutput.n90 CSoutput.n88 0.358259
R14426 CSoutput.n85 CSoutput.n83 0.358259
R14427 CSoutput.n83 CSoutput.n81 0.358259
R14428 CSoutput.n21 CSoutput.n20 0.169105
R14429 CSoutput.n21 CSoutput.n16 0.169105
R14430 CSoutput.n26 CSoutput.n16 0.169105
R14431 CSoutput.n27 CSoutput.n26 0.169105
R14432 CSoutput.n27 CSoutput.n14 0.169105
R14433 CSoutput.n32 CSoutput.n14 0.169105
R14434 CSoutput.n33 CSoutput.n32 0.169105
R14435 CSoutput.n34 CSoutput.n33 0.169105
R14436 CSoutput.n34 CSoutput.n12 0.169105
R14437 CSoutput.n39 CSoutput.n12 0.169105
R14438 CSoutput.n40 CSoutput.n39 0.169105
R14439 CSoutput.n40 CSoutput.n10 0.169105
R14440 CSoutput.n45 CSoutput.n10 0.169105
R14441 CSoutput.n46 CSoutput.n45 0.169105
R14442 CSoutput.n47 CSoutput.n46 0.169105
R14443 CSoutput.n47 CSoutput.n8 0.169105
R14444 CSoutput.n52 CSoutput.n8 0.169105
R14445 CSoutput.n53 CSoutput.n52 0.169105
R14446 CSoutput.n53 CSoutput.n6 0.169105
R14447 CSoutput.n58 CSoutput.n6 0.169105
R14448 CSoutput.n59 CSoutput.n58 0.169105
R14449 CSoutput.n60 CSoutput.n59 0.169105
R14450 CSoutput.n60 CSoutput.n4 0.169105
R14451 CSoutput.n66 CSoutput.n4 0.169105
R14452 CSoutput.n67 CSoutput.n66 0.169105
R14453 CSoutput.n68 CSoutput.n67 0.169105
R14454 CSoutput.n68 CSoutput.n2 0.169105
R14455 CSoutput.n73 CSoutput.n2 0.169105
R14456 CSoutput.n74 CSoutput.n73 0.169105
R14457 CSoutput.n74 CSoutput.n0 0.169105
R14458 CSoutput.n78 CSoutput.n0 0.169105
R14459 CSoutput.n195 CSoutput.n194 0.0910737
R14460 CSoutput.n246 CSoutput.n243 0.0723685
R14461 CSoutput.n200 CSoutput.n195 0.0522944
R14462 CSoutput.n243 CSoutput.n242 0.0499135
R14463 CSoutput.n194 CSoutput.n193 0.0499135
R14464 CSoutput.n228 CSoutput.n227 0.0464294
R14465 CSoutput.n236 CSoutput.n233 0.0391444
R14466 CSoutput.n195 CSoutput.t131 0.023435
R14467 CSoutput.n243 CSoutput.t130 0.02262
R14468 CSoutput.n194 CSoutput.t136 0.02262
R14469 CSoutput CSoutput.n349 0.0052
R14470 CSoutput.n165 CSoutput.n148 0.00365111
R14471 CSoutput.n168 CSoutput.n149 0.00365111
R14472 CSoutput.n151 CSoutput.n150 0.00365111
R14473 CSoutput.n193 CSoutput.n152 0.00365111
R14474 CSoutput.n157 CSoutput.n153 0.00365111
R14475 CSoutput.n240 CSoutput.n154 0.00365111
R14476 CSoutput.n231 CSoutput.n230 0.00365111
R14477 CSoutput.n211 CSoutput.n184 0.00365111
R14478 CSoutput.n213 CSoutput.n183 0.00365111
R14479 CSoutput.n201 CSoutput.n200 0.00365111
R14480 CSoutput.n207 CSoutput.n187 0.00365111
R14481 CSoutput.n209 CSoutput.n186 0.00365111
R14482 CSoutput.n131 CSoutput.n114 0.00365111
R14483 CSoutput.n134 CSoutput.n115 0.00365111
R14484 CSoutput.n117 CSoutput.n116 0.00365111
R14485 CSoutput.n227 CSoutput.n118 0.00365111
R14486 CSoutput.n123 CSoutput.n119 0.00365111
R14487 CSoutput.n250 CSoutput.n120 0.00365111
R14488 CSoutput.n162 CSoutput.n152 0.00340054
R14489 CSoutput.n155 CSoutput.n153 0.00340054
R14490 CSoutput.n240 CSoutput.n239 0.00340054
R14491 CSoutput.n235 CSoutput.n148 0.00340054
R14492 CSoutput.n164 CSoutput.n149 0.00340054
R14493 CSoutput.n167 CSoutput.n151 0.00340054
R14494 CSoutput.n206 CSoutput.n201 0.00340054
R14495 CSoutput.n208 CSoutput.n207 0.00340054
R14496 CSoutput.n210 CSoutput.n209 0.00340054
R14497 CSoutput.n232 CSoutput.n231 0.00340054
R14498 CSoutput.n212 CSoutput.n211 0.00340054
R14499 CSoutput.n214 CSoutput.n213 0.00340054
R14500 CSoutput.n128 CSoutput.n118 0.00340054
R14501 CSoutput.n121 CSoutput.n119 0.00340054
R14502 CSoutput.n250 CSoutput.n249 0.00340054
R14503 CSoutput.n245 CSoutput.n114 0.00340054
R14504 CSoutput.n130 CSoutput.n115 0.00340054
R14505 CSoutput.n133 CSoutput.n117 0.00340054
R14506 CSoutput.n163 CSoutput.n157 0.00252698
R14507 CSoutput.n156 CSoutput.n154 0.00252698
R14508 CSoutput.n238 CSoutput.n237 0.00252698
R14509 CSoutput.n166 CSoutput.n164 0.00252698
R14510 CSoutput.n169 CSoutput.n167 0.00252698
R14511 CSoutput.n242 CSoutput.n137 0.00252698
R14512 CSoutput.n163 CSoutput.n162 0.00252698
R14513 CSoutput.n156 CSoutput.n155 0.00252698
R14514 CSoutput.n239 CSoutput.n238 0.00252698
R14515 CSoutput.n166 CSoutput.n165 0.00252698
R14516 CSoutput.n169 CSoutput.n168 0.00252698
R14517 CSoutput.n150 CSoutput.n137 0.00252698
R14518 CSoutput.n217 CSoutput.n187 0.00252698
R14519 CSoutput.n216 CSoutput.n186 0.00252698
R14520 CSoutput.n215 CSoutput.n171 0.00252698
R14521 CSoutput.n212 CSoutput.n182 0.00252698
R14522 CSoutput.n219 CSoutput.n214 0.00252698
R14523 CSoutput.n228 CSoutput.n221 0.00252698
R14524 CSoutput.n217 CSoutput.n206 0.00252698
R14525 CSoutput.n216 CSoutput.n208 0.00252698
R14526 CSoutput.n215 CSoutput.n210 0.00252698
R14527 CSoutput.n230 CSoutput.n182 0.00252698
R14528 CSoutput.n219 CSoutput.n184 0.00252698
R14529 CSoutput.n221 CSoutput.n183 0.00252698
R14530 CSoutput.n129 CSoutput.n123 0.00252698
R14531 CSoutput.n122 CSoutput.n120 0.00252698
R14532 CSoutput.n248 CSoutput.n247 0.00252698
R14533 CSoutput.n132 CSoutput.n130 0.00252698
R14534 CSoutput.n135 CSoutput.n133 0.00252698
R14535 CSoutput.n252 CSoutput.n103 0.00252698
R14536 CSoutput.n129 CSoutput.n128 0.00252698
R14537 CSoutput.n122 CSoutput.n121 0.00252698
R14538 CSoutput.n249 CSoutput.n248 0.00252698
R14539 CSoutput.n132 CSoutput.n131 0.00252698
R14540 CSoutput.n135 CSoutput.n134 0.00252698
R14541 CSoutput.n116 CSoutput.n103 0.00252698
R14542 CSoutput.n237 CSoutput.n236 0.0020275
R14543 CSoutput.n236 CSoutput.n235 0.0020275
R14544 CSoutput.n233 CSoutput.n171 0.0020275
R14545 CSoutput.n233 CSoutput.n232 0.0020275
R14546 CSoutput.n247 CSoutput.n246 0.0020275
R14547 CSoutput.n246 CSoutput.n245 0.0020275
R14548 CSoutput.n147 CSoutput.n146 0.00166668
R14549 CSoutput.n229 CSoutput.n185 0.00166668
R14550 CSoutput.n113 CSoutput.n112 0.00166668
R14551 CSoutput.n251 CSoutput.n113 0.00133328
R14552 CSoutput.n185 CSoutput.n181 0.00133328
R14553 CSoutput.n241 CSoutput.n147 0.00133328
R14554 CSoutput.n244 CSoutput.n136 0.001
R14555 CSoutput.n222 CSoutput.n136 0.001
R14556 CSoutput.n124 CSoutput.n104 0.001
R14557 CSoutput.n223 CSoutput.n104 0.001
R14558 CSoutput.n125 CSoutput.n105 0.001
R14559 CSoutput.n224 CSoutput.n105 0.001
R14560 CSoutput.n126 CSoutput.n106 0.001
R14561 CSoutput.n225 CSoutput.n106 0.001
R14562 CSoutput.n127 CSoutput.n107 0.001
R14563 CSoutput.n226 CSoutput.n107 0.001
R14564 CSoutput.n220 CSoutput.n172 0.001
R14565 CSoutput.n220 CSoutput.n218 0.001
R14566 CSoutput.n202 CSoutput.n173 0.001
R14567 CSoutput.n196 CSoutput.n173 0.001
R14568 CSoutput.n203 CSoutput.n174 0.001
R14569 CSoutput.n197 CSoutput.n174 0.001
R14570 CSoutput.n204 CSoutput.n175 0.001
R14571 CSoutput.n198 CSoutput.n175 0.001
R14572 CSoutput.n205 CSoutput.n176 0.001
R14573 CSoutput.n199 CSoutput.n176 0.001
R14574 CSoutput.n234 CSoutput.n170 0.001
R14575 CSoutput.n188 CSoutput.n170 0.001
R14576 CSoutput.n158 CSoutput.n138 0.001
R14577 CSoutput.n189 CSoutput.n138 0.001
R14578 CSoutput.n159 CSoutput.n139 0.001
R14579 CSoutput.n190 CSoutput.n139 0.001
R14580 CSoutput.n160 CSoutput.n140 0.001
R14581 CSoutput.n191 CSoutput.n140 0.001
R14582 CSoutput.n161 CSoutput.n141 0.001
R14583 CSoutput.n192 CSoutput.n141 0.001
R14584 CSoutput.n192 CSoutput.n142 0.001
R14585 CSoutput.n191 CSoutput.n143 0.001
R14586 CSoutput.n190 CSoutput.n144 0.001
R14587 CSoutput.n189 CSoutput.t127 0.001
R14588 CSoutput.n188 CSoutput.n145 0.001
R14589 CSoutput.n161 CSoutput.n143 0.001
R14590 CSoutput.n160 CSoutput.n144 0.001
R14591 CSoutput.n159 CSoutput.t127 0.001
R14592 CSoutput.n158 CSoutput.n145 0.001
R14593 CSoutput.n234 CSoutput.n146 0.001
R14594 CSoutput.n199 CSoutput.n177 0.001
R14595 CSoutput.n198 CSoutput.n178 0.001
R14596 CSoutput.n197 CSoutput.n179 0.001
R14597 CSoutput.n196 CSoutput.t120 0.001
R14598 CSoutput.n218 CSoutput.n180 0.001
R14599 CSoutput.n205 CSoutput.n178 0.001
R14600 CSoutput.n204 CSoutput.n179 0.001
R14601 CSoutput.n203 CSoutput.t120 0.001
R14602 CSoutput.n202 CSoutput.n180 0.001
R14603 CSoutput.n229 CSoutput.n172 0.001
R14604 CSoutput.n226 CSoutput.n108 0.001
R14605 CSoutput.n225 CSoutput.n109 0.001
R14606 CSoutput.n224 CSoutput.n110 0.001
R14607 CSoutput.n223 CSoutput.t140 0.001
R14608 CSoutput.n222 CSoutput.n111 0.001
R14609 CSoutput.n127 CSoutput.n109 0.001
R14610 CSoutput.n126 CSoutput.n110 0.001
R14611 CSoutput.n125 CSoutput.t140 0.001
R14612 CSoutput.n124 CSoutput.n111 0.001
R14613 CSoutput.n244 CSoutput.n112 0.001
R14614 a_n5644_8799.n99 a_n5644_8799.t69 485.149
R14615 a_n5644_8799.n106 a_n5644_8799.t72 485.149
R14616 a_n5644_8799.n114 a_n5644_8799.t38 485.149
R14617 a_n5644_8799.n75 a_n5644_8799.t53 485.149
R14618 a_n5644_8799.n82 a_n5644_8799.t58 485.149
R14619 a_n5644_8799.n90 a_n5644_8799.t39 485.149
R14620 a_n5644_8799.n24 a_n5644_8799.t60 485.135
R14621 a_n5644_8799.n103 a_n5644_8799.t59 464.166
R14622 a_n5644_8799.n97 a_n5644_8799.t46 464.166
R14623 a_n5644_8799.n102 a_n5644_8799.t76 464.166
R14624 a_n5644_8799.n101 a_n5644_8799.t61 464.166
R14625 a_n5644_8799.n98 a_n5644_8799.t51 464.166
R14626 a_n5644_8799.n100 a_n5644_8799.t78 464.166
R14627 a_n5644_8799.n29 a_n5644_8799.t64 485.135
R14628 a_n5644_8799.n110 a_n5644_8799.t63 464.166
R14629 a_n5644_8799.n104 a_n5644_8799.t55 464.166
R14630 a_n5644_8799.n109 a_n5644_8799.t80 464.166
R14631 a_n5644_8799.n108 a_n5644_8799.t67 464.166
R14632 a_n5644_8799.n105 a_n5644_8799.t56 464.166
R14633 a_n5644_8799.n107 a_n5644_8799.t36 464.166
R14634 a_n5644_8799.n34 a_n5644_8799.t82 485.135
R14635 a_n5644_8799.n118 a_n5644_8799.t44 464.166
R14636 a_n5644_8799.n112 a_n5644_8799.t65 464.166
R14637 a_n5644_8799.n117 a_n5644_8799.t37 464.166
R14638 a_n5644_8799.n116 a_n5644_8799.t73 464.166
R14639 a_n5644_8799.n113 a_n5644_8799.t50 464.166
R14640 a_n5644_8799.n115 a_n5644_8799.t70 464.166
R14641 a_n5644_8799.n76 a_n5644_8799.t62 464.166
R14642 a_n5644_8799.n77 a_n5644_8799.t77 464.166
R14643 a_n5644_8799.n78 a_n5644_8799.t42 464.166
R14644 a_n5644_8799.n79 a_n5644_8799.t52 464.166
R14645 a_n5644_8799.n74 a_n5644_8799.t75 464.166
R14646 a_n5644_8799.n80 a_n5644_8799.t41 464.166
R14647 a_n5644_8799.n83 a_n5644_8799.t68 464.166
R14648 a_n5644_8799.n84 a_n5644_8799.t81 464.166
R14649 a_n5644_8799.n85 a_n5644_8799.t49 464.166
R14650 a_n5644_8799.n86 a_n5644_8799.t57 464.166
R14651 a_n5644_8799.n81 a_n5644_8799.t79 464.166
R14652 a_n5644_8799.n87 a_n5644_8799.t45 464.166
R14653 a_n5644_8799.n91 a_n5644_8799.t71 464.166
R14654 a_n5644_8799.n92 a_n5644_8799.t48 464.166
R14655 a_n5644_8799.n93 a_n5644_8799.t74 464.166
R14656 a_n5644_8799.n94 a_n5644_8799.t54 464.166
R14657 a_n5644_8799.n89 a_n5644_8799.t66 464.166
R14658 a_n5644_8799.n95 a_n5644_8799.t43 464.166
R14659 a_n5644_8799.n16 a_n5644_8799.n28 72.3034
R14660 a_n5644_8799.n28 a_n5644_8799.n98 16.6962
R14661 a_n5644_8799.n27 a_n5644_8799.n16 77.6622
R14662 a_n5644_8799.n101 a_n5644_8799.n27 5.97853
R14663 a_n5644_8799.n26 a_n5644_8799.n15 77.6622
R14664 a_n5644_8799.n15 a_n5644_8799.n25 72.3034
R14665 a_n5644_8799.n103 a_n5644_8799.n24 20.9683
R14666 a_n5644_8799.n17 a_n5644_8799.n24 70.1674
R14667 a_n5644_8799.n13 a_n5644_8799.n33 72.3034
R14668 a_n5644_8799.n33 a_n5644_8799.n105 16.6962
R14669 a_n5644_8799.n32 a_n5644_8799.n13 77.6622
R14670 a_n5644_8799.n108 a_n5644_8799.n32 5.97853
R14671 a_n5644_8799.n31 a_n5644_8799.n12 77.6622
R14672 a_n5644_8799.n12 a_n5644_8799.n30 72.3034
R14673 a_n5644_8799.n110 a_n5644_8799.n29 20.9683
R14674 a_n5644_8799.n14 a_n5644_8799.n29 70.1674
R14675 a_n5644_8799.n10 a_n5644_8799.n38 72.3034
R14676 a_n5644_8799.n38 a_n5644_8799.n113 16.6962
R14677 a_n5644_8799.n37 a_n5644_8799.n10 77.6622
R14678 a_n5644_8799.n116 a_n5644_8799.n37 5.97853
R14679 a_n5644_8799.n36 a_n5644_8799.n9 77.6622
R14680 a_n5644_8799.n9 a_n5644_8799.n35 72.3034
R14681 a_n5644_8799.n118 a_n5644_8799.n34 20.9683
R14682 a_n5644_8799.n11 a_n5644_8799.n34 70.1674
R14683 a_n5644_8799.n7 a_n5644_8799.n43 70.1674
R14684 a_n5644_8799.n80 a_n5644_8799.n43 20.9683
R14685 a_n5644_8799.n42 a_n5644_8799.n7 72.3034
R14686 a_n5644_8799.n42 a_n5644_8799.n74 16.6962
R14687 a_n5644_8799.n6 a_n5644_8799.n41 77.6622
R14688 a_n5644_8799.n79 a_n5644_8799.n41 5.97853
R14689 a_n5644_8799.n40 a_n5644_8799.n6 77.6622
R14690 a_n5644_8799.n39 a_n5644_8799.n77 16.6962
R14691 a_n5644_8799.n39 a_n5644_8799.n8 72.3034
R14692 a_n5644_8799.n4 a_n5644_8799.n48 70.1674
R14693 a_n5644_8799.n87 a_n5644_8799.n48 20.9683
R14694 a_n5644_8799.n47 a_n5644_8799.n4 72.3034
R14695 a_n5644_8799.n47 a_n5644_8799.n81 16.6962
R14696 a_n5644_8799.n3 a_n5644_8799.n46 77.6622
R14697 a_n5644_8799.n86 a_n5644_8799.n46 5.97853
R14698 a_n5644_8799.n45 a_n5644_8799.n3 77.6622
R14699 a_n5644_8799.n44 a_n5644_8799.n84 16.6962
R14700 a_n5644_8799.n44 a_n5644_8799.n5 72.3034
R14701 a_n5644_8799.n1 a_n5644_8799.n53 70.1674
R14702 a_n5644_8799.n95 a_n5644_8799.n53 20.9683
R14703 a_n5644_8799.n52 a_n5644_8799.n1 72.3034
R14704 a_n5644_8799.n52 a_n5644_8799.n89 16.6962
R14705 a_n5644_8799.n0 a_n5644_8799.n51 77.6622
R14706 a_n5644_8799.n94 a_n5644_8799.n51 5.97853
R14707 a_n5644_8799.n50 a_n5644_8799.n0 77.6622
R14708 a_n5644_8799.n49 a_n5644_8799.n92 16.6962
R14709 a_n5644_8799.n49 a_n5644_8799.n2 72.3034
R14710 a_n5644_8799.n18 a_n5644_8799.n54 98.9633
R14711 a_n5644_8799.n125 a_n5644_8799.n19 98.9632
R14712 a_n5644_8799.n19 a_n5644_8799.n124 98.6055
R14713 a_n5644_8799.n19 a_n5644_8799.n123 98.6055
R14714 a_n5644_8799.n18 a_n5644_8799.n56 98.6055
R14715 a_n5644_8799.n18 a_n5644_8799.n55 98.6055
R14716 a_n5644_8799.n59 a_n5644_8799.n57 81.4626
R14717 a_n5644_8799.n67 a_n5644_8799.n65 81.4626
R14718 a_n5644_8799.n63 a_n5644_8799.n61 81.4626
R14719 a_n5644_8799.n70 a_n5644_8799.n69 80.9324
R14720 a_n5644_8799.n72 a_n5644_8799.n71 80.9324
R14721 a_n5644_8799.n23 a_n5644_8799.n73 80.9324
R14722 a_n5644_8799.n22 a_n5644_8799.n60 80.9324
R14723 a_n5644_8799.n59 a_n5644_8799.n58 80.9324
R14724 a_n5644_8799.n67 a_n5644_8799.n66 80.9324
R14725 a_n5644_8799.n21 a_n5644_8799.n68 80.9324
R14726 a_n5644_8799.n20 a_n5644_8799.n64 80.9324
R14727 a_n5644_8799.n63 a_n5644_8799.n62 80.9324
R14728 a_n5644_8799.n16 a_n5644_8799.n99 70.4033
R14729 a_n5644_8799.n13 a_n5644_8799.n106 70.4033
R14730 a_n5644_8799.n10 a_n5644_8799.n114 70.4033
R14731 a_n5644_8799.n75 a_n5644_8799.n8 70.4033
R14732 a_n5644_8799.n82 a_n5644_8799.n5 70.4033
R14733 a_n5644_8799.n90 a_n5644_8799.n2 70.4033
R14734 a_n5644_8799.n102 a_n5644_8799.n101 48.2005
R14735 a_n5644_8799.n109 a_n5644_8799.n108 48.2005
R14736 a_n5644_8799.n117 a_n5644_8799.n116 48.2005
R14737 a_n5644_8799.n79 a_n5644_8799.n78 48.2005
R14738 a_n5644_8799.t40 a_n5644_8799.n43 485.135
R14739 a_n5644_8799.n86 a_n5644_8799.n85 48.2005
R14740 a_n5644_8799.t47 a_n5644_8799.n48 485.135
R14741 a_n5644_8799.n94 a_n5644_8799.n93 48.2005
R14742 a_n5644_8799.t83 a_n5644_8799.n53 485.135
R14743 a_n5644_8799.n25 a_n5644_8799.n97 16.6962
R14744 a_n5644_8799.n100 a_n5644_8799.n28 27.6507
R14745 a_n5644_8799.n30 a_n5644_8799.n104 16.6962
R14746 a_n5644_8799.n107 a_n5644_8799.n33 27.6507
R14747 a_n5644_8799.n35 a_n5644_8799.n112 16.6962
R14748 a_n5644_8799.n115 a_n5644_8799.n38 27.6507
R14749 a_n5644_8799.n80 a_n5644_8799.n42 27.6507
R14750 a_n5644_8799.n87 a_n5644_8799.n47 27.6507
R14751 a_n5644_8799.n95 a_n5644_8799.n52 27.6507
R14752 a_n5644_8799.n26 a_n5644_8799.n97 41.7634
R14753 a_n5644_8799.n31 a_n5644_8799.n104 41.7634
R14754 a_n5644_8799.n36 a_n5644_8799.n112 41.7634
R14755 a_n5644_8799.n77 a_n5644_8799.n40 41.7634
R14756 a_n5644_8799.n84 a_n5644_8799.n45 41.7634
R14757 a_n5644_8799.n92 a_n5644_8799.n50 41.7634
R14758 a_n5644_8799.n70 a_n5644_8799.n21 34.3237
R14759 a_n5644_8799.n100 a_n5644_8799.n99 20.9576
R14760 a_n5644_8799.n107 a_n5644_8799.n106 20.9576
R14761 a_n5644_8799.n115 a_n5644_8799.n114 20.9576
R14762 a_n5644_8799.n76 a_n5644_8799.n75 20.9576
R14763 a_n5644_8799.n83 a_n5644_8799.n82 20.9576
R14764 a_n5644_8799.n91 a_n5644_8799.n90 20.9576
R14765 a_n5644_8799.n26 a_n5644_8799.n102 5.97853
R14766 a_n5644_8799.n27 a_n5644_8799.n98 41.7634
R14767 a_n5644_8799.n31 a_n5644_8799.n109 5.97853
R14768 a_n5644_8799.n32 a_n5644_8799.n105 41.7634
R14769 a_n5644_8799.n36 a_n5644_8799.n117 5.97853
R14770 a_n5644_8799.n37 a_n5644_8799.n113 41.7634
R14771 a_n5644_8799.n78 a_n5644_8799.n40 5.97853
R14772 a_n5644_8799.n74 a_n5644_8799.n41 41.7634
R14773 a_n5644_8799.n85 a_n5644_8799.n45 5.97853
R14774 a_n5644_8799.n81 a_n5644_8799.n46 41.7634
R14775 a_n5644_8799.n93 a_n5644_8799.n50 5.97853
R14776 a_n5644_8799.n89 a_n5644_8799.n51 41.7634
R14777 a_n5644_8799.n19 a_n5644_8799.n122 31.5519
R14778 a_n5644_8799.n121 a_n5644_8799.n23 12.3339
R14779 a_n5644_8799.n122 a_n5644_8799.n121 11.4887
R14780 a_n5644_8799.n103 a_n5644_8799.n25 27.6507
R14781 a_n5644_8799.n110 a_n5644_8799.n30 27.6507
R14782 a_n5644_8799.n118 a_n5644_8799.n35 27.6507
R14783 a_n5644_8799.n39 a_n5644_8799.n76 27.6507
R14784 a_n5644_8799.n44 a_n5644_8799.n83 27.6507
R14785 a_n5644_8799.n49 a_n5644_8799.n91 27.6507
R14786 a_n5644_8799.n122 a_n5644_8799.n18 17.6132
R14787 a_n5644_8799.n111 a_n5644_8799.n17 9.05164
R14788 a_n5644_8799.n88 a_n5644_8799.n7 9.05164
R14789 a_n5644_8799.n120 a_n5644_8799.n96 6.93972
R14790 a_n5644_8799.n120 a_n5644_8799.n119 6.44309
R14791 a_n5644_8799.n111 a_n5644_8799.n14 4.94368
R14792 a_n5644_8799.n119 a_n5644_8799.n11 4.94368
R14793 a_n5644_8799.n88 a_n5644_8799.n4 4.94368
R14794 a_n5644_8799.n96 a_n5644_8799.n1 4.94368
R14795 a_n5644_8799.n119 a_n5644_8799.n111 4.10845
R14796 a_n5644_8799.n96 a_n5644_8799.n88 4.10845
R14797 a_n5644_8799.n124 a_n5644_8799.t18 3.61217
R14798 a_n5644_8799.n124 a_n5644_8799.t6 3.61217
R14799 a_n5644_8799.n123 a_n5644_8799.t14 3.61217
R14800 a_n5644_8799.n123 a_n5644_8799.t15 3.61217
R14801 a_n5644_8799.n56 a_n5644_8799.t13 3.61217
R14802 a_n5644_8799.n56 a_n5644_8799.t12 3.61217
R14803 a_n5644_8799.n55 a_n5644_8799.t23 3.61217
R14804 a_n5644_8799.n55 a_n5644_8799.t10 3.61217
R14805 a_n5644_8799.n54 a_n5644_8799.t7 3.61217
R14806 a_n5644_8799.n54 a_n5644_8799.t34 3.61217
R14807 a_n5644_8799.t2 a_n5644_8799.n125 3.61217
R14808 a_n5644_8799.n125 a_n5644_8799.t19 3.61217
R14809 a_n5644_8799.n121 a_n5644_8799.n120 3.4105
R14810 a_n5644_8799.n69 a_n5644_8799.t32 2.82907
R14811 a_n5644_8799.n69 a_n5644_8799.t25 2.82907
R14812 a_n5644_8799.n71 a_n5644_8799.t21 2.82907
R14813 a_n5644_8799.n71 a_n5644_8799.t35 2.82907
R14814 a_n5644_8799.n73 a_n5644_8799.t30 2.82907
R14815 a_n5644_8799.n73 a_n5644_8799.t4 2.82907
R14816 a_n5644_8799.n60 a_n5644_8799.t27 2.82907
R14817 a_n5644_8799.n60 a_n5644_8799.t17 2.82907
R14818 a_n5644_8799.n58 a_n5644_8799.t5 2.82907
R14819 a_n5644_8799.n58 a_n5644_8799.t3 2.82907
R14820 a_n5644_8799.n57 a_n5644_8799.t31 2.82907
R14821 a_n5644_8799.n57 a_n5644_8799.t24 2.82907
R14822 a_n5644_8799.n65 a_n5644_8799.t16 2.82907
R14823 a_n5644_8799.n65 a_n5644_8799.t8 2.82907
R14824 a_n5644_8799.n66 a_n5644_8799.t11 2.82907
R14825 a_n5644_8799.n66 a_n5644_8799.t22 2.82907
R14826 a_n5644_8799.n68 a_n5644_8799.t20 2.82907
R14827 a_n5644_8799.n68 a_n5644_8799.t1 2.82907
R14828 a_n5644_8799.n64 a_n5644_8799.t26 2.82907
R14829 a_n5644_8799.n64 a_n5644_8799.t29 2.82907
R14830 a_n5644_8799.n62 a_n5644_8799.t0 2.82907
R14831 a_n5644_8799.n62 a_n5644_8799.t28 2.82907
R14832 a_n5644_8799.n61 a_n5644_8799.t33 2.82907
R14833 a_n5644_8799.n61 a_n5644_8799.t9 2.82907
R14834 a_n5644_8799.n16 a_n5644_8799.n15 1.13686
R14835 a_n5644_8799.n13 a_n5644_8799.n12 1.13686
R14836 a_n5644_8799.n10 a_n5644_8799.n9 1.13686
R14837 a_n5644_8799.n7 a_n5644_8799.n6 1.13686
R14838 a_n5644_8799.n4 a_n5644_8799.n3 1.13686
R14839 a_n5644_8799.n1 a_n5644_8799.n0 1.13686
R14840 a_n5644_8799.n0 a_n5644_8799.n2 0.568682
R14841 a_n5644_8799.n3 a_n5644_8799.n5 0.568682
R14842 a_n5644_8799.n6 a_n5644_8799.n8 0.568682
R14843 a_n5644_8799.n9 a_n5644_8799.n11 0.568682
R14844 a_n5644_8799.n12 a_n5644_8799.n14 0.568682
R14845 a_n5644_8799.n15 a_n5644_8799.n17 0.568682
R14846 a_n5644_8799.n20 a_n5644_8799.n63 0.530672
R14847 a_n5644_8799.n21 a_n5644_8799.n67 0.530672
R14848 a_n5644_8799.n22 a_n5644_8799.n59 0.530672
R14849 a_n5644_8799.n23 a_n5644_8799.n72 0.530672
R14850 a_n5644_8799.n72 a_n5644_8799.n70 0.530672
R14851 a_n5644_8799.n23 a_n5644_8799.n22 0.530672
R14852 a_n5644_8799.n21 a_n5644_8799.n20 0.530672
R14853 vdd.n291 vdd.n255 756.745
R14854 vdd.n244 vdd.n208 756.745
R14855 vdd.n201 vdd.n165 756.745
R14856 vdd.n154 vdd.n118 756.745
R14857 vdd.n112 vdd.n76 756.745
R14858 vdd.n65 vdd.n29 756.745
R14859 vdd.n1106 vdd.n1070 756.745
R14860 vdd.n1153 vdd.n1117 756.745
R14861 vdd.n1016 vdd.n980 756.745
R14862 vdd.n1063 vdd.n1027 756.745
R14863 vdd.n927 vdd.n891 756.745
R14864 vdd.n974 vdd.n938 756.745
R14865 vdd.n1791 vdd.t61 640.208
R14866 vdd.n755 vdd.t46 640.208
R14867 vdd.n1765 vdd.t87 640.208
R14868 vdd.n747 vdd.t78 640.208
R14869 vdd.n2536 vdd.t29 640.208
R14870 vdd.n2256 vdd.t69 640.208
R14871 vdd.n622 vdd.t50 640.208
R14872 vdd.n2253 vdd.t54 640.208
R14873 vdd.n589 vdd.t58 640.208
R14874 vdd.n817 vdd.t65 640.208
R14875 vdd.n1320 vdd.t25 592.009
R14876 vdd.n1358 vdd.t72 592.009
R14877 vdd.n1254 vdd.t75 592.009
R14878 vdd.n1947 vdd.t21 592.009
R14879 vdd.n1584 vdd.t33 592.009
R14880 vdd.n1544 vdd.t40 592.009
R14881 vdd.n2908 vdd.t84 592.009
R14882 vdd.n405 vdd.t36 592.009
R14883 vdd.n365 vdd.t43 592.009
R14884 vdd.n557 vdd.t14 592.009
R14885 vdd.n2804 vdd.t18 592.009
R14886 vdd.n2711 vdd.t81 592.009
R14887 vdd.n292 vdd.n291 585
R14888 vdd.n290 vdd.n257 585
R14889 vdd.n289 vdd.n288 585
R14890 vdd.n260 vdd.n258 585
R14891 vdd.n283 vdd.n282 585
R14892 vdd.n281 vdd.n280 585
R14893 vdd.n264 vdd.n263 585
R14894 vdd.n275 vdd.n274 585
R14895 vdd.n273 vdd.n272 585
R14896 vdd.n268 vdd.n267 585
R14897 vdd.n245 vdd.n244 585
R14898 vdd.n243 vdd.n210 585
R14899 vdd.n242 vdd.n241 585
R14900 vdd.n213 vdd.n211 585
R14901 vdd.n236 vdd.n235 585
R14902 vdd.n234 vdd.n233 585
R14903 vdd.n217 vdd.n216 585
R14904 vdd.n228 vdd.n227 585
R14905 vdd.n226 vdd.n225 585
R14906 vdd.n221 vdd.n220 585
R14907 vdd.n202 vdd.n201 585
R14908 vdd.n200 vdd.n167 585
R14909 vdd.n199 vdd.n198 585
R14910 vdd.n170 vdd.n168 585
R14911 vdd.n193 vdd.n192 585
R14912 vdd.n191 vdd.n190 585
R14913 vdd.n174 vdd.n173 585
R14914 vdd.n185 vdd.n184 585
R14915 vdd.n183 vdd.n182 585
R14916 vdd.n178 vdd.n177 585
R14917 vdd.n155 vdd.n154 585
R14918 vdd.n153 vdd.n120 585
R14919 vdd.n152 vdd.n151 585
R14920 vdd.n123 vdd.n121 585
R14921 vdd.n146 vdd.n145 585
R14922 vdd.n144 vdd.n143 585
R14923 vdd.n127 vdd.n126 585
R14924 vdd.n138 vdd.n137 585
R14925 vdd.n136 vdd.n135 585
R14926 vdd.n131 vdd.n130 585
R14927 vdd.n113 vdd.n112 585
R14928 vdd.n111 vdd.n78 585
R14929 vdd.n110 vdd.n109 585
R14930 vdd.n81 vdd.n79 585
R14931 vdd.n104 vdd.n103 585
R14932 vdd.n102 vdd.n101 585
R14933 vdd.n85 vdd.n84 585
R14934 vdd.n96 vdd.n95 585
R14935 vdd.n94 vdd.n93 585
R14936 vdd.n89 vdd.n88 585
R14937 vdd.n66 vdd.n65 585
R14938 vdd.n64 vdd.n31 585
R14939 vdd.n63 vdd.n62 585
R14940 vdd.n34 vdd.n32 585
R14941 vdd.n57 vdd.n56 585
R14942 vdd.n55 vdd.n54 585
R14943 vdd.n38 vdd.n37 585
R14944 vdd.n49 vdd.n48 585
R14945 vdd.n47 vdd.n46 585
R14946 vdd.n42 vdd.n41 585
R14947 vdd.n1107 vdd.n1106 585
R14948 vdd.n1105 vdd.n1072 585
R14949 vdd.n1104 vdd.n1103 585
R14950 vdd.n1075 vdd.n1073 585
R14951 vdd.n1098 vdd.n1097 585
R14952 vdd.n1096 vdd.n1095 585
R14953 vdd.n1079 vdd.n1078 585
R14954 vdd.n1090 vdd.n1089 585
R14955 vdd.n1088 vdd.n1087 585
R14956 vdd.n1083 vdd.n1082 585
R14957 vdd.n1154 vdd.n1153 585
R14958 vdd.n1152 vdd.n1119 585
R14959 vdd.n1151 vdd.n1150 585
R14960 vdd.n1122 vdd.n1120 585
R14961 vdd.n1145 vdd.n1144 585
R14962 vdd.n1143 vdd.n1142 585
R14963 vdd.n1126 vdd.n1125 585
R14964 vdd.n1137 vdd.n1136 585
R14965 vdd.n1135 vdd.n1134 585
R14966 vdd.n1130 vdd.n1129 585
R14967 vdd.n1017 vdd.n1016 585
R14968 vdd.n1015 vdd.n982 585
R14969 vdd.n1014 vdd.n1013 585
R14970 vdd.n985 vdd.n983 585
R14971 vdd.n1008 vdd.n1007 585
R14972 vdd.n1006 vdd.n1005 585
R14973 vdd.n989 vdd.n988 585
R14974 vdd.n1000 vdd.n999 585
R14975 vdd.n998 vdd.n997 585
R14976 vdd.n993 vdd.n992 585
R14977 vdd.n1064 vdd.n1063 585
R14978 vdd.n1062 vdd.n1029 585
R14979 vdd.n1061 vdd.n1060 585
R14980 vdd.n1032 vdd.n1030 585
R14981 vdd.n1055 vdd.n1054 585
R14982 vdd.n1053 vdd.n1052 585
R14983 vdd.n1036 vdd.n1035 585
R14984 vdd.n1047 vdd.n1046 585
R14985 vdd.n1045 vdd.n1044 585
R14986 vdd.n1040 vdd.n1039 585
R14987 vdd.n928 vdd.n927 585
R14988 vdd.n926 vdd.n893 585
R14989 vdd.n925 vdd.n924 585
R14990 vdd.n896 vdd.n894 585
R14991 vdd.n919 vdd.n918 585
R14992 vdd.n917 vdd.n916 585
R14993 vdd.n900 vdd.n899 585
R14994 vdd.n911 vdd.n910 585
R14995 vdd.n909 vdd.n908 585
R14996 vdd.n904 vdd.n903 585
R14997 vdd.n975 vdd.n974 585
R14998 vdd.n973 vdd.n940 585
R14999 vdd.n972 vdd.n971 585
R15000 vdd.n943 vdd.n941 585
R15001 vdd.n966 vdd.n965 585
R15002 vdd.n964 vdd.n963 585
R15003 vdd.n947 vdd.n946 585
R15004 vdd.n958 vdd.n957 585
R15005 vdd.n956 vdd.n955 585
R15006 vdd.n951 vdd.n950 585
R15007 vdd.n3024 vdd.n330 515.122
R15008 vdd.n2906 vdd.n328 515.122
R15009 vdd.n515 vdd.n478 515.122
R15010 vdd.n2842 vdd.n479 515.122
R15011 vdd.n1942 vdd.n865 515.122
R15012 vdd.n1945 vdd.n1944 515.122
R15013 vdd.n1227 vdd.n1191 515.122
R15014 vdd.n1423 vdd.n1192 515.122
R15015 vdd.n269 vdd.t136 329.043
R15016 vdd.n222 vdd.t147 329.043
R15017 vdd.n179 vdd.t132 329.043
R15018 vdd.n132 vdd.t142 329.043
R15019 vdd.n90 vdd.t173 329.043
R15020 vdd.n43 vdd.t115 329.043
R15021 vdd.n1084 vdd.t171 329.043
R15022 vdd.n1131 vdd.t157 329.043
R15023 vdd.n994 vdd.t163 329.043
R15024 vdd.n1041 vdd.t150 329.043
R15025 vdd.n905 vdd.t113 329.043
R15026 vdd.n952 vdd.t172 329.043
R15027 vdd.n1320 vdd.t28 319.788
R15028 vdd.n1358 vdd.t74 319.788
R15029 vdd.n1254 vdd.t77 319.788
R15030 vdd.n1947 vdd.t23 319.788
R15031 vdd.n1584 vdd.t34 319.788
R15032 vdd.n1544 vdd.t41 319.788
R15033 vdd.n2908 vdd.t85 319.788
R15034 vdd.n405 vdd.t38 319.788
R15035 vdd.n365 vdd.t44 319.788
R15036 vdd.n557 vdd.t17 319.788
R15037 vdd.n2804 vdd.t20 319.788
R15038 vdd.n2711 vdd.t83 319.788
R15039 vdd.n1321 vdd.t27 303.69
R15040 vdd.n1359 vdd.t73 303.69
R15041 vdd.n1255 vdd.t76 303.69
R15042 vdd.n1948 vdd.t24 303.69
R15043 vdd.n1585 vdd.t35 303.69
R15044 vdd.n1545 vdd.t42 303.69
R15045 vdd.n2909 vdd.t86 303.69
R15046 vdd.n406 vdd.t39 303.69
R15047 vdd.n366 vdd.t45 303.69
R15048 vdd.n558 vdd.t16 303.69
R15049 vdd.n2805 vdd.t19 303.69
R15050 vdd.n2712 vdd.t82 303.69
R15051 vdd.n2479 vdd.n703 297.074
R15052 vdd.n2672 vdd.n599 297.074
R15053 vdd.n2609 vdd.n596 297.074
R15054 vdd.n2402 vdd.n704 297.074
R15055 vdd.n2217 vdd.n744 297.074
R15056 vdd.n2148 vdd.n2147 297.074
R15057 vdd.n1894 vdd.n840 297.074
R15058 vdd.n1990 vdd.n838 297.074
R15059 vdd.n2588 vdd.n597 297.074
R15060 vdd.n2675 vdd.n2674 297.074
R15061 vdd.n2251 vdd.n705 297.074
R15062 vdd.n2477 vdd.n706 297.074
R15063 vdd.n2145 vdd.n753 297.074
R15064 vdd.n751 vdd.n726 297.074
R15065 vdd.n1831 vdd.n841 297.074
R15066 vdd.n1988 vdd.n842 297.074
R15067 vdd.n2590 vdd.n597 185
R15068 vdd.n2673 vdd.n597 185
R15069 vdd.n2592 vdd.n2591 185
R15070 vdd.n2591 vdd.n595 185
R15071 vdd.n2593 vdd.n629 185
R15072 vdd.n2603 vdd.n629 185
R15073 vdd.n2594 vdd.n638 185
R15074 vdd.n638 vdd.n636 185
R15075 vdd.n2596 vdd.n2595 185
R15076 vdd.n2597 vdd.n2596 185
R15077 vdd.n2549 vdd.n637 185
R15078 vdd.n637 vdd.n633 185
R15079 vdd.n2548 vdd.n2547 185
R15080 vdd.n2547 vdd.n2546 185
R15081 vdd.n640 vdd.n639 185
R15082 vdd.n641 vdd.n640 185
R15083 vdd.n2539 vdd.n2538 185
R15084 vdd.n2540 vdd.n2539 185
R15085 vdd.n2535 vdd.n650 185
R15086 vdd.n650 vdd.n647 185
R15087 vdd.n2534 vdd.n2533 185
R15088 vdd.n2533 vdd.n2532 185
R15089 vdd.n652 vdd.n651 185
R15090 vdd.n660 vdd.n652 185
R15091 vdd.n2525 vdd.n2524 185
R15092 vdd.n2526 vdd.n2525 185
R15093 vdd.n2523 vdd.n661 185
R15094 vdd.n2374 vdd.n661 185
R15095 vdd.n2522 vdd.n2521 185
R15096 vdd.n2521 vdd.n2520 185
R15097 vdd.n663 vdd.n662 185
R15098 vdd.n664 vdd.n663 185
R15099 vdd.n2513 vdd.n2512 185
R15100 vdd.n2514 vdd.n2513 185
R15101 vdd.n2511 vdd.n673 185
R15102 vdd.n673 vdd.n670 185
R15103 vdd.n2510 vdd.n2509 185
R15104 vdd.n2509 vdd.n2508 185
R15105 vdd.n675 vdd.n674 185
R15106 vdd.n683 vdd.n675 185
R15107 vdd.n2501 vdd.n2500 185
R15108 vdd.n2502 vdd.n2501 185
R15109 vdd.n2499 vdd.n684 185
R15110 vdd.n690 vdd.n684 185
R15111 vdd.n2498 vdd.n2497 185
R15112 vdd.n2497 vdd.n2496 185
R15113 vdd.n686 vdd.n685 185
R15114 vdd.n687 vdd.n686 185
R15115 vdd.n2489 vdd.n2488 185
R15116 vdd.n2490 vdd.n2489 185
R15117 vdd.n2487 vdd.n696 185
R15118 vdd.n2395 vdd.n696 185
R15119 vdd.n2486 vdd.n2485 185
R15120 vdd.n2485 vdd.n2484 185
R15121 vdd.n698 vdd.n697 185
R15122 vdd.t3 vdd.n698 185
R15123 vdd.n2477 vdd.n2476 185
R15124 vdd.n2478 vdd.n2477 185
R15125 vdd.n2475 vdd.n706 185
R15126 vdd.n2474 vdd.n2473 185
R15127 vdd.n708 vdd.n707 185
R15128 vdd.n2260 vdd.n2259 185
R15129 vdd.n2262 vdd.n2261 185
R15130 vdd.n2264 vdd.n2263 185
R15131 vdd.n2266 vdd.n2265 185
R15132 vdd.n2268 vdd.n2267 185
R15133 vdd.n2270 vdd.n2269 185
R15134 vdd.n2272 vdd.n2271 185
R15135 vdd.n2274 vdd.n2273 185
R15136 vdd.n2276 vdd.n2275 185
R15137 vdd.n2278 vdd.n2277 185
R15138 vdd.n2280 vdd.n2279 185
R15139 vdd.n2282 vdd.n2281 185
R15140 vdd.n2284 vdd.n2283 185
R15141 vdd.n2286 vdd.n2285 185
R15142 vdd.n2288 vdd.n2287 185
R15143 vdd.n2290 vdd.n2289 185
R15144 vdd.n2292 vdd.n2291 185
R15145 vdd.n2294 vdd.n2293 185
R15146 vdd.n2296 vdd.n2295 185
R15147 vdd.n2298 vdd.n2297 185
R15148 vdd.n2300 vdd.n2299 185
R15149 vdd.n2302 vdd.n2301 185
R15150 vdd.n2304 vdd.n2303 185
R15151 vdd.n2306 vdd.n2305 185
R15152 vdd.n2308 vdd.n2307 185
R15153 vdd.n2310 vdd.n2309 185
R15154 vdd.n2312 vdd.n2311 185
R15155 vdd.n2314 vdd.n2313 185
R15156 vdd.n2316 vdd.n2315 185
R15157 vdd.n2318 vdd.n2317 185
R15158 vdd.n2320 vdd.n2319 185
R15159 vdd.n2321 vdd.n2251 185
R15160 vdd.n2471 vdd.n2251 185
R15161 vdd.n2676 vdd.n2675 185
R15162 vdd.n2677 vdd.n588 185
R15163 vdd.n2679 vdd.n2678 185
R15164 vdd.n2681 vdd.n586 185
R15165 vdd.n2683 vdd.n2682 185
R15166 vdd.n2684 vdd.n585 185
R15167 vdd.n2686 vdd.n2685 185
R15168 vdd.n2688 vdd.n583 185
R15169 vdd.n2690 vdd.n2689 185
R15170 vdd.n2691 vdd.n582 185
R15171 vdd.n2693 vdd.n2692 185
R15172 vdd.n2695 vdd.n580 185
R15173 vdd.n2697 vdd.n2696 185
R15174 vdd.n2698 vdd.n579 185
R15175 vdd.n2700 vdd.n2699 185
R15176 vdd.n2702 vdd.n578 185
R15177 vdd.n2703 vdd.n576 185
R15178 vdd.n2706 vdd.n2705 185
R15179 vdd.n577 vdd.n575 185
R15180 vdd.n2562 vdd.n2561 185
R15181 vdd.n2564 vdd.n2563 185
R15182 vdd.n2566 vdd.n2558 185
R15183 vdd.n2568 vdd.n2567 185
R15184 vdd.n2569 vdd.n2557 185
R15185 vdd.n2571 vdd.n2570 185
R15186 vdd.n2573 vdd.n2555 185
R15187 vdd.n2575 vdd.n2574 185
R15188 vdd.n2576 vdd.n2554 185
R15189 vdd.n2578 vdd.n2577 185
R15190 vdd.n2580 vdd.n2552 185
R15191 vdd.n2582 vdd.n2581 185
R15192 vdd.n2583 vdd.n2551 185
R15193 vdd.n2585 vdd.n2584 185
R15194 vdd.n2587 vdd.n2550 185
R15195 vdd.n2589 vdd.n2588 185
R15196 vdd.n2588 vdd.n484 185
R15197 vdd.n2674 vdd.n592 185
R15198 vdd.n2674 vdd.n2673 185
R15199 vdd.n2326 vdd.n594 185
R15200 vdd.n595 vdd.n594 185
R15201 vdd.n2327 vdd.n628 185
R15202 vdd.n2603 vdd.n628 185
R15203 vdd.n2329 vdd.n2328 185
R15204 vdd.n2328 vdd.n636 185
R15205 vdd.n2330 vdd.n635 185
R15206 vdd.n2597 vdd.n635 185
R15207 vdd.n2332 vdd.n2331 185
R15208 vdd.n2331 vdd.n633 185
R15209 vdd.n2333 vdd.n643 185
R15210 vdd.n2546 vdd.n643 185
R15211 vdd.n2335 vdd.n2334 185
R15212 vdd.n2334 vdd.n641 185
R15213 vdd.n2336 vdd.n649 185
R15214 vdd.n2540 vdd.n649 185
R15215 vdd.n2338 vdd.n2337 185
R15216 vdd.n2337 vdd.n647 185
R15217 vdd.n2339 vdd.n654 185
R15218 vdd.n2532 vdd.n654 185
R15219 vdd.n2341 vdd.n2340 185
R15220 vdd.n2340 vdd.n660 185
R15221 vdd.n2342 vdd.n659 185
R15222 vdd.n2526 vdd.n659 185
R15223 vdd.n2376 vdd.n2375 185
R15224 vdd.n2375 vdd.n2374 185
R15225 vdd.n2377 vdd.n666 185
R15226 vdd.n2520 vdd.n666 185
R15227 vdd.n2379 vdd.n2378 185
R15228 vdd.n2378 vdd.n664 185
R15229 vdd.n2380 vdd.n672 185
R15230 vdd.n2514 vdd.n672 185
R15231 vdd.n2382 vdd.n2381 185
R15232 vdd.n2381 vdd.n670 185
R15233 vdd.n2383 vdd.n677 185
R15234 vdd.n2508 vdd.n677 185
R15235 vdd.n2385 vdd.n2384 185
R15236 vdd.n2384 vdd.n683 185
R15237 vdd.n2386 vdd.n682 185
R15238 vdd.n2502 vdd.n682 185
R15239 vdd.n2388 vdd.n2387 185
R15240 vdd.n2387 vdd.n690 185
R15241 vdd.n2389 vdd.n689 185
R15242 vdd.n2496 vdd.n689 185
R15243 vdd.n2391 vdd.n2390 185
R15244 vdd.n2390 vdd.n687 185
R15245 vdd.n2392 vdd.n695 185
R15246 vdd.n2490 vdd.n695 185
R15247 vdd.n2394 vdd.n2393 185
R15248 vdd.n2395 vdd.n2394 185
R15249 vdd.n2325 vdd.n700 185
R15250 vdd.n2484 vdd.n700 185
R15251 vdd.n2324 vdd.n2323 185
R15252 vdd.n2323 vdd.t3 185
R15253 vdd.n2322 vdd.n705 185
R15254 vdd.n2478 vdd.n705 185
R15255 vdd.n1942 vdd.n1941 185
R15256 vdd.n1943 vdd.n1942 185
R15257 vdd.n866 vdd.n864 185
R15258 vdd.n1508 vdd.n864 185
R15259 vdd.n1511 vdd.n1510 185
R15260 vdd.n1510 vdd.n1509 185
R15261 vdd.n869 vdd.n868 185
R15262 vdd.n870 vdd.n869 185
R15263 vdd.n1497 vdd.n1496 185
R15264 vdd.n1498 vdd.n1497 185
R15265 vdd.n878 vdd.n877 185
R15266 vdd.n1489 vdd.n877 185
R15267 vdd.n1492 vdd.n1491 185
R15268 vdd.n1491 vdd.n1490 185
R15269 vdd.n881 vdd.n880 185
R15270 vdd.n888 vdd.n881 185
R15271 vdd.n1480 vdd.n1479 185
R15272 vdd.n1481 vdd.n1480 185
R15273 vdd.n890 vdd.n889 185
R15274 vdd.n889 vdd.n887 185
R15275 vdd.n1475 vdd.n1474 185
R15276 vdd.n1474 vdd.n1473 185
R15277 vdd.n1163 vdd.n1162 185
R15278 vdd.n1164 vdd.n1163 185
R15279 vdd.n1464 vdd.n1463 185
R15280 vdd.n1465 vdd.n1464 185
R15281 vdd.n1171 vdd.n1170 185
R15282 vdd.n1455 vdd.n1170 185
R15283 vdd.n1458 vdd.n1457 185
R15284 vdd.n1457 vdd.n1456 185
R15285 vdd.n1174 vdd.n1173 185
R15286 vdd.n1180 vdd.n1174 185
R15287 vdd.n1446 vdd.n1445 185
R15288 vdd.n1447 vdd.n1446 185
R15289 vdd.n1182 vdd.n1181 185
R15290 vdd.n1438 vdd.n1181 185
R15291 vdd.n1441 vdd.n1440 185
R15292 vdd.n1440 vdd.n1439 185
R15293 vdd.n1185 vdd.n1184 185
R15294 vdd.n1186 vdd.n1185 185
R15295 vdd.n1429 vdd.n1428 185
R15296 vdd.n1430 vdd.n1429 185
R15297 vdd.n1193 vdd.n1192 185
R15298 vdd.n1228 vdd.n1192 185
R15299 vdd.n1424 vdd.n1423 185
R15300 vdd.n1196 vdd.n1195 185
R15301 vdd.n1420 vdd.n1419 185
R15302 vdd.n1421 vdd.n1420 185
R15303 vdd.n1230 vdd.n1229 185
R15304 vdd.n1415 vdd.n1232 185
R15305 vdd.n1414 vdd.n1233 185
R15306 vdd.n1413 vdd.n1234 185
R15307 vdd.n1236 vdd.n1235 185
R15308 vdd.n1409 vdd.n1238 185
R15309 vdd.n1408 vdd.n1239 185
R15310 vdd.n1407 vdd.n1240 185
R15311 vdd.n1242 vdd.n1241 185
R15312 vdd.n1403 vdd.n1244 185
R15313 vdd.n1402 vdd.n1245 185
R15314 vdd.n1401 vdd.n1246 185
R15315 vdd.n1248 vdd.n1247 185
R15316 vdd.n1397 vdd.n1250 185
R15317 vdd.n1396 vdd.n1251 185
R15318 vdd.n1395 vdd.n1252 185
R15319 vdd.n1256 vdd.n1253 185
R15320 vdd.n1391 vdd.n1258 185
R15321 vdd.n1390 vdd.n1259 185
R15322 vdd.n1389 vdd.n1260 185
R15323 vdd.n1262 vdd.n1261 185
R15324 vdd.n1385 vdd.n1264 185
R15325 vdd.n1384 vdd.n1265 185
R15326 vdd.n1383 vdd.n1266 185
R15327 vdd.n1268 vdd.n1267 185
R15328 vdd.n1379 vdd.n1270 185
R15329 vdd.n1378 vdd.n1271 185
R15330 vdd.n1377 vdd.n1272 185
R15331 vdd.n1274 vdd.n1273 185
R15332 vdd.n1373 vdd.n1276 185
R15333 vdd.n1372 vdd.n1277 185
R15334 vdd.n1371 vdd.n1278 185
R15335 vdd.n1280 vdd.n1279 185
R15336 vdd.n1367 vdd.n1282 185
R15337 vdd.n1366 vdd.n1283 185
R15338 vdd.n1365 vdd.n1284 185
R15339 vdd.n1286 vdd.n1285 185
R15340 vdd.n1361 vdd.n1288 185
R15341 vdd.n1360 vdd.n1357 185
R15342 vdd.n1356 vdd.n1289 185
R15343 vdd.n1291 vdd.n1290 185
R15344 vdd.n1352 vdd.n1293 185
R15345 vdd.n1351 vdd.n1294 185
R15346 vdd.n1350 vdd.n1295 185
R15347 vdd.n1297 vdd.n1296 185
R15348 vdd.n1346 vdd.n1299 185
R15349 vdd.n1345 vdd.n1300 185
R15350 vdd.n1344 vdd.n1301 185
R15351 vdd.n1303 vdd.n1302 185
R15352 vdd.n1340 vdd.n1305 185
R15353 vdd.n1339 vdd.n1306 185
R15354 vdd.n1338 vdd.n1307 185
R15355 vdd.n1309 vdd.n1308 185
R15356 vdd.n1334 vdd.n1311 185
R15357 vdd.n1333 vdd.n1312 185
R15358 vdd.n1332 vdd.n1313 185
R15359 vdd.n1315 vdd.n1314 185
R15360 vdd.n1328 vdd.n1317 185
R15361 vdd.n1327 vdd.n1318 185
R15362 vdd.n1326 vdd.n1319 185
R15363 vdd.n1323 vdd.n1227 185
R15364 vdd.n1421 vdd.n1227 185
R15365 vdd.n1946 vdd.n1945 185
R15366 vdd.n1950 vdd.n859 185
R15367 vdd.n1613 vdd.n858 185
R15368 vdd.n1616 vdd.n1615 185
R15369 vdd.n1618 vdd.n1617 185
R15370 vdd.n1621 vdd.n1620 185
R15371 vdd.n1623 vdd.n1622 185
R15372 vdd.n1625 vdd.n1611 185
R15373 vdd.n1627 vdd.n1626 185
R15374 vdd.n1628 vdd.n1605 185
R15375 vdd.n1630 vdd.n1629 185
R15376 vdd.n1632 vdd.n1603 185
R15377 vdd.n1634 vdd.n1633 185
R15378 vdd.n1635 vdd.n1598 185
R15379 vdd.n1637 vdd.n1636 185
R15380 vdd.n1639 vdd.n1596 185
R15381 vdd.n1641 vdd.n1640 185
R15382 vdd.n1642 vdd.n1592 185
R15383 vdd.n1644 vdd.n1643 185
R15384 vdd.n1646 vdd.n1589 185
R15385 vdd.n1648 vdd.n1647 185
R15386 vdd.n1590 vdd.n1583 185
R15387 vdd.n1652 vdd.n1587 185
R15388 vdd.n1653 vdd.n1579 185
R15389 vdd.n1655 vdd.n1654 185
R15390 vdd.n1657 vdd.n1577 185
R15391 vdd.n1659 vdd.n1658 185
R15392 vdd.n1660 vdd.n1572 185
R15393 vdd.n1662 vdd.n1661 185
R15394 vdd.n1664 vdd.n1570 185
R15395 vdd.n1666 vdd.n1665 185
R15396 vdd.n1667 vdd.n1565 185
R15397 vdd.n1669 vdd.n1668 185
R15398 vdd.n1671 vdd.n1563 185
R15399 vdd.n1673 vdd.n1672 185
R15400 vdd.n1674 vdd.n1558 185
R15401 vdd.n1676 vdd.n1675 185
R15402 vdd.n1678 vdd.n1556 185
R15403 vdd.n1680 vdd.n1679 185
R15404 vdd.n1681 vdd.n1552 185
R15405 vdd.n1683 vdd.n1682 185
R15406 vdd.n1685 vdd.n1549 185
R15407 vdd.n1687 vdd.n1686 185
R15408 vdd.n1550 vdd.n1543 185
R15409 vdd.n1691 vdd.n1547 185
R15410 vdd.n1692 vdd.n1539 185
R15411 vdd.n1694 vdd.n1693 185
R15412 vdd.n1696 vdd.n1537 185
R15413 vdd.n1698 vdd.n1697 185
R15414 vdd.n1699 vdd.n1532 185
R15415 vdd.n1701 vdd.n1700 185
R15416 vdd.n1703 vdd.n1530 185
R15417 vdd.n1705 vdd.n1704 185
R15418 vdd.n1706 vdd.n1525 185
R15419 vdd.n1708 vdd.n1707 185
R15420 vdd.n1710 vdd.n1524 185
R15421 vdd.n1711 vdd.n1521 185
R15422 vdd.n1714 vdd.n1713 185
R15423 vdd.n1523 vdd.n1519 185
R15424 vdd.n1931 vdd.n1517 185
R15425 vdd.n1933 vdd.n1932 185
R15426 vdd.n1935 vdd.n1515 185
R15427 vdd.n1937 vdd.n1936 185
R15428 vdd.n1938 vdd.n865 185
R15429 vdd.n1944 vdd.n862 185
R15430 vdd.n1944 vdd.n1943 185
R15431 vdd.n873 vdd.n861 185
R15432 vdd.n1508 vdd.n861 185
R15433 vdd.n1507 vdd.n1506 185
R15434 vdd.n1509 vdd.n1507 185
R15435 vdd.n872 vdd.n871 185
R15436 vdd.n871 vdd.n870 185
R15437 vdd.n1500 vdd.n1499 185
R15438 vdd.n1499 vdd.n1498 185
R15439 vdd.n876 vdd.n875 185
R15440 vdd.n1489 vdd.n876 185
R15441 vdd.n1488 vdd.n1487 185
R15442 vdd.n1490 vdd.n1488 185
R15443 vdd.n883 vdd.n882 185
R15444 vdd.n888 vdd.n882 185
R15445 vdd.n1483 vdd.n1482 185
R15446 vdd.n1482 vdd.n1481 185
R15447 vdd.n886 vdd.n885 185
R15448 vdd.n887 vdd.n886 185
R15449 vdd.n1472 vdd.n1471 185
R15450 vdd.n1473 vdd.n1472 185
R15451 vdd.n1166 vdd.n1165 185
R15452 vdd.n1165 vdd.n1164 185
R15453 vdd.n1467 vdd.n1466 185
R15454 vdd.n1466 vdd.n1465 185
R15455 vdd.n1169 vdd.n1168 185
R15456 vdd.n1455 vdd.n1169 185
R15457 vdd.n1454 vdd.n1453 185
R15458 vdd.n1456 vdd.n1454 185
R15459 vdd.n1176 vdd.n1175 185
R15460 vdd.n1180 vdd.n1175 185
R15461 vdd.n1449 vdd.n1448 185
R15462 vdd.n1448 vdd.n1447 185
R15463 vdd.n1179 vdd.n1178 185
R15464 vdd.n1438 vdd.n1179 185
R15465 vdd.n1437 vdd.n1436 185
R15466 vdd.n1439 vdd.n1437 185
R15467 vdd.n1188 vdd.n1187 185
R15468 vdd.n1187 vdd.n1186 185
R15469 vdd.n1432 vdd.n1431 185
R15470 vdd.n1431 vdd.n1430 185
R15471 vdd.n1191 vdd.n1190 185
R15472 vdd.n1228 vdd.n1191 185
R15473 vdd.n746 vdd.n744 185
R15474 vdd.n2146 vdd.n744 185
R15475 vdd.n2068 vdd.n763 185
R15476 vdd.n763 vdd.t91 185
R15477 vdd.n2070 vdd.n2069 185
R15478 vdd.n2071 vdd.n2070 185
R15479 vdd.n2067 vdd.n762 185
R15480 vdd.n1770 vdd.n762 185
R15481 vdd.n2066 vdd.n2065 185
R15482 vdd.n2065 vdd.n2064 185
R15483 vdd.n765 vdd.n764 185
R15484 vdd.n766 vdd.n765 185
R15485 vdd.n2055 vdd.n2054 185
R15486 vdd.n2056 vdd.n2055 185
R15487 vdd.n2053 vdd.n776 185
R15488 vdd.n776 vdd.n773 185
R15489 vdd.n2052 vdd.n2051 185
R15490 vdd.n2051 vdd.n2050 185
R15491 vdd.n778 vdd.n777 185
R15492 vdd.n779 vdd.n778 185
R15493 vdd.n2043 vdd.n2042 185
R15494 vdd.n2044 vdd.n2043 185
R15495 vdd.n2041 vdd.n787 185
R15496 vdd.n792 vdd.n787 185
R15497 vdd.n2040 vdd.n2039 185
R15498 vdd.n2039 vdd.n2038 185
R15499 vdd.n789 vdd.n788 185
R15500 vdd.n798 vdd.n789 185
R15501 vdd.n2031 vdd.n2030 185
R15502 vdd.n2032 vdd.n2031 185
R15503 vdd.n2029 vdd.n799 185
R15504 vdd.n1871 vdd.n799 185
R15505 vdd.n2028 vdd.n2027 185
R15506 vdd.n2027 vdd.n2026 185
R15507 vdd.n801 vdd.n800 185
R15508 vdd.n802 vdd.n801 185
R15509 vdd.n2019 vdd.n2018 185
R15510 vdd.n2020 vdd.n2019 185
R15511 vdd.n2017 vdd.n811 185
R15512 vdd.n811 vdd.n808 185
R15513 vdd.n2016 vdd.n2015 185
R15514 vdd.n2015 vdd.n2014 185
R15515 vdd.n813 vdd.n812 185
R15516 vdd.n823 vdd.n813 185
R15517 vdd.n2006 vdd.n2005 185
R15518 vdd.n2007 vdd.n2006 185
R15519 vdd.n2004 vdd.n824 185
R15520 vdd.n824 vdd.n820 185
R15521 vdd.n2003 vdd.n2002 185
R15522 vdd.n2002 vdd.n2001 185
R15523 vdd.n826 vdd.n825 185
R15524 vdd.n827 vdd.n826 185
R15525 vdd.n1994 vdd.n1993 185
R15526 vdd.n1995 vdd.n1994 185
R15527 vdd.n1992 vdd.n836 185
R15528 vdd.n836 vdd.n833 185
R15529 vdd.n1991 vdd.n1990 185
R15530 vdd.n1990 vdd.n1989 185
R15531 vdd.n838 vdd.n837 185
R15532 vdd.n1726 vdd.n1725 185
R15533 vdd.n1727 vdd.n1723 185
R15534 vdd.n1723 vdd.n839 185
R15535 vdd.n1729 vdd.n1728 185
R15536 vdd.n1731 vdd.n1722 185
R15537 vdd.n1734 vdd.n1733 185
R15538 vdd.n1735 vdd.n1721 185
R15539 vdd.n1737 vdd.n1736 185
R15540 vdd.n1739 vdd.n1720 185
R15541 vdd.n1742 vdd.n1741 185
R15542 vdd.n1743 vdd.n1719 185
R15543 vdd.n1745 vdd.n1744 185
R15544 vdd.n1747 vdd.n1718 185
R15545 vdd.n1750 vdd.n1749 185
R15546 vdd.n1751 vdd.n1717 185
R15547 vdd.n1753 vdd.n1752 185
R15548 vdd.n1755 vdd.n1716 185
R15549 vdd.n1928 vdd.n1756 185
R15550 vdd.n1927 vdd.n1926 185
R15551 vdd.n1924 vdd.n1757 185
R15552 vdd.n1922 vdd.n1921 185
R15553 vdd.n1920 vdd.n1758 185
R15554 vdd.n1919 vdd.n1918 185
R15555 vdd.n1916 vdd.n1759 185
R15556 vdd.n1914 vdd.n1913 185
R15557 vdd.n1912 vdd.n1760 185
R15558 vdd.n1911 vdd.n1910 185
R15559 vdd.n1908 vdd.n1761 185
R15560 vdd.n1906 vdd.n1905 185
R15561 vdd.n1904 vdd.n1762 185
R15562 vdd.n1903 vdd.n1902 185
R15563 vdd.n1900 vdd.n1763 185
R15564 vdd.n1898 vdd.n1897 185
R15565 vdd.n1896 vdd.n1764 185
R15566 vdd.n1895 vdd.n1894 185
R15567 vdd.n2149 vdd.n2148 185
R15568 vdd.n2151 vdd.n2150 185
R15569 vdd.n2153 vdd.n2152 185
R15570 vdd.n2156 vdd.n2155 185
R15571 vdd.n2158 vdd.n2157 185
R15572 vdd.n2160 vdd.n2159 185
R15573 vdd.n2162 vdd.n2161 185
R15574 vdd.n2164 vdd.n2163 185
R15575 vdd.n2166 vdd.n2165 185
R15576 vdd.n2168 vdd.n2167 185
R15577 vdd.n2170 vdd.n2169 185
R15578 vdd.n2172 vdd.n2171 185
R15579 vdd.n2174 vdd.n2173 185
R15580 vdd.n2176 vdd.n2175 185
R15581 vdd.n2178 vdd.n2177 185
R15582 vdd.n2180 vdd.n2179 185
R15583 vdd.n2182 vdd.n2181 185
R15584 vdd.n2184 vdd.n2183 185
R15585 vdd.n2186 vdd.n2185 185
R15586 vdd.n2188 vdd.n2187 185
R15587 vdd.n2190 vdd.n2189 185
R15588 vdd.n2192 vdd.n2191 185
R15589 vdd.n2194 vdd.n2193 185
R15590 vdd.n2196 vdd.n2195 185
R15591 vdd.n2198 vdd.n2197 185
R15592 vdd.n2200 vdd.n2199 185
R15593 vdd.n2202 vdd.n2201 185
R15594 vdd.n2204 vdd.n2203 185
R15595 vdd.n2206 vdd.n2205 185
R15596 vdd.n2208 vdd.n2207 185
R15597 vdd.n2210 vdd.n2209 185
R15598 vdd.n2212 vdd.n2211 185
R15599 vdd.n2214 vdd.n2213 185
R15600 vdd.n2215 vdd.n745 185
R15601 vdd.n2217 vdd.n2216 185
R15602 vdd.n2218 vdd.n2217 185
R15603 vdd.n2147 vdd.n749 185
R15604 vdd.n2147 vdd.n2146 185
R15605 vdd.n1768 vdd.n750 185
R15606 vdd.t91 vdd.n750 185
R15607 vdd.n1769 vdd.n760 185
R15608 vdd.n2071 vdd.n760 185
R15609 vdd.n1772 vdd.n1771 185
R15610 vdd.n1771 vdd.n1770 185
R15611 vdd.n1773 vdd.n767 185
R15612 vdd.n2064 vdd.n767 185
R15613 vdd.n1775 vdd.n1774 185
R15614 vdd.n1774 vdd.n766 185
R15615 vdd.n1776 vdd.n774 185
R15616 vdd.n2056 vdd.n774 185
R15617 vdd.n1778 vdd.n1777 185
R15618 vdd.n1777 vdd.n773 185
R15619 vdd.n1779 vdd.n780 185
R15620 vdd.n2050 vdd.n780 185
R15621 vdd.n1781 vdd.n1780 185
R15622 vdd.n1780 vdd.n779 185
R15623 vdd.n1782 vdd.n785 185
R15624 vdd.n2044 vdd.n785 185
R15625 vdd.n1784 vdd.n1783 185
R15626 vdd.n1783 vdd.n792 185
R15627 vdd.n1785 vdd.n790 185
R15628 vdd.n2038 vdd.n790 185
R15629 vdd.n1787 vdd.n1786 185
R15630 vdd.n1786 vdd.n798 185
R15631 vdd.n1788 vdd.n796 185
R15632 vdd.n2032 vdd.n796 185
R15633 vdd.n1873 vdd.n1872 185
R15634 vdd.n1872 vdd.n1871 185
R15635 vdd.n1874 vdd.n803 185
R15636 vdd.n2026 vdd.n803 185
R15637 vdd.n1876 vdd.n1875 185
R15638 vdd.n1875 vdd.n802 185
R15639 vdd.n1877 vdd.n809 185
R15640 vdd.n2020 vdd.n809 185
R15641 vdd.n1879 vdd.n1878 185
R15642 vdd.n1878 vdd.n808 185
R15643 vdd.n1880 vdd.n814 185
R15644 vdd.n2014 vdd.n814 185
R15645 vdd.n1882 vdd.n1881 185
R15646 vdd.n1881 vdd.n823 185
R15647 vdd.n1883 vdd.n821 185
R15648 vdd.n2007 vdd.n821 185
R15649 vdd.n1885 vdd.n1884 185
R15650 vdd.n1884 vdd.n820 185
R15651 vdd.n1886 vdd.n828 185
R15652 vdd.n2001 vdd.n828 185
R15653 vdd.n1888 vdd.n1887 185
R15654 vdd.n1887 vdd.n827 185
R15655 vdd.n1889 vdd.n834 185
R15656 vdd.n1995 vdd.n834 185
R15657 vdd.n1891 vdd.n1890 185
R15658 vdd.n1890 vdd.n833 185
R15659 vdd.n1892 vdd.n840 185
R15660 vdd.n1989 vdd.n840 185
R15661 vdd.n3024 vdd.n3023 185
R15662 vdd.n3025 vdd.n3024 185
R15663 vdd.n325 vdd.n324 185
R15664 vdd.n3026 vdd.n325 185
R15665 vdd.n3029 vdd.n3028 185
R15666 vdd.n3028 vdd.n3027 185
R15667 vdd.n3030 vdd.n319 185
R15668 vdd.n319 vdd.n318 185
R15669 vdd.n3032 vdd.n3031 185
R15670 vdd.n3033 vdd.n3032 185
R15671 vdd.n314 vdd.n313 185
R15672 vdd.n3034 vdd.n314 185
R15673 vdd.n3037 vdd.n3036 185
R15674 vdd.n3036 vdd.n3035 185
R15675 vdd.n3038 vdd.n309 185
R15676 vdd.n309 vdd.n308 185
R15677 vdd.n3040 vdd.n3039 185
R15678 vdd.n3041 vdd.n3040 185
R15679 vdd.n303 vdd.n301 185
R15680 vdd.n3042 vdd.n303 185
R15681 vdd.n3045 vdd.n3044 185
R15682 vdd.n3044 vdd.n3043 185
R15683 vdd.n302 vdd.n300 185
R15684 vdd.n304 vdd.n302 185
R15685 vdd.n2881 vdd.n2880 185
R15686 vdd.n2882 vdd.n2881 185
R15687 vdd.n458 vdd.n457 185
R15688 vdd.n457 vdd.n456 185
R15689 vdd.n2876 vdd.n2875 185
R15690 vdd.n2875 vdd.n2874 185
R15691 vdd.n461 vdd.n460 185
R15692 vdd.n467 vdd.n461 185
R15693 vdd.n2865 vdd.n2864 185
R15694 vdd.n2866 vdd.n2865 185
R15695 vdd.n469 vdd.n468 185
R15696 vdd.n2857 vdd.n468 185
R15697 vdd.n2860 vdd.n2859 185
R15698 vdd.n2859 vdd.n2858 185
R15699 vdd.n472 vdd.n471 185
R15700 vdd.n473 vdd.n472 185
R15701 vdd.n2848 vdd.n2847 185
R15702 vdd.n2849 vdd.n2848 185
R15703 vdd.n480 vdd.n479 185
R15704 vdd.n516 vdd.n479 185
R15705 vdd.n2843 vdd.n2842 185
R15706 vdd.n483 vdd.n482 185
R15707 vdd.n2839 vdd.n2838 185
R15708 vdd.n2840 vdd.n2839 185
R15709 vdd.n518 vdd.n517 185
R15710 vdd.n522 vdd.n521 185
R15711 vdd.n2834 vdd.n523 185
R15712 vdd.n2833 vdd.n2832 185
R15713 vdd.n2831 vdd.n2830 185
R15714 vdd.n2829 vdd.n2828 185
R15715 vdd.n2827 vdd.n2826 185
R15716 vdd.n2825 vdd.n2824 185
R15717 vdd.n2823 vdd.n2822 185
R15718 vdd.n2821 vdd.n2820 185
R15719 vdd.n2819 vdd.n2818 185
R15720 vdd.n2817 vdd.n2816 185
R15721 vdd.n2815 vdd.n2814 185
R15722 vdd.n2813 vdd.n2812 185
R15723 vdd.n2811 vdd.n2810 185
R15724 vdd.n2809 vdd.n2808 185
R15725 vdd.n2807 vdd.n2806 185
R15726 vdd.n2798 vdd.n536 185
R15727 vdd.n2800 vdd.n2799 185
R15728 vdd.n2797 vdd.n2796 185
R15729 vdd.n2795 vdd.n2794 185
R15730 vdd.n2793 vdd.n2792 185
R15731 vdd.n2791 vdd.n2790 185
R15732 vdd.n2789 vdd.n2788 185
R15733 vdd.n2787 vdd.n2786 185
R15734 vdd.n2785 vdd.n2784 185
R15735 vdd.n2783 vdd.n2782 185
R15736 vdd.n2781 vdd.n2780 185
R15737 vdd.n2779 vdd.n2778 185
R15738 vdd.n2777 vdd.n2776 185
R15739 vdd.n2775 vdd.n2774 185
R15740 vdd.n2773 vdd.n2772 185
R15741 vdd.n2771 vdd.n2770 185
R15742 vdd.n2769 vdd.n2768 185
R15743 vdd.n2767 vdd.n2766 185
R15744 vdd.n2765 vdd.n2764 185
R15745 vdd.n2763 vdd.n2762 185
R15746 vdd.n2761 vdd.n2760 185
R15747 vdd.n2759 vdd.n2758 185
R15748 vdd.n2752 vdd.n556 185
R15749 vdd.n2754 vdd.n2753 185
R15750 vdd.n2751 vdd.n2750 185
R15751 vdd.n2749 vdd.n2748 185
R15752 vdd.n2747 vdd.n2746 185
R15753 vdd.n2745 vdd.n2744 185
R15754 vdd.n2743 vdd.n2742 185
R15755 vdd.n2741 vdd.n2740 185
R15756 vdd.n2739 vdd.n2738 185
R15757 vdd.n2737 vdd.n2736 185
R15758 vdd.n2735 vdd.n2734 185
R15759 vdd.n2733 vdd.n2732 185
R15760 vdd.n2731 vdd.n2730 185
R15761 vdd.n2729 vdd.n2728 185
R15762 vdd.n2727 vdd.n2726 185
R15763 vdd.n2725 vdd.n2724 185
R15764 vdd.n2723 vdd.n2722 185
R15765 vdd.n2721 vdd.n2720 185
R15766 vdd.n2719 vdd.n2718 185
R15767 vdd.n2717 vdd.n2716 185
R15768 vdd.n2715 vdd.n2714 185
R15769 vdd.n2710 vdd.n515 185
R15770 vdd.n2840 vdd.n515 185
R15771 vdd.n2907 vdd.n2906 185
R15772 vdd.n2911 vdd.n440 185
R15773 vdd.n2913 vdd.n2912 185
R15774 vdd.n2915 vdd.n438 185
R15775 vdd.n2917 vdd.n2916 185
R15776 vdd.n2918 vdd.n433 185
R15777 vdd.n2920 vdd.n2919 185
R15778 vdd.n2922 vdd.n431 185
R15779 vdd.n2924 vdd.n2923 185
R15780 vdd.n2925 vdd.n426 185
R15781 vdd.n2927 vdd.n2926 185
R15782 vdd.n2929 vdd.n424 185
R15783 vdd.n2931 vdd.n2930 185
R15784 vdd.n2932 vdd.n419 185
R15785 vdd.n2934 vdd.n2933 185
R15786 vdd.n2936 vdd.n417 185
R15787 vdd.n2938 vdd.n2937 185
R15788 vdd.n2939 vdd.n413 185
R15789 vdd.n2941 vdd.n2940 185
R15790 vdd.n2943 vdd.n410 185
R15791 vdd.n2945 vdd.n2944 185
R15792 vdd.n411 vdd.n404 185
R15793 vdd.n2949 vdd.n408 185
R15794 vdd.n2950 vdd.n400 185
R15795 vdd.n2952 vdd.n2951 185
R15796 vdd.n2954 vdd.n398 185
R15797 vdd.n2956 vdd.n2955 185
R15798 vdd.n2957 vdd.n393 185
R15799 vdd.n2959 vdd.n2958 185
R15800 vdd.n2961 vdd.n391 185
R15801 vdd.n2963 vdd.n2962 185
R15802 vdd.n2964 vdd.n386 185
R15803 vdd.n2966 vdd.n2965 185
R15804 vdd.n2968 vdd.n384 185
R15805 vdd.n2970 vdd.n2969 185
R15806 vdd.n2971 vdd.n379 185
R15807 vdd.n2973 vdd.n2972 185
R15808 vdd.n2975 vdd.n377 185
R15809 vdd.n2977 vdd.n2976 185
R15810 vdd.n2978 vdd.n373 185
R15811 vdd.n2980 vdd.n2979 185
R15812 vdd.n2982 vdd.n370 185
R15813 vdd.n2984 vdd.n2983 185
R15814 vdd.n371 vdd.n364 185
R15815 vdd.n2988 vdd.n368 185
R15816 vdd.n2989 vdd.n360 185
R15817 vdd.n2991 vdd.n2990 185
R15818 vdd.n2993 vdd.n358 185
R15819 vdd.n2995 vdd.n2994 185
R15820 vdd.n2996 vdd.n353 185
R15821 vdd.n2998 vdd.n2997 185
R15822 vdd.n3000 vdd.n351 185
R15823 vdd.n3002 vdd.n3001 185
R15824 vdd.n3003 vdd.n346 185
R15825 vdd.n3005 vdd.n3004 185
R15826 vdd.n3007 vdd.n344 185
R15827 vdd.n3009 vdd.n3008 185
R15828 vdd.n3010 vdd.n338 185
R15829 vdd.n3012 vdd.n3011 185
R15830 vdd.n3014 vdd.n337 185
R15831 vdd.n3015 vdd.n336 185
R15832 vdd.n3018 vdd.n3017 185
R15833 vdd.n3019 vdd.n334 185
R15834 vdd.n3020 vdd.n330 185
R15835 vdd.n2902 vdd.n328 185
R15836 vdd.n3025 vdd.n328 185
R15837 vdd.n2901 vdd.n327 185
R15838 vdd.n3026 vdd.n327 185
R15839 vdd.n2900 vdd.n326 185
R15840 vdd.n3027 vdd.n326 185
R15841 vdd.n446 vdd.n445 185
R15842 vdd.n445 vdd.n318 185
R15843 vdd.n2896 vdd.n317 185
R15844 vdd.n3033 vdd.n317 185
R15845 vdd.n2895 vdd.n316 185
R15846 vdd.n3034 vdd.n316 185
R15847 vdd.n2894 vdd.n315 185
R15848 vdd.n3035 vdd.n315 185
R15849 vdd.n449 vdd.n448 185
R15850 vdd.n448 vdd.n308 185
R15851 vdd.n2890 vdd.n307 185
R15852 vdd.n3041 vdd.n307 185
R15853 vdd.n2889 vdd.n306 185
R15854 vdd.n3042 vdd.n306 185
R15855 vdd.n2888 vdd.n305 185
R15856 vdd.n3043 vdd.n305 185
R15857 vdd.n455 vdd.n451 185
R15858 vdd.n455 vdd.n304 185
R15859 vdd.n2884 vdd.n2883 185
R15860 vdd.n2883 vdd.n2882 185
R15861 vdd.n454 vdd.n453 185
R15862 vdd.n456 vdd.n454 185
R15863 vdd.n2873 vdd.n2872 185
R15864 vdd.n2874 vdd.n2873 185
R15865 vdd.n463 vdd.n462 185
R15866 vdd.n467 vdd.n462 185
R15867 vdd.n2868 vdd.n2867 185
R15868 vdd.n2867 vdd.n2866 185
R15869 vdd.n466 vdd.n465 185
R15870 vdd.n2857 vdd.n466 185
R15871 vdd.n2856 vdd.n2855 185
R15872 vdd.n2858 vdd.n2856 185
R15873 vdd.n475 vdd.n474 185
R15874 vdd.n474 vdd.n473 185
R15875 vdd.n2851 vdd.n2850 185
R15876 vdd.n2850 vdd.n2849 185
R15877 vdd.n478 vdd.n477 185
R15878 vdd.n516 vdd.n478 185
R15879 vdd.n703 vdd.n702 185
R15880 vdd.n2469 vdd.n2468 185
R15881 vdd.n2467 vdd.n2252 185
R15882 vdd.n2471 vdd.n2252 185
R15883 vdd.n2466 vdd.n2465 185
R15884 vdd.n2464 vdd.n2463 185
R15885 vdd.n2462 vdd.n2461 185
R15886 vdd.n2460 vdd.n2459 185
R15887 vdd.n2458 vdd.n2457 185
R15888 vdd.n2456 vdd.n2455 185
R15889 vdd.n2454 vdd.n2453 185
R15890 vdd.n2452 vdd.n2451 185
R15891 vdd.n2450 vdd.n2449 185
R15892 vdd.n2448 vdd.n2447 185
R15893 vdd.n2446 vdd.n2445 185
R15894 vdd.n2444 vdd.n2443 185
R15895 vdd.n2442 vdd.n2441 185
R15896 vdd.n2440 vdd.n2439 185
R15897 vdd.n2438 vdd.n2437 185
R15898 vdd.n2436 vdd.n2435 185
R15899 vdd.n2434 vdd.n2433 185
R15900 vdd.n2432 vdd.n2431 185
R15901 vdd.n2430 vdd.n2429 185
R15902 vdd.n2428 vdd.n2427 185
R15903 vdd.n2426 vdd.n2425 185
R15904 vdd.n2424 vdd.n2423 185
R15905 vdd.n2422 vdd.n2421 185
R15906 vdd.n2420 vdd.n2419 185
R15907 vdd.n2418 vdd.n2417 185
R15908 vdd.n2416 vdd.n2415 185
R15909 vdd.n2414 vdd.n2413 185
R15910 vdd.n2412 vdd.n2411 185
R15911 vdd.n2410 vdd.n2409 185
R15912 vdd.n2407 vdd.n2406 185
R15913 vdd.n2405 vdd.n2404 185
R15914 vdd.n2403 vdd.n2402 185
R15915 vdd.n2609 vdd.n2608 185
R15916 vdd.n2611 vdd.n624 185
R15917 vdd.n2613 vdd.n2612 185
R15918 vdd.n2615 vdd.n621 185
R15919 vdd.n2617 vdd.n2616 185
R15920 vdd.n2619 vdd.n619 185
R15921 vdd.n2621 vdd.n2620 185
R15922 vdd.n2622 vdd.n618 185
R15923 vdd.n2624 vdd.n2623 185
R15924 vdd.n2626 vdd.n616 185
R15925 vdd.n2628 vdd.n2627 185
R15926 vdd.n2629 vdd.n615 185
R15927 vdd.n2631 vdd.n2630 185
R15928 vdd.n2633 vdd.n613 185
R15929 vdd.n2635 vdd.n2634 185
R15930 vdd.n2636 vdd.n612 185
R15931 vdd.n2638 vdd.n2637 185
R15932 vdd.n2640 vdd.n520 185
R15933 vdd.n2642 vdd.n2641 185
R15934 vdd.n2644 vdd.n610 185
R15935 vdd.n2646 vdd.n2645 185
R15936 vdd.n2647 vdd.n609 185
R15937 vdd.n2649 vdd.n2648 185
R15938 vdd.n2651 vdd.n607 185
R15939 vdd.n2653 vdd.n2652 185
R15940 vdd.n2654 vdd.n606 185
R15941 vdd.n2656 vdd.n2655 185
R15942 vdd.n2658 vdd.n604 185
R15943 vdd.n2660 vdd.n2659 185
R15944 vdd.n2661 vdd.n603 185
R15945 vdd.n2663 vdd.n2662 185
R15946 vdd.n2665 vdd.n602 185
R15947 vdd.n2666 vdd.n601 185
R15948 vdd.n2669 vdd.n2668 185
R15949 vdd.n2670 vdd.n599 185
R15950 vdd.n599 vdd.n484 185
R15951 vdd.n2607 vdd.n596 185
R15952 vdd.n2673 vdd.n596 185
R15953 vdd.n2606 vdd.n2605 185
R15954 vdd.n2605 vdd.n595 185
R15955 vdd.n2604 vdd.n626 185
R15956 vdd.n2604 vdd.n2603 185
R15957 vdd.n2358 vdd.n627 185
R15958 vdd.n636 vdd.n627 185
R15959 vdd.n2359 vdd.n634 185
R15960 vdd.n2597 vdd.n634 185
R15961 vdd.n2361 vdd.n2360 185
R15962 vdd.n2360 vdd.n633 185
R15963 vdd.n2362 vdd.n642 185
R15964 vdd.n2546 vdd.n642 185
R15965 vdd.n2364 vdd.n2363 185
R15966 vdd.n2363 vdd.n641 185
R15967 vdd.n2365 vdd.n648 185
R15968 vdd.n2540 vdd.n648 185
R15969 vdd.n2367 vdd.n2366 185
R15970 vdd.n2366 vdd.n647 185
R15971 vdd.n2368 vdd.n653 185
R15972 vdd.n2532 vdd.n653 185
R15973 vdd.n2370 vdd.n2369 185
R15974 vdd.n2369 vdd.n660 185
R15975 vdd.n2371 vdd.n658 185
R15976 vdd.n2526 vdd.n658 185
R15977 vdd.n2373 vdd.n2372 185
R15978 vdd.n2374 vdd.n2373 185
R15979 vdd.n2357 vdd.n665 185
R15980 vdd.n2520 vdd.n665 185
R15981 vdd.n2356 vdd.n2355 185
R15982 vdd.n2355 vdd.n664 185
R15983 vdd.n2354 vdd.n671 185
R15984 vdd.n2514 vdd.n671 185
R15985 vdd.n2353 vdd.n2352 185
R15986 vdd.n2352 vdd.n670 185
R15987 vdd.n2351 vdd.n676 185
R15988 vdd.n2508 vdd.n676 185
R15989 vdd.n2350 vdd.n2349 185
R15990 vdd.n2349 vdd.n683 185
R15991 vdd.n2348 vdd.n681 185
R15992 vdd.n2502 vdd.n681 185
R15993 vdd.n2347 vdd.n2346 185
R15994 vdd.n2346 vdd.n690 185
R15995 vdd.n2345 vdd.n688 185
R15996 vdd.n2496 vdd.n688 185
R15997 vdd.n2344 vdd.n2343 185
R15998 vdd.n2343 vdd.n687 185
R15999 vdd.n2255 vdd.n694 185
R16000 vdd.n2490 vdd.n694 185
R16001 vdd.n2397 vdd.n2396 185
R16002 vdd.n2396 vdd.n2395 185
R16003 vdd.n2398 vdd.n699 185
R16004 vdd.n2484 vdd.n699 185
R16005 vdd.n2400 vdd.n2399 185
R16006 vdd.n2399 vdd.t3 185
R16007 vdd.n2401 vdd.n704 185
R16008 vdd.n2478 vdd.n704 185
R16009 vdd.n2480 vdd.n2479 185
R16010 vdd.n2479 vdd.n2478 185
R16011 vdd.n2481 vdd.n701 185
R16012 vdd.n701 vdd.t3 185
R16013 vdd.n2483 vdd.n2482 185
R16014 vdd.n2484 vdd.n2483 185
R16015 vdd.n693 vdd.n692 185
R16016 vdd.n2395 vdd.n693 185
R16017 vdd.n2492 vdd.n2491 185
R16018 vdd.n2491 vdd.n2490 185
R16019 vdd.n2493 vdd.n691 185
R16020 vdd.n691 vdd.n687 185
R16021 vdd.n2495 vdd.n2494 185
R16022 vdd.n2496 vdd.n2495 185
R16023 vdd.n680 vdd.n679 185
R16024 vdd.n690 vdd.n680 185
R16025 vdd.n2504 vdd.n2503 185
R16026 vdd.n2503 vdd.n2502 185
R16027 vdd.n2505 vdd.n678 185
R16028 vdd.n683 vdd.n678 185
R16029 vdd.n2507 vdd.n2506 185
R16030 vdd.n2508 vdd.n2507 185
R16031 vdd.n669 vdd.n668 185
R16032 vdd.n670 vdd.n669 185
R16033 vdd.n2516 vdd.n2515 185
R16034 vdd.n2515 vdd.n2514 185
R16035 vdd.n2517 vdd.n667 185
R16036 vdd.n667 vdd.n664 185
R16037 vdd.n2519 vdd.n2518 185
R16038 vdd.n2520 vdd.n2519 185
R16039 vdd.n657 vdd.n656 185
R16040 vdd.n2374 vdd.n657 185
R16041 vdd.n2528 vdd.n2527 185
R16042 vdd.n2527 vdd.n2526 185
R16043 vdd.n2529 vdd.n655 185
R16044 vdd.n660 vdd.n655 185
R16045 vdd.n2531 vdd.n2530 185
R16046 vdd.n2532 vdd.n2531 185
R16047 vdd.n646 vdd.n645 185
R16048 vdd.n647 vdd.n646 185
R16049 vdd.n2542 vdd.n2541 185
R16050 vdd.n2541 vdd.n2540 185
R16051 vdd.n2543 vdd.n644 185
R16052 vdd.n644 vdd.n641 185
R16053 vdd.n2545 vdd.n2544 185
R16054 vdd.n2546 vdd.n2545 185
R16055 vdd.n632 vdd.n631 185
R16056 vdd.n633 vdd.n632 185
R16057 vdd.n2599 vdd.n2598 185
R16058 vdd.n2598 vdd.n2597 185
R16059 vdd.n2600 vdd.n630 185
R16060 vdd.n636 vdd.n630 185
R16061 vdd.n2602 vdd.n2601 185
R16062 vdd.n2603 vdd.n2602 185
R16063 vdd.n600 vdd.n598 185
R16064 vdd.n598 vdd.n595 185
R16065 vdd.n2672 vdd.n2671 185
R16066 vdd.n2673 vdd.n2672 185
R16067 vdd.n2145 vdd.n2144 185
R16068 vdd.n2146 vdd.n2145 185
R16069 vdd.n754 vdd.n752 185
R16070 vdd.n752 vdd.t91 185
R16071 vdd.n2060 vdd.n761 185
R16072 vdd.n2071 vdd.n761 185
R16073 vdd.n2061 vdd.n770 185
R16074 vdd.n1770 vdd.n770 185
R16075 vdd.n2063 vdd.n2062 185
R16076 vdd.n2064 vdd.n2063 185
R16077 vdd.n2059 vdd.n769 185
R16078 vdd.n769 vdd.n766 185
R16079 vdd.n2058 vdd.n2057 185
R16080 vdd.n2057 vdd.n2056 185
R16081 vdd.n772 vdd.n771 185
R16082 vdd.n773 vdd.n772 185
R16083 vdd.n2049 vdd.n2048 185
R16084 vdd.n2050 vdd.n2049 185
R16085 vdd.n2047 vdd.n782 185
R16086 vdd.n782 vdd.n779 185
R16087 vdd.n2046 vdd.n2045 185
R16088 vdd.n2045 vdd.n2044 185
R16089 vdd.n784 vdd.n783 185
R16090 vdd.n792 vdd.n784 185
R16091 vdd.n2037 vdd.n2036 185
R16092 vdd.n2038 vdd.n2037 185
R16093 vdd.n2035 vdd.n793 185
R16094 vdd.n798 vdd.n793 185
R16095 vdd.n2034 vdd.n2033 185
R16096 vdd.n2033 vdd.n2032 185
R16097 vdd.n795 vdd.n794 185
R16098 vdd.n1871 vdd.n795 185
R16099 vdd.n2025 vdd.n2024 185
R16100 vdd.n2026 vdd.n2025 185
R16101 vdd.n2023 vdd.n805 185
R16102 vdd.n805 vdd.n802 185
R16103 vdd.n2022 vdd.n2021 185
R16104 vdd.n2021 vdd.n2020 185
R16105 vdd.n807 vdd.n806 185
R16106 vdd.n808 vdd.n807 185
R16107 vdd.n2013 vdd.n2012 185
R16108 vdd.n2014 vdd.n2013 185
R16109 vdd.n2010 vdd.n816 185
R16110 vdd.n823 vdd.n816 185
R16111 vdd.n2009 vdd.n2008 185
R16112 vdd.n2008 vdd.n2007 185
R16113 vdd.n819 vdd.n818 185
R16114 vdd.n820 vdd.n819 185
R16115 vdd.n2000 vdd.n1999 185
R16116 vdd.n2001 vdd.n2000 185
R16117 vdd.n1998 vdd.n830 185
R16118 vdd.n830 vdd.n827 185
R16119 vdd.n1997 vdd.n1996 185
R16120 vdd.n1996 vdd.n1995 185
R16121 vdd.n832 vdd.n831 185
R16122 vdd.n833 vdd.n832 185
R16123 vdd.n1988 vdd.n1987 185
R16124 vdd.n1989 vdd.n1988 185
R16125 vdd.n2076 vdd.n726 185
R16126 vdd.n2218 vdd.n726 185
R16127 vdd.n2078 vdd.n2077 185
R16128 vdd.n2080 vdd.n2079 185
R16129 vdd.n2082 vdd.n2081 185
R16130 vdd.n2084 vdd.n2083 185
R16131 vdd.n2086 vdd.n2085 185
R16132 vdd.n2088 vdd.n2087 185
R16133 vdd.n2090 vdd.n2089 185
R16134 vdd.n2092 vdd.n2091 185
R16135 vdd.n2094 vdd.n2093 185
R16136 vdd.n2096 vdd.n2095 185
R16137 vdd.n2098 vdd.n2097 185
R16138 vdd.n2100 vdd.n2099 185
R16139 vdd.n2102 vdd.n2101 185
R16140 vdd.n2104 vdd.n2103 185
R16141 vdd.n2106 vdd.n2105 185
R16142 vdd.n2108 vdd.n2107 185
R16143 vdd.n2110 vdd.n2109 185
R16144 vdd.n2112 vdd.n2111 185
R16145 vdd.n2114 vdd.n2113 185
R16146 vdd.n2116 vdd.n2115 185
R16147 vdd.n2118 vdd.n2117 185
R16148 vdd.n2120 vdd.n2119 185
R16149 vdd.n2122 vdd.n2121 185
R16150 vdd.n2124 vdd.n2123 185
R16151 vdd.n2126 vdd.n2125 185
R16152 vdd.n2128 vdd.n2127 185
R16153 vdd.n2130 vdd.n2129 185
R16154 vdd.n2132 vdd.n2131 185
R16155 vdd.n2134 vdd.n2133 185
R16156 vdd.n2136 vdd.n2135 185
R16157 vdd.n2138 vdd.n2137 185
R16158 vdd.n2140 vdd.n2139 185
R16159 vdd.n2142 vdd.n2141 185
R16160 vdd.n2143 vdd.n753 185
R16161 vdd.n2075 vdd.n751 185
R16162 vdd.n2146 vdd.n751 185
R16163 vdd.n2074 vdd.n2073 185
R16164 vdd.n2073 vdd.t91 185
R16165 vdd.n2072 vdd.n758 185
R16166 vdd.n2072 vdd.n2071 185
R16167 vdd.n1852 vdd.n759 185
R16168 vdd.n1770 vdd.n759 185
R16169 vdd.n1853 vdd.n768 185
R16170 vdd.n2064 vdd.n768 185
R16171 vdd.n1855 vdd.n1854 185
R16172 vdd.n1854 vdd.n766 185
R16173 vdd.n1856 vdd.n775 185
R16174 vdd.n2056 vdd.n775 185
R16175 vdd.n1858 vdd.n1857 185
R16176 vdd.n1857 vdd.n773 185
R16177 vdd.n1859 vdd.n781 185
R16178 vdd.n2050 vdd.n781 185
R16179 vdd.n1861 vdd.n1860 185
R16180 vdd.n1860 vdd.n779 185
R16181 vdd.n1862 vdd.n786 185
R16182 vdd.n2044 vdd.n786 185
R16183 vdd.n1864 vdd.n1863 185
R16184 vdd.n1863 vdd.n792 185
R16185 vdd.n1865 vdd.n791 185
R16186 vdd.n2038 vdd.n791 185
R16187 vdd.n1867 vdd.n1866 185
R16188 vdd.n1866 vdd.n798 185
R16189 vdd.n1868 vdd.n797 185
R16190 vdd.n2032 vdd.n797 185
R16191 vdd.n1870 vdd.n1869 185
R16192 vdd.n1871 vdd.n1870 185
R16193 vdd.n1851 vdd.n804 185
R16194 vdd.n2026 vdd.n804 185
R16195 vdd.n1850 vdd.n1849 185
R16196 vdd.n1849 vdd.n802 185
R16197 vdd.n1848 vdd.n810 185
R16198 vdd.n2020 vdd.n810 185
R16199 vdd.n1847 vdd.n1846 185
R16200 vdd.n1846 vdd.n808 185
R16201 vdd.n1845 vdd.n815 185
R16202 vdd.n2014 vdd.n815 185
R16203 vdd.n1844 vdd.n1843 185
R16204 vdd.n1843 vdd.n823 185
R16205 vdd.n1842 vdd.n822 185
R16206 vdd.n2007 vdd.n822 185
R16207 vdd.n1841 vdd.n1840 185
R16208 vdd.n1840 vdd.n820 185
R16209 vdd.n1839 vdd.n829 185
R16210 vdd.n2001 vdd.n829 185
R16211 vdd.n1838 vdd.n1837 185
R16212 vdd.n1837 vdd.n827 185
R16213 vdd.n1836 vdd.n835 185
R16214 vdd.n1995 vdd.n835 185
R16215 vdd.n1835 vdd.n1834 185
R16216 vdd.n1834 vdd.n833 185
R16217 vdd.n1833 vdd.n841 185
R16218 vdd.n1989 vdd.n841 185
R16219 vdd.n1986 vdd.n842 185
R16220 vdd.n1985 vdd.n1984 185
R16221 vdd.n1982 vdd.n843 185
R16222 vdd.n1980 vdd.n1979 185
R16223 vdd.n1978 vdd.n844 185
R16224 vdd.n1977 vdd.n1976 185
R16225 vdd.n1974 vdd.n845 185
R16226 vdd.n1972 vdd.n1971 185
R16227 vdd.n1970 vdd.n846 185
R16228 vdd.n1969 vdd.n1968 185
R16229 vdd.n1966 vdd.n847 185
R16230 vdd.n1964 vdd.n1963 185
R16231 vdd.n1962 vdd.n848 185
R16232 vdd.n1961 vdd.n1960 185
R16233 vdd.n1958 vdd.n849 185
R16234 vdd.n1956 vdd.n1955 185
R16235 vdd.n1954 vdd.n850 185
R16236 vdd.n1953 vdd.n852 185
R16237 vdd.n1798 vdd.n853 185
R16238 vdd.n1801 vdd.n1800 185
R16239 vdd.n1803 vdd.n1802 185
R16240 vdd.n1805 vdd.n1797 185
R16241 vdd.n1808 vdd.n1807 185
R16242 vdd.n1809 vdd.n1796 185
R16243 vdd.n1811 vdd.n1810 185
R16244 vdd.n1813 vdd.n1795 185
R16245 vdd.n1816 vdd.n1815 185
R16246 vdd.n1817 vdd.n1794 185
R16247 vdd.n1819 vdd.n1818 185
R16248 vdd.n1821 vdd.n1793 185
R16249 vdd.n1824 vdd.n1823 185
R16250 vdd.n1825 vdd.n1790 185
R16251 vdd.n1828 vdd.n1827 185
R16252 vdd.n1830 vdd.n1789 185
R16253 vdd.n1832 vdd.n1831 185
R16254 vdd.n1831 vdd.n839 185
R16255 vdd.n291 vdd.n290 171.744
R16256 vdd.n290 vdd.n289 171.744
R16257 vdd.n289 vdd.n258 171.744
R16258 vdd.n282 vdd.n258 171.744
R16259 vdd.n282 vdd.n281 171.744
R16260 vdd.n281 vdd.n263 171.744
R16261 vdd.n274 vdd.n263 171.744
R16262 vdd.n274 vdd.n273 171.744
R16263 vdd.n273 vdd.n267 171.744
R16264 vdd.n244 vdd.n243 171.744
R16265 vdd.n243 vdd.n242 171.744
R16266 vdd.n242 vdd.n211 171.744
R16267 vdd.n235 vdd.n211 171.744
R16268 vdd.n235 vdd.n234 171.744
R16269 vdd.n234 vdd.n216 171.744
R16270 vdd.n227 vdd.n216 171.744
R16271 vdd.n227 vdd.n226 171.744
R16272 vdd.n226 vdd.n220 171.744
R16273 vdd.n201 vdd.n200 171.744
R16274 vdd.n200 vdd.n199 171.744
R16275 vdd.n199 vdd.n168 171.744
R16276 vdd.n192 vdd.n168 171.744
R16277 vdd.n192 vdd.n191 171.744
R16278 vdd.n191 vdd.n173 171.744
R16279 vdd.n184 vdd.n173 171.744
R16280 vdd.n184 vdd.n183 171.744
R16281 vdd.n183 vdd.n177 171.744
R16282 vdd.n154 vdd.n153 171.744
R16283 vdd.n153 vdd.n152 171.744
R16284 vdd.n152 vdd.n121 171.744
R16285 vdd.n145 vdd.n121 171.744
R16286 vdd.n145 vdd.n144 171.744
R16287 vdd.n144 vdd.n126 171.744
R16288 vdd.n137 vdd.n126 171.744
R16289 vdd.n137 vdd.n136 171.744
R16290 vdd.n136 vdd.n130 171.744
R16291 vdd.n112 vdd.n111 171.744
R16292 vdd.n111 vdd.n110 171.744
R16293 vdd.n110 vdd.n79 171.744
R16294 vdd.n103 vdd.n79 171.744
R16295 vdd.n103 vdd.n102 171.744
R16296 vdd.n102 vdd.n84 171.744
R16297 vdd.n95 vdd.n84 171.744
R16298 vdd.n95 vdd.n94 171.744
R16299 vdd.n94 vdd.n88 171.744
R16300 vdd.n65 vdd.n64 171.744
R16301 vdd.n64 vdd.n63 171.744
R16302 vdd.n63 vdd.n32 171.744
R16303 vdd.n56 vdd.n32 171.744
R16304 vdd.n56 vdd.n55 171.744
R16305 vdd.n55 vdd.n37 171.744
R16306 vdd.n48 vdd.n37 171.744
R16307 vdd.n48 vdd.n47 171.744
R16308 vdd.n47 vdd.n41 171.744
R16309 vdd.n1106 vdd.n1105 171.744
R16310 vdd.n1105 vdd.n1104 171.744
R16311 vdd.n1104 vdd.n1073 171.744
R16312 vdd.n1097 vdd.n1073 171.744
R16313 vdd.n1097 vdd.n1096 171.744
R16314 vdd.n1096 vdd.n1078 171.744
R16315 vdd.n1089 vdd.n1078 171.744
R16316 vdd.n1089 vdd.n1088 171.744
R16317 vdd.n1088 vdd.n1082 171.744
R16318 vdd.n1153 vdd.n1152 171.744
R16319 vdd.n1152 vdd.n1151 171.744
R16320 vdd.n1151 vdd.n1120 171.744
R16321 vdd.n1144 vdd.n1120 171.744
R16322 vdd.n1144 vdd.n1143 171.744
R16323 vdd.n1143 vdd.n1125 171.744
R16324 vdd.n1136 vdd.n1125 171.744
R16325 vdd.n1136 vdd.n1135 171.744
R16326 vdd.n1135 vdd.n1129 171.744
R16327 vdd.n1016 vdd.n1015 171.744
R16328 vdd.n1015 vdd.n1014 171.744
R16329 vdd.n1014 vdd.n983 171.744
R16330 vdd.n1007 vdd.n983 171.744
R16331 vdd.n1007 vdd.n1006 171.744
R16332 vdd.n1006 vdd.n988 171.744
R16333 vdd.n999 vdd.n988 171.744
R16334 vdd.n999 vdd.n998 171.744
R16335 vdd.n998 vdd.n992 171.744
R16336 vdd.n1063 vdd.n1062 171.744
R16337 vdd.n1062 vdd.n1061 171.744
R16338 vdd.n1061 vdd.n1030 171.744
R16339 vdd.n1054 vdd.n1030 171.744
R16340 vdd.n1054 vdd.n1053 171.744
R16341 vdd.n1053 vdd.n1035 171.744
R16342 vdd.n1046 vdd.n1035 171.744
R16343 vdd.n1046 vdd.n1045 171.744
R16344 vdd.n1045 vdd.n1039 171.744
R16345 vdd.n927 vdd.n926 171.744
R16346 vdd.n926 vdd.n925 171.744
R16347 vdd.n925 vdd.n894 171.744
R16348 vdd.n918 vdd.n894 171.744
R16349 vdd.n918 vdd.n917 171.744
R16350 vdd.n917 vdd.n899 171.744
R16351 vdd.n910 vdd.n899 171.744
R16352 vdd.n910 vdd.n909 171.744
R16353 vdd.n909 vdd.n903 171.744
R16354 vdd.n974 vdd.n973 171.744
R16355 vdd.n973 vdd.n972 171.744
R16356 vdd.n972 vdd.n941 171.744
R16357 vdd.n965 vdd.n941 171.744
R16358 vdd.n965 vdd.n964 171.744
R16359 vdd.n964 vdd.n946 171.744
R16360 vdd.n957 vdd.n946 171.744
R16361 vdd.n957 vdd.n956 171.744
R16362 vdd.n956 vdd.n950 171.744
R16363 vdd.n3017 vdd.n334 146.341
R16364 vdd.n3015 vdd.n3014 146.341
R16365 vdd.n3012 vdd.n338 146.341
R16366 vdd.n3008 vdd.n3007 146.341
R16367 vdd.n3005 vdd.n346 146.341
R16368 vdd.n3001 vdd.n3000 146.341
R16369 vdd.n2998 vdd.n353 146.341
R16370 vdd.n2994 vdd.n2993 146.341
R16371 vdd.n2991 vdd.n360 146.341
R16372 vdd.n371 vdd.n368 146.341
R16373 vdd.n2983 vdd.n2982 146.341
R16374 vdd.n2980 vdd.n373 146.341
R16375 vdd.n2976 vdd.n2975 146.341
R16376 vdd.n2973 vdd.n379 146.341
R16377 vdd.n2969 vdd.n2968 146.341
R16378 vdd.n2966 vdd.n386 146.341
R16379 vdd.n2962 vdd.n2961 146.341
R16380 vdd.n2959 vdd.n393 146.341
R16381 vdd.n2955 vdd.n2954 146.341
R16382 vdd.n2952 vdd.n400 146.341
R16383 vdd.n411 vdd.n408 146.341
R16384 vdd.n2944 vdd.n2943 146.341
R16385 vdd.n2941 vdd.n413 146.341
R16386 vdd.n2937 vdd.n2936 146.341
R16387 vdd.n2934 vdd.n419 146.341
R16388 vdd.n2930 vdd.n2929 146.341
R16389 vdd.n2927 vdd.n426 146.341
R16390 vdd.n2923 vdd.n2922 146.341
R16391 vdd.n2920 vdd.n433 146.341
R16392 vdd.n2916 vdd.n2915 146.341
R16393 vdd.n2913 vdd.n440 146.341
R16394 vdd.n2850 vdd.n478 146.341
R16395 vdd.n2850 vdd.n474 146.341
R16396 vdd.n2856 vdd.n474 146.341
R16397 vdd.n2856 vdd.n466 146.341
R16398 vdd.n2867 vdd.n466 146.341
R16399 vdd.n2867 vdd.n462 146.341
R16400 vdd.n2873 vdd.n462 146.341
R16401 vdd.n2873 vdd.n454 146.341
R16402 vdd.n2883 vdd.n454 146.341
R16403 vdd.n2883 vdd.n455 146.341
R16404 vdd.n455 vdd.n305 146.341
R16405 vdd.n306 vdd.n305 146.341
R16406 vdd.n307 vdd.n306 146.341
R16407 vdd.n448 vdd.n307 146.341
R16408 vdd.n448 vdd.n315 146.341
R16409 vdd.n316 vdd.n315 146.341
R16410 vdd.n317 vdd.n316 146.341
R16411 vdd.n445 vdd.n317 146.341
R16412 vdd.n445 vdd.n326 146.341
R16413 vdd.n327 vdd.n326 146.341
R16414 vdd.n328 vdd.n327 146.341
R16415 vdd.n2839 vdd.n483 146.341
R16416 vdd.n2839 vdd.n517 146.341
R16417 vdd.n523 vdd.n522 146.341
R16418 vdd.n2832 vdd.n2831 146.341
R16419 vdd.n2828 vdd.n2827 146.341
R16420 vdd.n2824 vdd.n2823 146.341
R16421 vdd.n2820 vdd.n2819 146.341
R16422 vdd.n2816 vdd.n2815 146.341
R16423 vdd.n2812 vdd.n2811 146.341
R16424 vdd.n2808 vdd.n2807 146.341
R16425 vdd.n2799 vdd.n2798 146.341
R16426 vdd.n2796 vdd.n2795 146.341
R16427 vdd.n2792 vdd.n2791 146.341
R16428 vdd.n2788 vdd.n2787 146.341
R16429 vdd.n2784 vdd.n2783 146.341
R16430 vdd.n2780 vdd.n2779 146.341
R16431 vdd.n2776 vdd.n2775 146.341
R16432 vdd.n2772 vdd.n2771 146.341
R16433 vdd.n2768 vdd.n2767 146.341
R16434 vdd.n2764 vdd.n2763 146.341
R16435 vdd.n2760 vdd.n2759 146.341
R16436 vdd.n2753 vdd.n2752 146.341
R16437 vdd.n2750 vdd.n2749 146.341
R16438 vdd.n2746 vdd.n2745 146.341
R16439 vdd.n2742 vdd.n2741 146.341
R16440 vdd.n2738 vdd.n2737 146.341
R16441 vdd.n2734 vdd.n2733 146.341
R16442 vdd.n2730 vdd.n2729 146.341
R16443 vdd.n2726 vdd.n2725 146.341
R16444 vdd.n2722 vdd.n2721 146.341
R16445 vdd.n2718 vdd.n2717 146.341
R16446 vdd.n2714 vdd.n515 146.341
R16447 vdd.n2848 vdd.n479 146.341
R16448 vdd.n2848 vdd.n472 146.341
R16449 vdd.n2859 vdd.n472 146.341
R16450 vdd.n2859 vdd.n468 146.341
R16451 vdd.n2865 vdd.n468 146.341
R16452 vdd.n2865 vdd.n461 146.341
R16453 vdd.n2875 vdd.n461 146.341
R16454 vdd.n2875 vdd.n457 146.341
R16455 vdd.n2881 vdd.n457 146.341
R16456 vdd.n2881 vdd.n302 146.341
R16457 vdd.n3044 vdd.n302 146.341
R16458 vdd.n3044 vdd.n303 146.341
R16459 vdd.n3040 vdd.n303 146.341
R16460 vdd.n3040 vdd.n309 146.341
R16461 vdd.n3036 vdd.n309 146.341
R16462 vdd.n3036 vdd.n314 146.341
R16463 vdd.n3032 vdd.n314 146.341
R16464 vdd.n3032 vdd.n319 146.341
R16465 vdd.n3028 vdd.n319 146.341
R16466 vdd.n3028 vdd.n325 146.341
R16467 vdd.n3024 vdd.n325 146.341
R16468 vdd.n1936 vdd.n1935 146.341
R16469 vdd.n1933 vdd.n1517 146.341
R16470 vdd.n1713 vdd.n1523 146.341
R16471 vdd.n1711 vdd.n1710 146.341
R16472 vdd.n1708 vdd.n1525 146.341
R16473 vdd.n1704 vdd.n1703 146.341
R16474 vdd.n1701 vdd.n1532 146.341
R16475 vdd.n1697 vdd.n1696 146.341
R16476 vdd.n1694 vdd.n1539 146.341
R16477 vdd.n1550 vdd.n1547 146.341
R16478 vdd.n1686 vdd.n1685 146.341
R16479 vdd.n1683 vdd.n1552 146.341
R16480 vdd.n1679 vdd.n1678 146.341
R16481 vdd.n1676 vdd.n1558 146.341
R16482 vdd.n1672 vdd.n1671 146.341
R16483 vdd.n1669 vdd.n1565 146.341
R16484 vdd.n1665 vdd.n1664 146.341
R16485 vdd.n1662 vdd.n1572 146.341
R16486 vdd.n1658 vdd.n1657 146.341
R16487 vdd.n1655 vdd.n1579 146.341
R16488 vdd.n1590 vdd.n1587 146.341
R16489 vdd.n1647 vdd.n1646 146.341
R16490 vdd.n1644 vdd.n1592 146.341
R16491 vdd.n1640 vdd.n1639 146.341
R16492 vdd.n1637 vdd.n1598 146.341
R16493 vdd.n1633 vdd.n1632 146.341
R16494 vdd.n1630 vdd.n1605 146.341
R16495 vdd.n1626 vdd.n1625 146.341
R16496 vdd.n1623 vdd.n1620 146.341
R16497 vdd.n1618 vdd.n1615 146.341
R16498 vdd.n1613 vdd.n859 146.341
R16499 vdd.n1431 vdd.n1191 146.341
R16500 vdd.n1431 vdd.n1187 146.341
R16501 vdd.n1437 vdd.n1187 146.341
R16502 vdd.n1437 vdd.n1179 146.341
R16503 vdd.n1448 vdd.n1179 146.341
R16504 vdd.n1448 vdd.n1175 146.341
R16505 vdd.n1454 vdd.n1175 146.341
R16506 vdd.n1454 vdd.n1169 146.341
R16507 vdd.n1466 vdd.n1169 146.341
R16508 vdd.n1466 vdd.n1165 146.341
R16509 vdd.n1472 vdd.n1165 146.341
R16510 vdd.n1472 vdd.n886 146.341
R16511 vdd.n1482 vdd.n886 146.341
R16512 vdd.n1482 vdd.n882 146.341
R16513 vdd.n1488 vdd.n882 146.341
R16514 vdd.n1488 vdd.n876 146.341
R16515 vdd.n1499 vdd.n876 146.341
R16516 vdd.n1499 vdd.n871 146.341
R16517 vdd.n1507 vdd.n871 146.341
R16518 vdd.n1507 vdd.n861 146.341
R16519 vdd.n1944 vdd.n861 146.341
R16520 vdd.n1420 vdd.n1196 146.341
R16521 vdd.n1420 vdd.n1229 146.341
R16522 vdd.n1233 vdd.n1232 146.341
R16523 vdd.n1235 vdd.n1234 146.341
R16524 vdd.n1239 vdd.n1238 146.341
R16525 vdd.n1241 vdd.n1240 146.341
R16526 vdd.n1245 vdd.n1244 146.341
R16527 vdd.n1247 vdd.n1246 146.341
R16528 vdd.n1251 vdd.n1250 146.341
R16529 vdd.n1253 vdd.n1252 146.341
R16530 vdd.n1259 vdd.n1258 146.341
R16531 vdd.n1261 vdd.n1260 146.341
R16532 vdd.n1265 vdd.n1264 146.341
R16533 vdd.n1267 vdd.n1266 146.341
R16534 vdd.n1271 vdd.n1270 146.341
R16535 vdd.n1273 vdd.n1272 146.341
R16536 vdd.n1277 vdd.n1276 146.341
R16537 vdd.n1279 vdd.n1278 146.341
R16538 vdd.n1283 vdd.n1282 146.341
R16539 vdd.n1285 vdd.n1284 146.341
R16540 vdd.n1357 vdd.n1288 146.341
R16541 vdd.n1290 vdd.n1289 146.341
R16542 vdd.n1294 vdd.n1293 146.341
R16543 vdd.n1296 vdd.n1295 146.341
R16544 vdd.n1300 vdd.n1299 146.341
R16545 vdd.n1302 vdd.n1301 146.341
R16546 vdd.n1306 vdd.n1305 146.341
R16547 vdd.n1308 vdd.n1307 146.341
R16548 vdd.n1312 vdd.n1311 146.341
R16549 vdd.n1314 vdd.n1313 146.341
R16550 vdd.n1318 vdd.n1317 146.341
R16551 vdd.n1319 vdd.n1227 146.341
R16552 vdd.n1429 vdd.n1192 146.341
R16553 vdd.n1429 vdd.n1185 146.341
R16554 vdd.n1440 vdd.n1185 146.341
R16555 vdd.n1440 vdd.n1181 146.341
R16556 vdd.n1446 vdd.n1181 146.341
R16557 vdd.n1446 vdd.n1174 146.341
R16558 vdd.n1457 vdd.n1174 146.341
R16559 vdd.n1457 vdd.n1170 146.341
R16560 vdd.n1464 vdd.n1170 146.341
R16561 vdd.n1464 vdd.n1163 146.341
R16562 vdd.n1474 vdd.n1163 146.341
R16563 vdd.n1474 vdd.n889 146.341
R16564 vdd.n1480 vdd.n889 146.341
R16565 vdd.n1480 vdd.n881 146.341
R16566 vdd.n1491 vdd.n881 146.341
R16567 vdd.n1491 vdd.n877 146.341
R16568 vdd.n1497 vdd.n877 146.341
R16569 vdd.n1497 vdd.n869 146.341
R16570 vdd.n1510 vdd.n869 146.341
R16571 vdd.n1510 vdd.n864 146.341
R16572 vdd.n1942 vdd.n864 146.341
R16573 vdd.n863 vdd.n839 141.707
R16574 vdd.n2840 vdd.n484 141.707
R16575 vdd.n1791 vdd.t64 127.284
R16576 vdd.n755 vdd.t48 127.284
R16577 vdd.n1765 vdd.t89 127.284
R16578 vdd.n747 vdd.t79 127.284
R16579 vdd.n2536 vdd.t31 127.284
R16580 vdd.n2536 vdd.t32 127.284
R16581 vdd.n2256 vdd.t71 127.284
R16582 vdd.n622 vdd.t52 127.284
R16583 vdd.n2253 vdd.t57 127.284
R16584 vdd.n589 vdd.t59 127.284
R16585 vdd.n817 vdd.t67 127.284
R16586 vdd.n817 vdd.t68 127.284
R16587 vdd.n22 vdd.n20 117.314
R16588 vdd.n17 vdd.n15 117.314
R16589 vdd.n27 vdd.n26 116.927
R16590 vdd.n24 vdd.n23 116.927
R16591 vdd.n22 vdd.n21 116.927
R16592 vdd.n17 vdd.n16 116.927
R16593 vdd.n19 vdd.n18 116.927
R16594 vdd.n27 vdd.n25 116.927
R16595 vdd.n1792 vdd.t63 111.188
R16596 vdd.n756 vdd.t49 111.188
R16597 vdd.n1766 vdd.t88 111.188
R16598 vdd.n748 vdd.t80 111.188
R16599 vdd.n2257 vdd.t70 111.188
R16600 vdd.n623 vdd.t53 111.188
R16601 vdd.n2254 vdd.t56 111.188
R16602 vdd.n590 vdd.t60 111.188
R16603 vdd.n2479 vdd.n701 99.5127
R16604 vdd.n2483 vdd.n701 99.5127
R16605 vdd.n2483 vdd.n693 99.5127
R16606 vdd.n2491 vdd.n693 99.5127
R16607 vdd.n2491 vdd.n691 99.5127
R16608 vdd.n2495 vdd.n691 99.5127
R16609 vdd.n2495 vdd.n680 99.5127
R16610 vdd.n2503 vdd.n680 99.5127
R16611 vdd.n2503 vdd.n678 99.5127
R16612 vdd.n2507 vdd.n678 99.5127
R16613 vdd.n2507 vdd.n669 99.5127
R16614 vdd.n2515 vdd.n669 99.5127
R16615 vdd.n2515 vdd.n667 99.5127
R16616 vdd.n2519 vdd.n667 99.5127
R16617 vdd.n2519 vdd.n657 99.5127
R16618 vdd.n2527 vdd.n657 99.5127
R16619 vdd.n2527 vdd.n655 99.5127
R16620 vdd.n2531 vdd.n655 99.5127
R16621 vdd.n2531 vdd.n646 99.5127
R16622 vdd.n2541 vdd.n646 99.5127
R16623 vdd.n2541 vdd.n644 99.5127
R16624 vdd.n2545 vdd.n644 99.5127
R16625 vdd.n2545 vdd.n632 99.5127
R16626 vdd.n2598 vdd.n632 99.5127
R16627 vdd.n2598 vdd.n630 99.5127
R16628 vdd.n2602 vdd.n630 99.5127
R16629 vdd.n2602 vdd.n598 99.5127
R16630 vdd.n2672 vdd.n598 99.5127
R16631 vdd.n2668 vdd.n599 99.5127
R16632 vdd.n2666 vdd.n2665 99.5127
R16633 vdd.n2663 vdd.n603 99.5127
R16634 vdd.n2659 vdd.n2658 99.5127
R16635 vdd.n2656 vdd.n606 99.5127
R16636 vdd.n2652 vdd.n2651 99.5127
R16637 vdd.n2649 vdd.n609 99.5127
R16638 vdd.n2645 vdd.n2644 99.5127
R16639 vdd.n2642 vdd.n2640 99.5127
R16640 vdd.n2638 vdd.n612 99.5127
R16641 vdd.n2634 vdd.n2633 99.5127
R16642 vdd.n2631 vdd.n615 99.5127
R16643 vdd.n2627 vdd.n2626 99.5127
R16644 vdd.n2624 vdd.n618 99.5127
R16645 vdd.n2620 vdd.n2619 99.5127
R16646 vdd.n2617 vdd.n621 99.5127
R16647 vdd.n2612 vdd.n2611 99.5127
R16648 vdd.n2399 vdd.n704 99.5127
R16649 vdd.n2399 vdd.n699 99.5127
R16650 vdd.n2396 vdd.n699 99.5127
R16651 vdd.n2396 vdd.n694 99.5127
R16652 vdd.n2343 vdd.n694 99.5127
R16653 vdd.n2343 vdd.n688 99.5127
R16654 vdd.n2346 vdd.n688 99.5127
R16655 vdd.n2346 vdd.n681 99.5127
R16656 vdd.n2349 vdd.n681 99.5127
R16657 vdd.n2349 vdd.n676 99.5127
R16658 vdd.n2352 vdd.n676 99.5127
R16659 vdd.n2352 vdd.n671 99.5127
R16660 vdd.n2355 vdd.n671 99.5127
R16661 vdd.n2355 vdd.n665 99.5127
R16662 vdd.n2373 vdd.n665 99.5127
R16663 vdd.n2373 vdd.n658 99.5127
R16664 vdd.n2369 vdd.n658 99.5127
R16665 vdd.n2369 vdd.n653 99.5127
R16666 vdd.n2366 vdd.n653 99.5127
R16667 vdd.n2366 vdd.n648 99.5127
R16668 vdd.n2363 vdd.n648 99.5127
R16669 vdd.n2363 vdd.n642 99.5127
R16670 vdd.n2360 vdd.n642 99.5127
R16671 vdd.n2360 vdd.n634 99.5127
R16672 vdd.n634 vdd.n627 99.5127
R16673 vdd.n2604 vdd.n627 99.5127
R16674 vdd.n2605 vdd.n2604 99.5127
R16675 vdd.n2605 vdd.n596 99.5127
R16676 vdd.n2469 vdd.n2252 99.5127
R16677 vdd.n2465 vdd.n2252 99.5127
R16678 vdd.n2463 vdd.n2462 99.5127
R16679 vdd.n2459 vdd.n2458 99.5127
R16680 vdd.n2455 vdd.n2454 99.5127
R16681 vdd.n2451 vdd.n2450 99.5127
R16682 vdd.n2447 vdd.n2446 99.5127
R16683 vdd.n2443 vdd.n2442 99.5127
R16684 vdd.n2439 vdd.n2438 99.5127
R16685 vdd.n2435 vdd.n2434 99.5127
R16686 vdd.n2431 vdd.n2430 99.5127
R16687 vdd.n2427 vdd.n2426 99.5127
R16688 vdd.n2423 vdd.n2422 99.5127
R16689 vdd.n2419 vdd.n2418 99.5127
R16690 vdd.n2415 vdd.n2414 99.5127
R16691 vdd.n2411 vdd.n2410 99.5127
R16692 vdd.n2406 vdd.n2405 99.5127
R16693 vdd.n2217 vdd.n745 99.5127
R16694 vdd.n2213 vdd.n2212 99.5127
R16695 vdd.n2209 vdd.n2208 99.5127
R16696 vdd.n2205 vdd.n2204 99.5127
R16697 vdd.n2201 vdd.n2200 99.5127
R16698 vdd.n2197 vdd.n2196 99.5127
R16699 vdd.n2193 vdd.n2192 99.5127
R16700 vdd.n2189 vdd.n2188 99.5127
R16701 vdd.n2185 vdd.n2184 99.5127
R16702 vdd.n2181 vdd.n2180 99.5127
R16703 vdd.n2177 vdd.n2176 99.5127
R16704 vdd.n2173 vdd.n2172 99.5127
R16705 vdd.n2169 vdd.n2168 99.5127
R16706 vdd.n2165 vdd.n2164 99.5127
R16707 vdd.n2161 vdd.n2160 99.5127
R16708 vdd.n2157 vdd.n2156 99.5127
R16709 vdd.n2152 vdd.n2151 99.5127
R16710 vdd.n1890 vdd.n840 99.5127
R16711 vdd.n1890 vdd.n834 99.5127
R16712 vdd.n1887 vdd.n834 99.5127
R16713 vdd.n1887 vdd.n828 99.5127
R16714 vdd.n1884 vdd.n828 99.5127
R16715 vdd.n1884 vdd.n821 99.5127
R16716 vdd.n1881 vdd.n821 99.5127
R16717 vdd.n1881 vdd.n814 99.5127
R16718 vdd.n1878 vdd.n814 99.5127
R16719 vdd.n1878 vdd.n809 99.5127
R16720 vdd.n1875 vdd.n809 99.5127
R16721 vdd.n1875 vdd.n803 99.5127
R16722 vdd.n1872 vdd.n803 99.5127
R16723 vdd.n1872 vdd.n796 99.5127
R16724 vdd.n1786 vdd.n796 99.5127
R16725 vdd.n1786 vdd.n790 99.5127
R16726 vdd.n1783 vdd.n790 99.5127
R16727 vdd.n1783 vdd.n785 99.5127
R16728 vdd.n1780 vdd.n785 99.5127
R16729 vdd.n1780 vdd.n780 99.5127
R16730 vdd.n1777 vdd.n780 99.5127
R16731 vdd.n1777 vdd.n774 99.5127
R16732 vdd.n1774 vdd.n774 99.5127
R16733 vdd.n1774 vdd.n767 99.5127
R16734 vdd.n1771 vdd.n767 99.5127
R16735 vdd.n1771 vdd.n760 99.5127
R16736 vdd.n760 vdd.n750 99.5127
R16737 vdd.n2147 vdd.n750 99.5127
R16738 vdd.n1725 vdd.n1723 99.5127
R16739 vdd.n1729 vdd.n1723 99.5127
R16740 vdd.n1733 vdd.n1731 99.5127
R16741 vdd.n1737 vdd.n1721 99.5127
R16742 vdd.n1741 vdd.n1739 99.5127
R16743 vdd.n1745 vdd.n1719 99.5127
R16744 vdd.n1749 vdd.n1747 99.5127
R16745 vdd.n1753 vdd.n1717 99.5127
R16746 vdd.n1756 vdd.n1755 99.5127
R16747 vdd.n1926 vdd.n1924 99.5127
R16748 vdd.n1922 vdd.n1758 99.5127
R16749 vdd.n1918 vdd.n1916 99.5127
R16750 vdd.n1914 vdd.n1760 99.5127
R16751 vdd.n1910 vdd.n1908 99.5127
R16752 vdd.n1906 vdd.n1762 99.5127
R16753 vdd.n1902 vdd.n1900 99.5127
R16754 vdd.n1898 vdd.n1764 99.5127
R16755 vdd.n1990 vdd.n836 99.5127
R16756 vdd.n1994 vdd.n836 99.5127
R16757 vdd.n1994 vdd.n826 99.5127
R16758 vdd.n2002 vdd.n826 99.5127
R16759 vdd.n2002 vdd.n824 99.5127
R16760 vdd.n2006 vdd.n824 99.5127
R16761 vdd.n2006 vdd.n813 99.5127
R16762 vdd.n2015 vdd.n813 99.5127
R16763 vdd.n2015 vdd.n811 99.5127
R16764 vdd.n2019 vdd.n811 99.5127
R16765 vdd.n2019 vdd.n801 99.5127
R16766 vdd.n2027 vdd.n801 99.5127
R16767 vdd.n2027 vdd.n799 99.5127
R16768 vdd.n2031 vdd.n799 99.5127
R16769 vdd.n2031 vdd.n789 99.5127
R16770 vdd.n2039 vdd.n789 99.5127
R16771 vdd.n2039 vdd.n787 99.5127
R16772 vdd.n2043 vdd.n787 99.5127
R16773 vdd.n2043 vdd.n778 99.5127
R16774 vdd.n2051 vdd.n778 99.5127
R16775 vdd.n2051 vdd.n776 99.5127
R16776 vdd.n2055 vdd.n776 99.5127
R16777 vdd.n2055 vdd.n765 99.5127
R16778 vdd.n2065 vdd.n765 99.5127
R16779 vdd.n2065 vdd.n762 99.5127
R16780 vdd.n2070 vdd.n762 99.5127
R16781 vdd.n2070 vdd.n763 99.5127
R16782 vdd.n763 vdd.n744 99.5127
R16783 vdd.n2588 vdd.n2587 99.5127
R16784 vdd.n2585 vdd.n2551 99.5127
R16785 vdd.n2581 vdd.n2580 99.5127
R16786 vdd.n2578 vdd.n2554 99.5127
R16787 vdd.n2574 vdd.n2573 99.5127
R16788 vdd.n2571 vdd.n2557 99.5127
R16789 vdd.n2567 vdd.n2566 99.5127
R16790 vdd.n2564 vdd.n2561 99.5127
R16791 vdd.n2705 vdd.n577 99.5127
R16792 vdd.n2703 vdd.n2702 99.5127
R16793 vdd.n2700 vdd.n579 99.5127
R16794 vdd.n2696 vdd.n2695 99.5127
R16795 vdd.n2693 vdd.n582 99.5127
R16796 vdd.n2689 vdd.n2688 99.5127
R16797 vdd.n2686 vdd.n585 99.5127
R16798 vdd.n2682 vdd.n2681 99.5127
R16799 vdd.n2679 vdd.n588 99.5127
R16800 vdd.n2323 vdd.n705 99.5127
R16801 vdd.n2323 vdd.n700 99.5127
R16802 vdd.n2394 vdd.n700 99.5127
R16803 vdd.n2394 vdd.n695 99.5127
R16804 vdd.n2390 vdd.n695 99.5127
R16805 vdd.n2390 vdd.n689 99.5127
R16806 vdd.n2387 vdd.n689 99.5127
R16807 vdd.n2387 vdd.n682 99.5127
R16808 vdd.n2384 vdd.n682 99.5127
R16809 vdd.n2384 vdd.n677 99.5127
R16810 vdd.n2381 vdd.n677 99.5127
R16811 vdd.n2381 vdd.n672 99.5127
R16812 vdd.n2378 vdd.n672 99.5127
R16813 vdd.n2378 vdd.n666 99.5127
R16814 vdd.n2375 vdd.n666 99.5127
R16815 vdd.n2375 vdd.n659 99.5127
R16816 vdd.n2340 vdd.n659 99.5127
R16817 vdd.n2340 vdd.n654 99.5127
R16818 vdd.n2337 vdd.n654 99.5127
R16819 vdd.n2337 vdd.n649 99.5127
R16820 vdd.n2334 vdd.n649 99.5127
R16821 vdd.n2334 vdd.n643 99.5127
R16822 vdd.n2331 vdd.n643 99.5127
R16823 vdd.n2331 vdd.n635 99.5127
R16824 vdd.n2328 vdd.n635 99.5127
R16825 vdd.n2328 vdd.n628 99.5127
R16826 vdd.n628 vdd.n594 99.5127
R16827 vdd.n2674 vdd.n594 99.5127
R16828 vdd.n2473 vdd.n708 99.5127
R16829 vdd.n2261 vdd.n2260 99.5127
R16830 vdd.n2265 vdd.n2264 99.5127
R16831 vdd.n2269 vdd.n2268 99.5127
R16832 vdd.n2273 vdd.n2272 99.5127
R16833 vdd.n2277 vdd.n2276 99.5127
R16834 vdd.n2281 vdd.n2280 99.5127
R16835 vdd.n2285 vdd.n2284 99.5127
R16836 vdd.n2289 vdd.n2288 99.5127
R16837 vdd.n2293 vdd.n2292 99.5127
R16838 vdd.n2297 vdd.n2296 99.5127
R16839 vdd.n2301 vdd.n2300 99.5127
R16840 vdd.n2305 vdd.n2304 99.5127
R16841 vdd.n2309 vdd.n2308 99.5127
R16842 vdd.n2313 vdd.n2312 99.5127
R16843 vdd.n2317 vdd.n2316 99.5127
R16844 vdd.n2319 vdd.n2251 99.5127
R16845 vdd.n2477 vdd.n698 99.5127
R16846 vdd.n2485 vdd.n698 99.5127
R16847 vdd.n2485 vdd.n696 99.5127
R16848 vdd.n2489 vdd.n696 99.5127
R16849 vdd.n2489 vdd.n686 99.5127
R16850 vdd.n2497 vdd.n686 99.5127
R16851 vdd.n2497 vdd.n684 99.5127
R16852 vdd.n2501 vdd.n684 99.5127
R16853 vdd.n2501 vdd.n675 99.5127
R16854 vdd.n2509 vdd.n675 99.5127
R16855 vdd.n2509 vdd.n673 99.5127
R16856 vdd.n2513 vdd.n673 99.5127
R16857 vdd.n2513 vdd.n663 99.5127
R16858 vdd.n2521 vdd.n663 99.5127
R16859 vdd.n2521 vdd.n661 99.5127
R16860 vdd.n2525 vdd.n661 99.5127
R16861 vdd.n2525 vdd.n652 99.5127
R16862 vdd.n2533 vdd.n652 99.5127
R16863 vdd.n2533 vdd.n650 99.5127
R16864 vdd.n2539 vdd.n650 99.5127
R16865 vdd.n2539 vdd.n640 99.5127
R16866 vdd.n2547 vdd.n640 99.5127
R16867 vdd.n2547 vdd.n637 99.5127
R16868 vdd.n2596 vdd.n637 99.5127
R16869 vdd.n2596 vdd.n638 99.5127
R16870 vdd.n638 vdd.n629 99.5127
R16871 vdd.n2591 vdd.n629 99.5127
R16872 vdd.n2591 vdd.n597 99.5127
R16873 vdd.n2141 vdd.n2140 99.5127
R16874 vdd.n2137 vdd.n2136 99.5127
R16875 vdd.n2133 vdd.n2132 99.5127
R16876 vdd.n2129 vdd.n2128 99.5127
R16877 vdd.n2125 vdd.n2124 99.5127
R16878 vdd.n2121 vdd.n2120 99.5127
R16879 vdd.n2117 vdd.n2116 99.5127
R16880 vdd.n2113 vdd.n2112 99.5127
R16881 vdd.n2109 vdd.n2108 99.5127
R16882 vdd.n2105 vdd.n2104 99.5127
R16883 vdd.n2101 vdd.n2100 99.5127
R16884 vdd.n2097 vdd.n2096 99.5127
R16885 vdd.n2093 vdd.n2092 99.5127
R16886 vdd.n2089 vdd.n2088 99.5127
R16887 vdd.n2085 vdd.n2084 99.5127
R16888 vdd.n2081 vdd.n2080 99.5127
R16889 vdd.n2077 vdd.n726 99.5127
R16890 vdd.n1834 vdd.n841 99.5127
R16891 vdd.n1834 vdd.n835 99.5127
R16892 vdd.n1837 vdd.n835 99.5127
R16893 vdd.n1837 vdd.n829 99.5127
R16894 vdd.n1840 vdd.n829 99.5127
R16895 vdd.n1840 vdd.n822 99.5127
R16896 vdd.n1843 vdd.n822 99.5127
R16897 vdd.n1843 vdd.n815 99.5127
R16898 vdd.n1846 vdd.n815 99.5127
R16899 vdd.n1846 vdd.n810 99.5127
R16900 vdd.n1849 vdd.n810 99.5127
R16901 vdd.n1849 vdd.n804 99.5127
R16902 vdd.n1870 vdd.n804 99.5127
R16903 vdd.n1870 vdd.n797 99.5127
R16904 vdd.n1866 vdd.n797 99.5127
R16905 vdd.n1866 vdd.n791 99.5127
R16906 vdd.n1863 vdd.n791 99.5127
R16907 vdd.n1863 vdd.n786 99.5127
R16908 vdd.n1860 vdd.n786 99.5127
R16909 vdd.n1860 vdd.n781 99.5127
R16910 vdd.n1857 vdd.n781 99.5127
R16911 vdd.n1857 vdd.n775 99.5127
R16912 vdd.n1854 vdd.n775 99.5127
R16913 vdd.n1854 vdd.n768 99.5127
R16914 vdd.n768 vdd.n759 99.5127
R16915 vdd.n2072 vdd.n759 99.5127
R16916 vdd.n2073 vdd.n2072 99.5127
R16917 vdd.n2073 vdd.n751 99.5127
R16918 vdd.n1984 vdd.n1982 99.5127
R16919 vdd.n1980 vdd.n844 99.5127
R16920 vdd.n1976 vdd.n1974 99.5127
R16921 vdd.n1972 vdd.n846 99.5127
R16922 vdd.n1968 vdd.n1966 99.5127
R16923 vdd.n1964 vdd.n848 99.5127
R16924 vdd.n1960 vdd.n1958 99.5127
R16925 vdd.n1956 vdd.n850 99.5127
R16926 vdd.n1798 vdd.n852 99.5127
R16927 vdd.n1803 vdd.n1800 99.5127
R16928 vdd.n1807 vdd.n1805 99.5127
R16929 vdd.n1811 vdd.n1796 99.5127
R16930 vdd.n1815 vdd.n1813 99.5127
R16931 vdd.n1819 vdd.n1794 99.5127
R16932 vdd.n1823 vdd.n1821 99.5127
R16933 vdd.n1828 vdd.n1790 99.5127
R16934 vdd.n1831 vdd.n1830 99.5127
R16935 vdd.n1988 vdd.n832 99.5127
R16936 vdd.n1996 vdd.n832 99.5127
R16937 vdd.n1996 vdd.n830 99.5127
R16938 vdd.n2000 vdd.n830 99.5127
R16939 vdd.n2000 vdd.n819 99.5127
R16940 vdd.n2008 vdd.n819 99.5127
R16941 vdd.n2008 vdd.n816 99.5127
R16942 vdd.n2013 vdd.n816 99.5127
R16943 vdd.n2013 vdd.n807 99.5127
R16944 vdd.n2021 vdd.n807 99.5127
R16945 vdd.n2021 vdd.n805 99.5127
R16946 vdd.n2025 vdd.n805 99.5127
R16947 vdd.n2025 vdd.n795 99.5127
R16948 vdd.n2033 vdd.n795 99.5127
R16949 vdd.n2033 vdd.n793 99.5127
R16950 vdd.n2037 vdd.n793 99.5127
R16951 vdd.n2037 vdd.n784 99.5127
R16952 vdd.n2045 vdd.n784 99.5127
R16953 vdd.n2045 vdd.n782 99.5127
R16954 vdd.n2049 vdd.n782 99.5127
R16955 vdd.n2049 vdd.n772 99.5127
R16956 vdd.n2057 vdd.n772 99.5127
R16957 vdd.n2057 vdd.n769 99.5127
R16958 vdd.n2063 vdd.n769 99.5127
R16959 vdd.n2063 vdd.n770 99.5127
R16960 vdd.n770 vdd.n761 99.5127
R16961 vdd.n761 vdd.n752 99.5127
R16962 vdd.n2145 vdd.n752 99.5127
R16963 vdd.n9 vdd.n7 98.9633
R16964 vdd.n2 vdd.n0 98.9633
R16965 vdd.n9 vdd.n8 98.6055
R16966 vdd.n11 vdd.n10 98.6055
R16967 vdd.n13 vdd.n12 98.6055
R16968 vdd.n6 vdd.n5 98.6055
R16969 vdd.n4 vdd.n3 98.6055
R16970 vdd.n2 vdd.n1 98.6055
R16971 vdd.t136 vdd.n267 85.8723
R16972 vdd.t147 vdd.n220 85.8723
R16973 vdd.t132 vdd.n177 85.8723
R16974 vdd.t142 vdd.n130 85.8723
R16975 vdd.t173 vdd.n88 85.8723
R16976 vdd.t115 vdd.n41 85.8723
R16977 vdd.t171 vdd.n1082 85.8723
R16978 vdd.t157 vdd.n1129 85.8723
R16979 vdd.t163 vdd.n992 85.8723
R16980 vdd.t150 vdd.n1039 85.8723
R16981 vdd.t113 vdd.n903 85.8723
R16982 vdd.t172 vdd.n950 85.8723
R16983 vdd.n2537 vdd.n2536 78.546
R16984 vdd.n2011 vdd.n817 78.546
R16985 vdd.n254 vdd.n253 75.1835
R16986 vdd.n252 vdd.n251 75.1835
R16987 vdd.n250 vdd.n249 75.1835
R16988 vdd.n164 vdd.n163 75.1835
R16989 vdd.n162 vdd.n161 75.1835
R16990 vdd.n160 vdd.n159 75.1835
R16991 vdd.n75 vdd.n74 75.1835
R16992 vdd.n73 vdd.n72 75.1835
R16993 vdd.n71 vdd.n70 75.1835
R16994 vdd.n1112 vdd.n1111 75.1835
R16995 vdd.n1114 vdd.n1113 75.1835
R16996 vdd.n1116 vdd.n1115 75.1835
R16997 vdd.n1022 vdd.n1021 75.1835
R16998 vdd.n1024 vdd.n1023 75.1835
R16999 vdd.n1026 vdd.n1025 75.1835
R17000 vdd.n933 vdd.n932 75.1835
R17001 vdd.n935 vdd.n934 75.1835
R17002 vdd.n937 vdd.n936 75.1835
R17003 vdd.n2472 vdd.n2471 72.8958
R17004 vdd.n2471 vdd.n2235 72.8958
R17005 vdd.n2471 vdd.n2236 72.8958
R17006 vdd.n2471 vdd.n2237 72.8958
R17007 vdd.n2471 vdd.n2238 72.8958
R17008 vdd.n2471 vdd.n2239 72.8958
R17009 vdd.n2471 vdd.n2240 72.8958
R17010 vdd.n2471 vdd.n2241 72.8958
R17011 vdd.n2471 vdd.n2242 72.8958
R17012 vdd.n2471 vdd.n2243 72.8958
R17013 vdd.n2471 vdd.n2244 72.8958
R17014 vdd.n2471 vdd.n2245 72.8958
R17015 vdd.n2471 vdd.n2246 72.8958
R17016 vdd.n2471 vdd.n2247 72.8958
R17017 vdd.n2471 vdd.n2248 72.8958
R17018 vdd.n2471 vdd.n2249 72.8958
R17019 vdd.n2471 vdd.n2250 72.8958
R17020 vdd.n593 vdd.n484 72.8958
R17021 vdd.n2680 vdd.n484 72.8958
R17022 vdd.n587 vdd.n484 72.8958
R17023 vdd.n2687 vdd.n484 72.8958
R17024 vdd.n584 vdd.n484 72.8958
R17025 vdd.n2694 vdd.n484 72.8958
R17026 vdd.n581 vdd.n484 72.8958
R17027 vdd.n2701 vdd.n484 72.8958
R17028 vdd.n2704 vdd.n484 72.8958
R17029 vdd.n2560 vdd.n484 72.8958
R17030 vdd.n2565 vdd.n484 72.8958
R17031 vdd.n2559 vdd.n484 72.8958
R17032 vdd.n2572 vdd.n484 72.8958
R17033 vdd.n2556 vdd.n484 72.8958
R17034 vdd.n2579 vdd.n484 72.8958
R17035 vdd.n2553 vdd.n484 72.8958
R17036 vdd.n2586 vdd.n484 72.8958
R17037 vdd.n1724 vdd.n839 72.8958
R17038 vdd.n1730 vdd.n839 72.8958
R17039 vdd.n1732 vdd.n839 72.8958
R17040 vdd.n1738 vdd.n839 72.8958
R17041 vdd.n1740 vdd.n839 72.8958
R17042 vdd.n1746 vdd.n839 72.8958
R17043 vdd.n1748 vdd.n839 72.8958
R17044 vdd.n1754 vdd.n839 72.8958
R17045 vdd.n1925 vdd.n839 72.8958
R17046 vdd.n1923 vdd.n839 72.8958
R17047 vdd.n1917 vdd.n839 72.8958
R17048 vdd.n1915 vdd.n839 72.8958
R17049 vdd.n1909 vdd.n839 72.8958
R17050 vdd.n1907 vdd.n839 72.8958
R17051 vdd.n1901 vdd.n839 72.8958
R17052 vdd.n1899 vdd.n839 72.8958
R17053 vdd.n1893 vdd.n839 72.8958
R17054 vdd.n2218 vdd.n727 72.8958
R17055 vdd.n2218 vdd.n728 72.8958
R17056 vdd.n2218 vdd.n729 72.8958
R17057 vdd.n2218 vdd.n730 72.8958
R17058 vdd.n2218 vdd.n731 72.8958
R17059 vdd.n2218 vdd.n732 72.8958
R17060 vdd.n2218 vdd.n733 72.8958
R17061 vdd.n2218 vdd.n734 72.8958
R17062 vdd.n2218 vdd.n735 72.8958
R17063 vdd.n2218 vdd.n736 72.8958
R17064 vdd.n2218 vdd.n737 72.8958
R17065 vdd.n2218 vdd.n738 72.8958
R17066 vdd.n2218 vdd.n739 72.8958
R17067 vdd.n2218 vdd.n740 72.8958
R17068 vdd.n2218 vdd.n741 72.8958
R17069 vdd.n2218 vdd.n742 72.8958
R17070 vdd.n2218 vdd.n743 72.8958
R17071 vdd.n2471 vdd.n2470 72.8958
R17072 vdd.n2471 vdd.n2219 72.8958
R17073 vdd.n2471 vdd.n2220 72.8958
R17074 vdd.n2471 vdd.n2221 72.8958
R17075 vdd.n2471 vdd.n2222 72.8958
R17076 vdd.n2471 vdd.n2223 72.8958
R17077 vdd.n2471 vdd.n2224 72.8958
R17078 vdd.n2471 vdd.n2225 72.8958
R17079 vdd.n2471 vdd.n2226 72.8958
R17080 vdd.n2471 vdd.n2227 72.8958
R17081 vdd.n2471 vdd.n2228 72.8958
R17082 vdd.n2471 vdd.n2229 72.8958
R17083 vdd.n2471 vdd.n2230 72.8958
R17084 vdd.n2471 vdd.n2231 72.8958
R17085 vdd.n2471 vdd.n2232 72.8958
R17086 vdd.n2471 vdd.n2233 72.8958
R17087 vdd.n2471 vdd.n2234 72.8958
R17088 vdd.n2610 vdd.n484 72.8958
R17089 vdd.n625 vdd.n484 72.8958
R17090 vdd.n2618 vdd.n484 72.8958
R17091 vdd.n620 vdd.n484 72.8958
R17092 vdd.n2625 vdd.n484 72.8958
R17093 vdd.n617 vdd.n484 72.8958
R17094 vdd.n2632 vdd.n484 72.8958
R17095 vdd.n614 vdd.n484 72.8958
R17096 vdd.n2639 vdd.n484 72.8958
R17097 vdd.n2643 vdd.n484 72.8958
R17098 vdd.n611 vdd.n484 72.8958
R17099 vdd.n2650 vdd.n484 72.8958
R17100 vdd.n608 vdd.n484 72.8958
R17101 vdd.n2657 vdd.n484 72.8958
R17102 vdd.n605 vdd.n484 72.8958
R17103 vdd.n2664 vdd.n484 72.8958
R17104 vdd.n2667 vdd.n484 72.8958
R17105 vdd.n2218 vdd.n725 72.8958
R17106 vdd.n2218 vdd.n724 72.8958
R17107 vdd.n2218 vdd.n723 72.8958
R17108 vdd.n2218 vdd.n722 72.8958
R17109 vdd.n2218 vdd.n721 72.8958
R17110 vdd.n2218 vdd.n720 72.8958
R17111 vdd.n2218 vdd.n719 72.8958
R17112 vdd.n2218 vdd.n718 72.8958
R17113 vdd.n2218 vdd.n717 72.8958
R17114 vdd.n2218 vdd.n716 72.8958
R17115 vdd.n2218 vdd.n715 72.8958
R17116 vdd.n2218 vdd.n714 72.8958
R17117 vdd.n2218 vdd.n713 72.8958
R17118 vdd.n2218 vdd.n712 72.8958
R17119 vdd.n2218 vdd.n711 72.8958
R17120 vdd.n2218 vdd.n710 72.8958
R17121 vdd.n2218 vdd.n709 72.8958
R17122 vdd.n1983 vdd.n839 72.8958
R17123 vdd.n1981 vdd.n839 72.8958
R17124 vdd.n1975 vdd.n839 72.8958
R17125 vdd.n1973 vdd.n839 72.8958
R17126 vdd.n1967 vdd.n839 72.8958
R17127 vdd.n1965 vdd.n839 72.8958
R17128 vdd.n1959 vdd.n839 72.8958
R17129 vdd.n1957 vdd.n839 72.8958
R17130 vdd.n851 vdd.n839 72.8958
R17131 vdd.n1799 vdd.n839 72.8958
R17132 vdd.n1804 vdd.n839 72.8958
R17133 vdd.n1806 vdd.n839 72.8958
R17134 vdd.n1812 vdd.n839 72.8958
R17135 vdd.n1814 vdd.n839 72.8958
R17136 vdd.n1820 vdd.n839 72.8958
R17137 vdd.n1822 vdd.n839 72.8958
R17138 vdd.n1829 vdd.n839 72.8958
R17139 vdd.n1422 vdd.n1421 66.2847
R17140 vdd.n1421 vdd.n1197 66.2847
R17141 vdd.n1421 vdd.n1198 66.2847
R17142 vdd.n1421 vdd.n1199 66.2847
R17143 vdd.n1421 vdd.n1200 66.2847
R17144 vdd.n1421 vdd.n1201 66.2847
R17145 vdd.n1421 vdd.n1202 66.2847
R17146 vdd.n1421 vdd.n1203 66.2847
R17147 vdd.n1421 vdd.n1204 66.2847
R17148 vdd.n1421 vdd.n1205 66.2847
R17149 vdd.n1421 vdd.n1206 66.2847
R17150 vdd.n1421 vdd.n1207 66.2847
R17151 vdd.n1421 vdd.n1208 66.2847
R17152 vdd.n1421 vdd.n1209 66.2847
R17153 vdd.n1421 vdd.n1210 66.2847
R17154 vdd.n1421 vdd.n1211 66.2847
R17155 vdd.n1421 vdd.n1212 66.2847
R17156 vdd.n1421 vdd.n1213 66.2847
R17157 vdd.n1421 vdd.n1214 66.2847
R17158 vdd.n1421 vdd.n1215 66.2847
R17159 vdd.n1421 vdd.n1216 66.2847
R17160 vdd.n1421 vdd.n1217 66.2847
R17161 vdd.n1421 vdd.n1218 66.2847
R17162 vdd.n1421 vdd.n1219 66.2847
R17163 vdd.n1421 vdd.n1220 66.2847
R17164 vdd.n1421 vdd.n1221 66.2847
R17165 vdd.n1421 vdd.n1222 66.2847
R17166 vdd.n1421 vdd.n1223 66.2847
R17167 vdd.n1421 vdd.n1224 66.2847
R17168 vdd.n1421 vdd.n1225 66.2847
R17169 vdd.n1421 vdd.n1226 66.2847
R17170 vdd.n863 vdd.n860 66.2847
R17171 vdd.n1614 vdd.n863 66.2847
R17172 vdd.n1619 vdd.n863 66.2847
R17173 vdd.n1624 vdd.n863 66.2847
R17174 vdd.n1612 vdd.n863 66.2847
R17175 vdd.n1631 vdd.n863 66.2847
R17176 vdd.n1604 vdd.n863 66.2847
R17177 vdd.n1638 vdd.n863 66.2847
R17178 vdd.n1597 vdd.n863 66.2847
R17179 vdd.n1645 vdd.n863 66.2847
R17180 vdd.n1591 vdd.n863 66.2847
R17181 vdd.n1586 vdd.n863 66.2847
R17182 vdd.n1656 vdd.n863 66.2847
R17183 vdd.n1578 vdd.n863 66.2847
R17184 vdd.n1663 vdd.n863 66.2847
R17185 vdd.n1571 vdd.n863 66.2847
R17186 vdd.n1670 vdd.n863 66.2847
R17187 vdd.n1564 vdd.n863 66.2847
R17188 vdd.n1677 vdd.n863 66.2847
R17189 vdd.n1557 vdd.n863 66.2847
R17190 vdd.n1684 vdd.n863 66.2847
R17191 vdd.n1551 vdd.n863 66.2847
R17192 vdd.n1546 vdd.n863 66.2847
R17193 vdd.n1695 vdd.n863 66.2847
R17194 vdd.n1538 vdd.n863 66.2847
R17195 vdd.n1702 vdd.n863 66.2847
R17196 vdd.n1531 vdd.n863 66.2847
R17197 vdd.n1709 vdd.n863 66.2847
R17198 vdd.n1712 vdd.n863 66.2847
R17199 vdd.n1522 vdd.n863 66.2847
R17200 vdd.n1934 vdd.n863 66.2847
R17201 vdd.n1516 vdd.n863 66.2847
R17202 vdd.n2841 vdd.n2840 66.2847
R17203 vdd.n2840 vdd.n485 66.2847
R17204 vdd.n2840 vdd.n486 66.2847
R17205 vdd.n2840 vdd.n487 66.2847
R17206 vdd.n2840 vdd.n488 66.2847
R17207 vdd.n2840 vdd.n489 66.2847
R17208 vdd.n2840 vdd.n490 66.2847
R17209 vdd.n2840 vdd.n491 66.2847
R17210 vdd.n2840 vdd.n492 66.2847
R17211 vdd.n2840 vdd.n493 66.2847
R17212 vdd.n2840 vdd.n494 66.2847
R17213 vdd.n2840 vdd.n495 66.2847
R17214 vdd.n2840 vdd.n496 66.2847
R17215 vdd.n2840 vdd.n497 66.2847
R17216 vdd.n2840 vdd.n498 66.2847
R17217 vdd.n2840 vdd.n499 66.2847
R17218 vdd.n2840 vdd.n500 66.2847
R17219 vdd.n2840 vdd.n501 66.2847
R17220 vdd.n2840 vdd.n502 66.2847
R17221 vdd.n2840 vdd.n503 66.2847
R17222 vdd.n2840 vdd.n504 66.2847
R17223 vdd.n2840 vdd.n505 66.2847
R17224 vdd.n2840 vdd.n506 66.2847
R17225 vdd.n2840 vdd.n507 66.2847
R17226 vdd.n2840 vdd.n508 66.2847
R17227 vdd.n2840 vdd.n509 66.2847
R17228 vdd.n2840 vdd.n510 66.2847
R17229 vdd.n2840 vdd.n511 66.2847
R17230 vdd.n2840 vdd.n512 66.2847
R17231 vdd.n2840 vdd.n513 66.2847
R17232 vdd.n2840 vdd.n514 66.2847
R17233 vdd.n2905 vdd.n329 66.2847
R17234 vdd.n2914 vdd.n329 66.2847
R17235 vdd.n439 vdd.n329 66.2847
R17236 vdd.n2921 vdd.n329 66.2847
R17237 vdd.n432 vdd.n329 66.2847
R17238 vdd.n2928 vdd.n329 66.2847
R17239 vdd.n425 vdd.n329 66.2847
R17240 vdd.n2935 vdd.n329 66.2847
R17241 vdd.n418 vdd.n329 66.2847
R17242 vdd.n2942 vdd.n329 66.2847
R17243 vdd.n412 vdd.n329 66.2847
R17244 vdd.n407 vdd.n329 66.2847
R17245 vdd.n2953 vdd.n329 66.2847
R17246 vdd.n399 vdd.n329 66.2847
R17247 vdd.n2960 vdd.n329 66.2847
R17248 vdd.n392 vdd.n329 66.2847
R17249 vdd.n2967 vdd.n329 66.2847
R17250 vdd.n385 vdd.n329 66.2847
R17251 vdd.n2974 vdd.n329 66.2847
R17252 vdd.n378 vdd.n329 66.2847
R17253 vdd.n2981 vdd.n329 66.2847
R17254 vdd.n372 vdd.n329 66.2847
R17255 vdd.n367 vdd.n329 66.2847
R17256 vdd.n2992 vdd.n329 66.2847
R17257 vdd.n359 vdd.n329 66.2847
R17258 vdd.n2999 vdd.n329 66.2847
R17259 vdd.n352 vdd.n329 66.2847
R17260 vdd.n3006 vdd.n329 66.2847
R17261 vdd.n345 vdd.n329 66.2847
R17262 vdd.n3013 vdd.n329 66.2847
R17263 vdd.n3016 vdd.n329 66.2847
R17264 vdd.n333 vdd.n329 66.2847
R17265 vdd.n334 vdd.n333 52.4337
R17266 vdd.n3016 vdd.n3015 52.4337
R17267 vdd.n3013 vdd.n3012 52.4337
R17268 vdd.n3008 vdd.n345 52.4337
R17269 vdd.n3006 vdd.n3005 52.4337
R17270 vdd.n3001 vdd.n352 52.4337
R17271 vdd.n2999 vdd.n2998 52.4337
R17272 vdd.n2994 vdd.n359 52.4337
R17273 vdd.n2992 vdd.n2991 52.4337
R17274 vdd.n368 vdd.n367 52.4337
R17275 vdd.n2983 vdd.n372 52.4337
R17276 vdd.n2981 vdd.n2980 52.4337
R17277 vdd.n2976 vdd.n378 52.4337
R17278 vdd.n2974 vdd.n2973 52.4337
R17279 vdd.n2969 vdd.n385 52.4337
R17280 vdd.n2967 vdd.n2966 52.4337
R17281 vdd.n2962 vdd.n392 52.4337
R17282 vdd.n2960 vdd.n2959 52.4337
R17283 vdd.n2955 vdd.n399 52.4337
R17284 vdd.n2953 vdd.n2952 52.4337
R17285 vdd.n408 vdd.n407 52.4337
R17286 vdd.n2944 vdd.n412 52.4337
R17287 vdd.n2942 vdd.n2941 52.4337
R17288 vdd.n2937 vdd.n418 52.4337
R17289 vdd.n2935 vdd.n2934 52.4337
R17290 vdd.n2930 vdd.n425 52.4337
R17291 vdd.n2928 vdd.n2927 52.4337
R17292 vdd.n2923 vdd.n432 52.4337
R17293 vdd.n2921 vdd.n2920 52.4337
R17294 vdd.n2916 vdd.n439 52.4337
R17295 vdd.n2914 vdd.n2913 52.4337
R17296 vdd.n2906 vdd.n2905 52.4337
R17297 vdd.n2842 vdd.n2841 52.4337
R17298 vdd.n517 vdd.n485 52.4337
R17299 vdd.n523 vdd.n486 52.4337
R17300 vdd.n2831 vdd.n487 52.4337
R17301 vdd.n2827 vdd.n488 52.4337
R17302 vdd.n2823 vdd.n489 52.4337
R17303 vdd.n2819 vdd.n490 52.4337
R17304 vdd.n2815 vdd.n491 52.4337
R17305 vdd.n2811 vdd.n492 52.4337
R17306 vdd.n2807 vdd.n493 52.4337
R17307 vdd.n2799 vdd.n494 52.4337
R17308 vdd.n2795 vdd.n495 52.4337
R17309 vdd.n2791 vdd.n496 52.4337
R17310 vdd.n2787 vdd.n497 52.4337
R17311 vdd.n2783 vdd.n498 52.4337
R17312 vdd.n2779 vdd.n499 52.4337
R17313 vdd.n2775 vdd.n500 52.4337
R17314 vdd.n2771 vdd.n501 52.4337
R17315 vdd.n2767 vdd.n502 52.4337
R17316 vdd.n2763 vdd.n503 52.4337
R17317 vdd.n2759 vdd.n504 52.4337
R17318 vdd.n2753 vdd.n505 52.4337
R17319 vdd.n2749 vdd.n506 52.4337
R17320 vdd.n2745 vdd.n507 52.4337
R17321 vdd.n2741 vdd.n508 52.4337
R17322 vdd.n2737 vdd.n509 52.4337
R17323 vdd.n2733 vdd.n510 52.4337
R17324 vdd.n2729 vdd.n511 52.4337
R17325 vdd.n2725 vdd.n512 52.4337
R17326 vdd.n2721 vdd.n513 52.4337
R17327 vdd.n2717 vdd.n514 52.4337
R17328 vdd.n1936 vdd.n1516 52.4337
R17329 vdd.n1934 vdd.n1933 52.4337
R17330 vdd.n1523 vdd.n1522 52.4337
R17331 vdd.n1712 vdd.n1711 52.4337
R17332 vdd.n1709 vdd.n1708 52.4337
R17333 vdd.n1704 vdd.n1531 52.4337
R17334 vdd.n1702 vdd.n1701 52.4337
R17335 vdd.n1697 vdd.n1538 52.4337
R17336 vdd.n1695 vdd.n1694 52.4337
R17337 vdd.n1547 vdd.n1546 52.4337
R17338 vdd.n1686 vdd.n1551 52.4337
R17339 vdd.n1684 vdd.n1683 52.4337
R17340 vdd.n1679 vdd.n1557 52.4337
R17341 vdd.n1677 vdd.n1676 52.4337
R17342 vdd.n1672 vdd.n1564 52.4337
R17343 vdd.n1670 vdd.n1669 52.4337
R17344 vdd.n1665 vdd.n1571 52.4337
R17345 vdd.n1663 vdd.n1662 52.4337
R17346 vdd.n1658 vdd.n1578 52.4337
R17347 vdd.n1656 vdd.n1655 52.4337
R17348 vdd.n1587 vdd.n1586 52.4337
R17349 vdd.n1647 vdd.n1591 52.4337
R17350 vdd.n1645 vdd.n1644 52.4337
R17351 vdd.n1640 vdd.n1597 52.4337
R17352 vdd.n1638 vdd.n1637 52.4337
R17353 vdd.n1633 vdd.n1604 52.4337
R17354 vdd.n1631 vdd.n1630 52.4337
R17355 vdd.n1626 vdd.n1612 52.4337
R17356 vdd.n1624 vdd.n1623 52.4337
R17357 vdd.n1619 vdd.n1618 52.4337
R17358 vdd.n1614 vdd.n1613 52.4337
R17359 vdd.n1945 vdd.n860 52.4337
R17360 vdd.n1423 vdd.n1422 52.4337
R17361 vdd.n1229 vdd.n1197 52.4337
R17362 vdd.n1233 vdd.n1198 52.4337
R17363 vdd.n1235 vdd.n1199 52.4337
R17364 vdd.n1239 vdd.n1200 52.4337
R17365 vdd.n1241 vdd.n1201 52.4337
R17366 vdd.n1245 vdd.n1202 52.4337
R17367 vdd.n1247 vdd.n1203 52.4337
R17368 vdd.n1251 vdd.n1204 52.4337
R17369 vdd.n1253 vdd.n1205 52.4337
R17370 vdd.n1259 vdd.n1206 52.4337
R17371 vdd.n1261 vdd.n1207 52.4337
R17372 vdd.n1265 vdd.n1208 52.4337
R17373 vdd.n1267 vdd.n1209 52.4337
R17374 vdd.n1271 vdd.n1210 52.4337
R17375 vdd.n1273 vdd.n1211 52.4337
R17376 vdd.n1277 vdd.n1212 52.4337
R17377 vdd.n1279 vdd.n1213 52.4337
R17378 vdd.n1283 vdd.n1214 52.4337
R17379 vdd.n1285 vdd.n1215 52.4337
R17380 vdd.n1357 vdd.n1216 52.4337
R17381 vdd.n1290 vdd.n1217 52.4337
R17382 vdd.n1294 vdd.n1218 52.4337
R17383 vdd.n1296 vdd.n1219 52.4337
R17384 vdd.n1300 vdd.n1220 52.4337
R17385 vdd.n1302 vdd.n1221 52.4337
R17386 vdd.n1306 vdd.n1222 52.4337
R17387 vdd.n1308 vdd.n1223 52.4337
R17388 vdd.n1312 vdd.n1224 52.4337
R17389 vdd.n1314 vdd.n1225 52.4337
R17390 vdd.n1318 vdd.n1226 52.4337
R17391 vdd.n1422 vdd.n1196 52.4337
R17392 vdd.n1232 vdd.n1197 52.4337
R17393 vdd.n1234 vdd.n1198 52.4337
R17394 vdd.n1238 vdd.n1199 52.4337
R17395 vdd.n1240 vdd.n1200 52.4337
R17396 vdd.n1244 vdd.n1201 52.4337
R17397 vdd.n1246 vdd.n1202 52.4337
R17398 vdd.n1250 vdd.n1203 52.4337
R17399 vdd.n1252 vdd.n1204 52.4337
R17400 vdd.n1258 vdd.n1205 52.4337
R17401 vdd.n1260 vdd.n1206 52.4337
R17402 vdd.n1264 vdd.n1207 52.4337
R17403 vdd.n1266 vdd.n1208 52.4337
R17404 vdd.n1270 vdd.n1209 52.4337
R17405 vdd.n1272 vdd.n1210 52.4337
R17406 vdd.n1276 vdd.n1211 52.4337
R17407 vdd.n1278 vdd.n1212 52.4337
R17408 vdd.n1282 vdd.n1213 52.4337
R17409 vdd.n1284 vdd.n1214 52.4337
R17410 vdd.n1288 vdd.n1215 52.4337
R17411 vdd.n1289 vdd.n1216 52.4337
R17412 vdd.n1293 vdd.n1217 52.4337
R17413 vdd.n1295 vdd.n1218 52.4337
R17414 vdd.n1299 vdd.n1219 52.4337
R17415 vdd.n1301 vdd.n1220 52.4337
R17416 vdd.n1305 vdd.n1221 52.4337
R17417 vdd.n1307 vdd.n1222 52.4337
R17418 vdd.n1311 vdd.n1223 52.4337
R17419 vdd.n1313 vdd.n1224 52.4337
R17420 vdd.n1317 vdd.n1225 52.4337
R17421 vdd.n1319 vdd.n1226 52.4337
R17422 vdd.n860 vdd.n859 52.4337
R17423 vdd.n1615 vdd.n1614 52.4337
R17424 vdd.n1620 vdd.n1619 52.4337
R17425 vdd.n1625 vdd.n1624 52.4337
R17426 vdd.n1612 vdd.n1605 52.4337
R17427 vdd.n1632 vdd.n1631 52.4337
R17428 vdd.n1604 vdd.n1598 52.4337
R17429 vdd.n1639 vdd.n1638 52.4337
R17430 vdd.n1597 vdd.n1592 52.4337
R17431 vdd.n1646 vdd.n1645 52.4337
R17432 vdd.n1591 vdd.n1590 52.4337
R17433 vdd.n1586 vdd.n1579 52.4337
R17434 vdd.n1657 vdd.n1656 52.4337
R17435 vdd.n1578 vdd.n1572 52.4337
R17436 vdd.n1664 vdd.n1663 52.4337
R17437 vdd.n1571 vdd.n1565 52.4337
R17438 vdd.n1671 vdd.n1670 52.4337
R17439 vdd.n1564 vdd.n1558 52.4337
R17440 vdd.n1678 vdd.n1677 52.4337
R17441 vdd.n1557 vdd.n1552 52.4337
R17442 vdd.n1685 vdd.n1684 52.4337
R17443 vdd.n1551 vdd.n1550 52.4337
R17444 vdd.n1546 vdd.n1539 52.4337
R17445 vdd.n1696 vdd.n1695 52.4337
R17446 vdd.n1538 vdd.n1532 52.4337
R17447 vdd.n1703 vdd.n1702 52.4337
R17448 vdd.n1531 vdd.n1525 52.4337
R17449 vdd.n1710 vdd.n1709 52.4337
R17450 vdd.n1713 vdd.n1712 52.4337
R17451 vdd.n1522 vdd.n1517 52.4337
R17452 vdd.n1935 vdd.n1934 52.4337
R17453 vdd.n1516 vdd.n865 52.4337
R17454 vdd.n2841 vdd.n483 52.4337
R17455 vdd.n522 vdd.n485 52.4337
R17456 vdd.n2832 vdd.n486 52.4337
R17457 vdd.n2828 vdd.n487 52.4337
R17458 vdd.n2824 vdd.n488 52.4337
R17459 vdd.n2820 vdd.n489 52.4337
R17460 vdd.n2816 vdd.n490 52.4337
R17461 vdd.n2812 vdd.n491 52.4337
R17462 vdd.n2808 vdd.n492 52.4337
R17463 vdd.n2798 vdd.n493 52.4337
R17464 vdd.n2796 vdd.n494 52.4337
R17465 vdd.n2792 vdd.n495 52.4337
R17466 vdd.n2788 vdd.n496 52.4337
R17467 vdd.n2784 vdd.n497 52.4337
R17468 vdd.n2780 vdd.n498 52.4337
R17469 vdd.n2776 vdd.n499 52.4337
R17470 vdd.n2772 vdd.n500 52.4337
R17471 vdd.n2768 vdd.n501 52.4337
R17472 vdd.n2764 vdd.n502 52.4337
R17473 vdd.n2760 vdd.n503 52.4337
R17474 vdd.n2752 vdd.n504 52.4337
R17475 vdd.n2750 vdd.n505 52.4337
R17476 vdd.n2746 vdd.n506 52.4337
R17477 vdd.n2742 vdd.n507 52.4337
R17478 vdd.n2738 vdd.n508 52.4337
R17479 vdd.n2734 vdd.n509 52.4337
R17480 vdd.n2730 vdd.n510 52.4337
R17481 vdd.n2726 vdd.n511 52.4337
R17482 vdd.n2722 vdd.n512 52.4337
R17483 vdd.n2718 vdd.n513 52.4337
R17484 vdd.n2714 vdd.n514 52.4337
R17485 vdd.n2905 vdd.n440 52.4337
R17486 vdd.n2915 vdd.n2914 52.4337
R17487 vdd.n439 vdd.n433 52.4337
R17488 vdd.n2922 vdd.n2921 52.4337
R17489 vdd.n432 vdd.n426 52.4337
R17490 vdd.n2929 vdd.n2928 52.4337
R17491 vdd.n425 vdd.n419 52.4337
R17492 vdd.n2936 vdd.n2935 52.4337
R17493 vdd.n418 vdd.n413 52.4337
R17494 vdd.n2943 vdd.n2942 52.4337
R17495 vdd.n412 vdd.n411 52.4337
R17496 vdd.n407 vdd.n400 52.4337
R17497 vdd.n2954 vdd.n2953 52.4337
R17498 vdd.n399 vdd.n393 52.4337
R17499 vdd.n2961 vdd.n2960 52.4337
R17500 vdd.n392 vdd.n386 52.4337
R17501 vdd.n2968 vdd.n2967 52.4337
R17502 vdd.n385 vdd.n379 52.4337
R17503 vdd.n2975 vdd.n2974 52.4337
R17504 vdd.n378 vdd.n373 52.4337
R17505 vdd.n2982 vdd.n2981 52.4337
R17506 vdd.n372 vdd.n371 52.4337
R17507 vdd.n367 vdd.n360 52.4337
R17508 vdd.n2993 vdd.n2992 52.4337
R17509 vdd.n359 vdd.n353 52.4337
R17510 vdd.n3000 vdd.n2999 52.4337
R17511 vdd.n352 vdd.n346 52.4337
R17512 vdd.n3007 vdd.n3006 52.4337
R17513 vdd.n345 vdd.n338 52.4337
R17514 vdd.n3014 vdd.n3013 52.4337
R17515 vdd.n3017 vdd.n3016 52.4337
R17516 vdd.n333 vdd.n330 52.4337
R17517 vdd.t98 vdd.t192 51.4683
R17518 vdd.n250 vdd.n248 42.0461
R17519 vdd.n160 vdd.n158 42.0461
R17520 vdd.n71 vdd.n69 42.0461
R17521 vdd.n1112 vdd.n1110 42.0461
R17522 vdd.n1022 vdd.n1020 42.0461
R17523 vdd.n933 vdd.n931 42.0461
R17524 vdd.n296 vdd.n295 41.6884
R17525 vdd.n206 vdd.n205 41.6884
R17526 vdd.n117 vdd.n116 41.6884
R17527 vdd.n1158 vdd.n1157 41.6884
R17528 vdd.n1068 vdd.n1067 41.6884
R17529 vdd.n979 vdd.n978 41.6884
R17530 vdd.n1322 vdd.n1321 41.1157
R17531 vdd.n1360 vdd.n1359 41.1157
R17532 vdd.n1256 vdd.n1255 41.1157
R17533 vdd.n2910 vdd.n2909 41.1157
R17534 vdd.n2949 vdd.n406 41.1157
R17535 vdd.n2988 vdd.n366 41.1157
R17536 vdd.n2667 vdd.n2666 39.2114
R17537 vdd.n2664 vdd.n2663 39.2114
R17538 vdd.n2659 vdd.n605 39.2114
R17539 vdd.n2657 vdd.n2656 39.2114
R17540 vdd.n2652 vdd.n608 39.2114
R17541 vdd.n2650 vdd.n2649 39.2114
R17542 vdd.n2645 vdd.n611 39.2114
R17543 vdd.n2643 vdd.n2642 39.2114
R17544 vdd.n2639 vdd.n2638 39.2114
R17545 vdd.n2634 vdd.n614 39.2114
R17546 vdd.n2632 vdd.n2631 39.2114
R17547 vdd.n2627 vdd.n617 39.2114
R17548 vdd.n2625 vdd.n2624 39.2114
R17549 vdd.n2620 vdd.n620 39.2114
R17550 vdd.n2618 vdd.n2617 39.2114
R17551 vdd.n2612 vdd.n625 39.2114
R17552 vdd.n2610 vdd.n2609 39.2114
R17553 vdd.n2470 vdd.n703 39.2114
R17554 vdd.n2465 vdd.n2219 39.2114
R17555 vdd.n2462 vdd.n2220 39.2114
R17556 vdd.n2458 vdd.n2221 39.2114
R17557 vdd.n2454 vdd.n2222 39.2114
R17558 vdd.n2450 vdd.n2223 39.2114
R17559 vdd.n2446 vdd.n2224 39.2114
R17560 vdd.n2442 vdd.n2225 39.2114
R17561 vdd.n2438 vdd.n2226 39.2114
R17562 vdd.n2434 vdd.n2227 39.2114
R17563 vdd.n2430 vdd.n2228 39.2114
R17564 vdd.n2426 vdd.n2229 39.2114
R17565 vdd.n2422 vdd.n2230 39.2114
R17566 vdd.n2418 vdd.n2231 39.2114
R17567 vdd.n2414 vdd.n2232 39.2114
R17568 vdd.n2410 vdd.n2233 39.2114
R17569 vdd.n2405 vdd.n2234 39.2114
R17570 vdd.n2213 vdd.n743 39.2114
R17571 vdd.n2209 vdd.n742 39.2114
R17572 vdd.n2205 vdd.n741 39.2114
R17573 vdd.n2201 vdd.n740 39.2114
R17574 vdd.n2197 vdd.n739 39.2114
R17575 vdd.n2193 vdd.n738 39.2114
R17576 vdd.n2189 vdd.n737 39.2114
R17577 vdd.n2185 vdd.n736 39.2114
R17578 vdd.n2181 vdd.n735 39.2114
R17579 vdd.n2177 vdd.n734 39.2114
R17580 vdd.n2173 vdd.n733 39.2114
R17581 vdd.n2169 vdd.n732 39.2114
R17582 vdd.n2165 vdd.n731 39.2114
R17583 vdd.n2161 vdd.n730 39.2114
R17584 vdd.n2157 vdd.n729 39.2114
R17585 vdd.n2152 vdd.n728 39.2114
R17586 vdd.n2148 vdd.n727 39.2114
R17587 vdd.n1724 vdd.n838 39.2114
R17588 vdd.n1730 vdd.n1729 39.2114
R17589 vdd.n1733 vdd.n1732 39.2114
R17590 vdd.n1738 vdd.n1737 39.2114
R17591 vdd.n1741 vdd.n1740 39.2114
R17592 vdd.n1746 vdd.n1745 39.2114
R17593 vdd.n1749 vdd.n1748 39.2114
R17594 vdd.n1754 vdd.n1753 39.2114
R17595 vdd.n1925 vdd.n1756 39.2114
R17596 vdd.n1924 vdd.n1923 39.2114
R17597 vdd.n1917 vdd.n1758 39.2114
R17598 vdd.n1916 vdd.n1915 39.2114
R17599 vdd.n1909 vdd.n1760 39.2114
R17600 vdd.n1908 vdd.n1907 39.2114
R17601 vdd.n1901 vdd.n1762 39.2114
R17602 vdd.n1900 vdd.n1899 39.2114
R17603 vdd.n1893 vdd.n1764 39.2114
R17604 vdd.n2586 vdd.n2585 39.2114
R17605 vdd.n2581 vdd.n2553 39.2114
R17606 vdd.n2579 vdd.n2578 39.2114
R17607 vdd.n2574 vdd.n2556 39.2114
R17608 vdd.n2572 vdd.n2571 39.2114
R17609 vdd.n2567 vdd.n2559 39.2114
R17610 vdd.n2565 vdd.n2564 39.2114
R17611 vdd.n2560 vdd.n577 39.2114
R17612 vdd.n2704 vdd.n2703 39.2114
R17613 vdd.n2701 vdd.n2700 39.2114
R17614 vdd.n2696 vdd.n581 39.2114
R17615 vdd.n2694 vdd.n2693 39.2114
R17616 vdd.n2689 vdd.n584 39.2114
R17617 vdd.n2687 vdd.n2686 39.2114
R17618 vdd.n2682 vdd.n587 39.2114
R17619 vdd.n2680 vdd.n2679 39.2114
R17620 vdd.n2675 vdd.n593 39.2114
R17621 vdd.n2472 vdd.n706 39.2114
R17622 vdd.n2235 vdd.n708 39.2114
R17623 vdd.n2261 vdd.n2236 39.2114
R17624 vdd.n2265 vdd.n2237 39.2114
R17625 vdd.n2269 vdd.n2238 39.2114
R17626 vdd.n2273 vdd.n2239 39.2114
R17627 vdd.n2277 vdd.n2240 39.2114
R17628 vdd.n2281 vdd.n2241 39.2114
R17629 vdd.n2285 vdd.n2242 39.2114
R17630 vdd.n2289 vdd.n2243 39.2114
R17631 vdd.n2293 vdd.n2244 39.2114
R17632 vdd.n2297 vdd.n2245 39.2114
R17633 vdd.n2301 vdd.n2246 39.2114
R17634 vdd.n2305 vdd.n2247 39.2114
R17635 vdd.n2309 vdd.n2248 39.2114
R17636 vdd.n2313 vdd.n2249 39.2114
R17637 vdd.n2317 vdd.n2250 39.2114
R17638 vdd.n2473 vdd.n2472 39.2114
R17639 vdd.n2260 vdd.n2235 39.2114
R17640 vdd.n2264 vdd.n2236 39.2114
R17641 vdd.n2268 vdd.n2237 39.2114
R17642 vdd.n2272 vdd.n2238 39.2114
R17643 vdd.n2276 vdd.n2239 39.2114
R17644 vdd.n2280 vdd.n2240 39.2114
R17645 vdd.n2284 vdd.n2241 39.2114
R17646 vdd.n2288 vdd.n2242 39.2114
R17647 vdd.n2292 vdd.n2243 39.2114
R17648 vdd.n2296 vdd.n2244 39.2114
R17649 vdd.n2300 vdd.n2245 39.2114
R17650 vdd.n2304 vdd.n2246 39.2114
R17651 vdd.n2308 vdd.n2247 39.2114
R17652 vdd.n2312 vdd.n2248 39.2114
R17653 vdd.n2316 vdd.n2249 39.2114
R17654 vdd.n2319 vdd.n2250 39.2114
R17655 vdd.n593 vdd.n588 39.2114
R17656 vdd.n2681 vdd.n2680 39.2114
R17657 vdd.n587 vdd.n585 39.2114
R17658 vdd.n2688 vdd.n2687 39.2114
R17659 vdd.n584 vdd.n582 39.2114
R17660 vdd.n2695 vdd.n2694 39.2114
R17661 vdd.n581 vdd.n579 39.2114
R17662 vdd.n2702 vdd.n2701 39.2114
R17663 vdd.n2705 vdd.n2704 39.2114
R17664 vdd.n2561 vdd.n2560 39.2114
R17665 vdd.n2566 vdd.n2565 39.2114
R17666 vdd.n2559 vdd.n2557 39.2114
R17667 vdd.n2573 vdd.n2572 39.2114
R17668 vdd.n2556 vdd.n2554 39.2114
R17669 vdd.n2580 vdd.n2579 39.2114
R17670 vdd.n2553 vdd.n2551 39.2114
R17671 vdd.n2587 vdd.n2586 39.2114
R17672 vdd.n1725 vdd.n1724 39.2114
R17673 vdd.n1731 vdd.n1730 39.2114
R17674 vdd.n1732 vdd.n1721 39.2114
R17675 vdd.n1739 vdd.n1738 39.2114
R17676 vdd.n1740 vdd.n1719 39.2114
R17677 vdd.n1747 vdd.n1746 39.2114
R17678 vdd.n1748 vdd.n1717 39.2114
R17679 vdd.n1755 vdd.n1754 39.2114
R17680 vdd.n1926 vdd.n1925 39.2114
R17681 vdd.n1923 vdd.n1922 39.2114
R17682 vdd.n1918 vdd.n1917 39.2114
R17683 vdd.n1915 vdd.n1914 39.2114
R17684 vdd.n1910 vdd.n1909 39.2114
R17685 vdd.n1907 vdd.n1906 39.2114
R17686 vdd.n1902 vdd.n1901 39.2114
R17687 vdd.n1899 vdd.n1898 39.2114
R17688 vdd.n1894 vdd.n1893 39.2114
R17689 vdd.n2151 vdd.n727 39.2114
R17690 vdd.n2156 vdd.n728 39.2114
R17691 vdd.n2160 vdd.n729 39.2114
R17692 vdd.n2164 vdd.n730 39.2114
R17693 vdd.n2168 vdd.n731 39.2114
R17694 vdd.n2172 vdd.n732 39.2114
R17695 vdd.n2176 vdd.n733 39.2114
R17696 vdd.n2180 vdd.n734 39.2114
R17697 vdd.n2184 vdd.n735 39.2114
R17698 vdd.n2188 vdd.n736 39.2114
R17699 vdd.n2192 vdd.n737 39.2114
R17700 vdd.n2196 vdd.n738 39.2114
R17701 vdd.n2200 vdd.n739 39.2114
R17702 vdd.n2204 vdd.n740 39.2114
R17703 vdd.n2208 vdd.n741 39.2114
R17704 vdd.n2212 vdd.n742 39.2114
R17705 vdd.n745 vdd.n743 39.2114
R17706 vdd.n2470 vdd.n2469 39.2114
R17707 vdd.n2463 vdd.n2219 39.2114
R17708 vdd.n2459 vdd.n2220 39.2114
R17709 vdd.n2455 vdd.n2221 39.2114
R17710 vdd.n2451 vdd.n2222 39.2114
R17711 vdd.n2447 vdd.n2223 39.2114
R17712 vdd.n2443 vdd.n2224 39.2114
R17713 vdd.n2439 vdd.n2225 39.2114
R17714 vdd.n2435 vdd.n2226 39.2114
R17715 vdd.n2431 vdd.n2227 39.2114
R17716 vdd.n2427 vdd.n2228 39.2114
R17717 vdd.n2423 vdd.n2229 39.2114
R17718 vdd.n2419 vdd.n2230 39.2114
R17719 vdd.n2415 vdd.n2231 39.2114
R17720 vdd.n2411 vdd.n2232 39.2114
R17721 vdd.n2406 vdd.n2233 39.2114
R17722 vdd.n2402 vdd.n2234 39.2114
R17723 vdd.n2611 vdd.n2610 39.2114
R17724 vdd.n625 vdd.n621 39.2114
R17725 vdd.n2619 vdd.n2618 39.2114
R17726 vdd.n620 vdd.n618 39.2114
R17727 vdd.n2626 vdd.n2625 39.2114
R17728 vdd.n617 vdd.n615 39.2114
R17729 vdd.n2633 vdd.n2632 39.2114
R17730 vdd.n614 vdd.n612 39.2114
R17731 vdd.n2640 vdd.n2639 39.2114
R17732 vdd.n2644 vdd.n2643 39.2114
R17733 vdd.n611 vdd.n609 39.2114
R17734 vdd.n2651 vdd.n2650 39.2114
R17735 vdd.n608 vdd.n606 39.2114
R17736 vdd.n2658 vdd.n2657 39.2114
R17737 vdd.n605 vdd.n603 39.2114
R17738 vdd.n2665 vdd.n2664 39.2114
R17739 vdd.n2668 vdd.n2667 39.2114
R17740 vdd.n753 vdd.n709 39.2114
R17741 vdd.n2140 vdd.n710 39.2114
R17742 vdd.n2136 vdd.n711 39.2114
R17743 vdd.n2132 vdd.n712 39.2114
R17744 vdd.n2128 vdd.n713 39.2114
R17745 vdd.n2124 vdd.n714 39.2114
R17746 vdd.n2120 vdd.n715 39.2114
R17747 vdd.n2116 vdd.n716 39.2114
R17748 vdd.n2112 vdd.n717 39.2114
R17749 vdd.n2108 vdd.n718 39.2114
R17750 vdd.n2104 vdd.n719 39.2114
R17751 vdd.n2100 vdd.n720 39.2114
R17752 vdd.n2096 vdd.n721 39.2114
R17753 vdd.n2092 vdd.n722 39.2114
R17754 vdd.n2088 vdd.n723 39.2114
R17755 vdd.n2084 vdd.n724 39.2114
R17756 vdd.n2080 vdd.n725 39.2114
R17757 vdd.n1983 vdd.n842 39.2114
R17758 vdd.n1982 vdd.n1981 39.2114
R17759 vdd.n1975 vdd.n844 39.2114
R17760 vdd.n1974 vdd.n1973 39.2114
R17761 vdd.n1967 vdd.n846 39.2114
R17762 vdd.n1966 vdd.n1965 39.2114
R17763 vdd.n1959 vdd.n848 39.2114
R17764 vdd.n1958 vdd.n1957 39.2114
R17765 vdd.n851 vdd.n850 39.2114
R17766 vdd.n1799 vdd.n1798 39.2114
R17767 vdd.n1804 vdd.n1803 39.2114
R17768 vdd.n1807 vdd.n1806 39.2114
R17769 vdd.n1812 vdd.n1811 39.2114
R17770 vdd.n1815 vdd.n1814 39.2114
R17771 vdd.n1820 vdd.n1819 39.2114
R17772 vdd.n1823 vdd.n1822 39.2114
R17773 vdd.n1829 vdd.n1828 39.2114
R17774 vdd.n2077 vdd.n725 39.2114
R17775 vdd.n2081 vdd.n724 39.2114
R17776 vdd.n2085 vdd.n723 39.2114
R17777 vdd.n2089 vdd.n722 39.2114
R17778 vdd.n2093 vdd.n721 39.2114
R17779 vdd.n2097 vdd.n720 39.2114
R17780 vdd.n2101 vdd.n719 39.2114
R17781 vdd.n2105 vdd.n718 39.2114
R17782 vdd.n2109 vdd.n717 39.2114
R17783 vdd.n2113 vdd.n716 39.2114
R17784 vdd.n2117 vdd.n715 39.2114
R17785 vdd.n2121 vdd.n714 39.2114
R17786 vdd.n2125 vdd.n713 39.2114
R17787 vdd.n2129 vdd.n712 39.2114
R17788 vdd.n2133 vdd.n711 39.2114
R17789 vdd.n2137 vdd.n710 39.2114
R17790 vdd.n2141 vdd.n709 39.2114
R17791 vdd.n1984 vdd.n1983 39.2114
R17792 vdd.n1981 vdd.n1980 39.2114
R17793 vdd.n1976 vdd.n1975 39.2114
R17794 vdd.n1973 vdd.n1972 39.2114
R17795 vdd.n1968 vdd.n1967 39.2114
R17796 vdd.n1965 vdd.n1964 39.2114
R17797 vdd.n1960 vdd.n1959 39.2114
R17798 vdd.n1957 vdd.n1956 39.2114
R17799 vdd.n852 vdd.n851 39.2114
R17800 vdd.n1800 vdd.n1799 39.2114
R17801 vdd.n1805 vdd.n1804 39.2114
R17802 vdd.n1806 vdd.n1796 39.2114
R17803 vdd.n1813 vdd.n1812 39.2114
R17804 vdd.n1814 vdd.n1794 39.2114
R17805 vdd.n1821 vdd.n1820 39.2114
R17806 vdd.n1822 vdd.n1790 39.2114
R17807 vdd.n1830 vdd.n1829 39.2114
R17808 vdd.n1949 vdd.n1948 37.2369
R17809 vdd.n1652 vdd.n1585 37.2369
R17810 vdd.n1691 vdd.n1545 37.2369
R17811 vdd.n2758 vdd.n558 37.2369
R17812 vdd.n2806 vdd.n2805 37.2369
R17813 vdd.n2713 vdd.n2712 37.2369
R17814 vdd.n1991 vdd.n837 31.6883
R17815 vdd.n2216 vdd.n746 31.6883
R17816 vdd.n2149 vdd.n749 31.6883
R17817 vdd.n1895 vdd.n1892 31.6883
R17818 vdd.n2403 vdd.n2401 31.6883
R17819 vdd.n2608 vdd.n2607 31.6883
R17820 vdd.n2480 vdd.n702 31.6883
R17821 vdd.n2671 vdd.n2670 31.6883
R17822 vdd.n2590 vdd.n2589 31.6883
R17823 vdd.n2676 vdd.n592 31.6883
R17824 vdd.n2322 vdd.n2321 31.6883
R17825 vdd.n2476 vdd.n2475 31.6883
R17826 vdd.n1987 vdd.n1986 31.6883
R17827 vdd.n2144 vdd.n2143 31.6883
R17828 vdd.n2076 vdd.n2075 31.6883
R17829 vdd.n1833 vdd.n1832 31.6883
R17830 vdd.n1826 vdd.n1792 30.449
R17831 vdd.n757 vdd.n756 30.449
R17832 vdd.n1767 vdd.n1766 30.449
R17833 vdd.n2154 vdd.n748 30.449
R17834 vdd.n2258 vdd.n2257 30.449
R17835 vdd.n2614 vdd.n623 30.449
R17836 vdd.n2408 vdd.n2254 30.449
R17837 vdd.n591 vdd.n590 30.449
R17838 vdd.n1421 vdd.n1228 22.6735
R17839 vdd.n1943 vdd.n863 22.6735
R17840 vdd.n2840 vdd.n516 22.6735
R17841 vdd.n3025 vdd.n329 22.6735
R17842 vdd.n1432 vdd.n1190 19.3944
R17843 vdd.n1432 vdd.n1188 19.3944
R17844 vdd.n1436 vdd.n1188 19.3944
R17845 vdd.n1436 vdd.n1178 19.3944
R17846 vdd.n1449 vdd.n1178 19.3944
R17847 vdd.n1449 vdd.n1176 19.3944
R17848 vdd.n1453 vdd.n1176 19.3944
R17849 vdd.n1453 vdd.n1168 19.3944
R17850 vdd.n1467 vdd.n1168 19.3944
R17851 vdd.n1467 vdd.n1166 19.3944
R17852 vdd.n1471 vdd.n1166 19.3944
R17853 vdd.n1471 vdd.n885 19.3944
R17854 vdd.n1483 vdd.n885 19.3944
R17855 vdd.n1483 vdd.n883 19.3944
R17856 vdd.n1487 vdd.n883 19.3944
R17857 vdd.n1487 vdd.n875 19.3944
R17858 vdd.n1500 vdd.n875 19.3944
R17859 vdd.n1500 vdd.n872 19.3944
R17860 vdd.n1506 vdd.n872 19.3944
R17861 vdd.n1506 vdd.n873 19.3944
R17862 vdd.n873 vdd.n862 19.3944
R17863 vdd.n1356 vdd.n1291 19.3944
R17864 vdd.n1352 vdd.n1291 19.3944
R17865 vdd.n1352 vdd.n1351 19.3944
R17866 vdd.n1351 vdd.n1350 19.3944
R17867 vdd.n1350 vdd.n1297 19.3944
R17868 vdd.n1346 vdd.n1297 19.3944
R17869 vdd.n1346 vdd.n1345 19.3944
R17870 vdd.n1345 vdd.n1344 19.3944
R17871 vdd.n1344 vdd.n1303 19.3944
R17872 vdd.n1340 vdd.n1303 19.3944
R17873 vdd.n1340 vdd.n1339 19.3944
R17874 vdd.n1339 vdd.n1338 19.3944
R17875 vdd.n1338 vdd.n1309 19.3944
R17876 vdd.n1334 vdd.n1309 19.3944
R17877 vdd.n1334 vdd.n1333 19.3944
R17878 vdd.n1333 vdd.n1332 19.3944
R17879 vdd.n1332 vdd.n1315 19.3944
R17880 vdd.n1328 vdd.n1315 19.3944
R17881 vdd.n1328 vdd.n1327 19.3944
R17882 vdd.n1327 vdd.n1326 19.3944
R17883 vdd.n1391 vdd.n1390 19.3944
R17884 vdd.n1390 vdd.n1389 19.3944
R17885 vdd.n1389 vdd.n1262 19.3944
R17886 vdd.n1385 vdd.n1262 19.3944
R17887 vdd.n1385 vdd.n1384 19.3944
R17888 vdd.n1384 vdd.n1383 19.3944
R17889 vdd.n1383 vdd.n1268 19.3944
R17890 vdd.n1379 vdd.n1268 19.3944
R17891 vdd.n1379 vdd.n1378 19.3944
R17892 vdd.n1378 vdd.n1377 19.3944
R17893 vdd.n1377 vdd.n1274 19.3944
R17894 vdd.n1373 vdd.n1274 19.3944
R17895 vdd.n1373 vdd.n1372 19.3944
R17896 vdd.n1372 vdd.n1371 19.3944
R17897 vdd.n1371 vdd.n1280 19.3944
R17898 vdd.n1367 vdd.n1280 19.3944
R17899 vdd.n1367 vdd.n1366 19.3944
R17900 vdd.n1366 vdd.n1365 19.3944
R17901 vdd.n1365 vdd.n1286 19.3944
R17902 vdd.n1361 vdd.n1286 19.3944
R17903 vdd.n1424 vdd.n1195 19.3944
R17904 vdd.n1419 vdd.n1195 19.3944
R17905 vdd.n1419 vdd.n1230 19.3944
R17906 vdd.n1415 vdd.n1230 19.3944
R17907 vdd.n1415 vdd.n1414 19.3944
R17908 vdd.n1414 vdd.n1413 19.3944
R17909 vdd.n1413 vdd.n1236 19.3944
R17910 vdd.n1409 vdd.n1236 19.3944
R17911 vdd.n1409 vdd.n1408 19.3944
R17912 vdd.n1408 vdd.n1407 19.3944
R17913 vdd.n1407 vdd.n1242 19.3944
R17914 vdd.n1403 vdd.n1242 19.3944
R17915 vdd.n1403 vdd.n1402 19.3944
R17916 vdd.n1402 vdd.n1401 19.3944
R17917 vdd.n1401 vdd.n1248 19.3944
R17918 vdd.n1397 vdd.n1248 19.3944
R17919 vdd.n1397 vdd.n1396 19.3944
R17920 vdd.n1396 vdd.n1395 19.3944
R17921 vdd.n1648 vdd.n1583 19.3944
R17922 vdd.n1648 vdd.n1589 19.3944
R17923 vdd.n1643 vdd.n1589 19.3944
R17924 vdd.n1643 vdd.n1642 19.3944
R17925 vdd.n1642 vdd.n1641 19.3944
R17926 vdd.n1641 vdd.n1596 19.3944
R17927 vdd.n1636 vdd.n1596 19.3944
R17928 vdd.n1636 vdd.n1635 19.3944
R17929 vdd.n1635 vdd.n1634 19.3944
R17930 vdd.n1634 vdd.n1603 19.3944
R17931 vdd.n1629 vdd.n1603 19.3944
R17932 vdd.n1629 vdd.n1628 19.3944
R17933 vdd.n1628 vdd.n1627 19.3944
R17934 vdd.n1627 vdd.n1611 19.3944
R17935 vdd.n1622 vdd.n1611 19.3944
R17936 vdd.n1622 vdd.n1621 19.3944
R17937 vdd.n1617 vdd.n1616 19.3944
R17938 vdd.n1950 vdd.n858 19.3944
R17939 vdd.n1687 vdd.n1543 19.3944
R17940 vdd.n1687 vdd.n1549 19.3944
R17941 vdd.n1682 vdd.n1549 19.3944
R17942 vdd.n1682 vdd.n1681 19.3944
R17943 vdd.n1681 vdd.n1680 19.3944
R17944 vdd.n1680 vdd.n1556 19.3944
R17945 vdd.n1675 vdd.n1556 19.3944
R17946 vdd.n1675 vdd.n1674 19.3944
R17947 vdd.n1674 vdd.n1673 19.3944
R17948 vdd.n1673 vdd.n1563 19.3944
R17949 vdd.n1668 vdd.n1563 19.3944
R17950 vdd.n1668 vdd.n1667 19.3944
R17951 vdd.n1667 vdd.n1666 19.3944
R17952 vdd.n1666 vdd.n1570 19.3944
R17953 vdd.n1661 vdd.n1570 19.3944
R17954 vdd.n1661 vdd.n1660 19.3944
R17955 vdd.n1660 vdd.n1659 19.3944
R17956 vdd.n1659 vdd.n1577 19.3944
R17957 vdd.n1654 vdd.n1577 19.3944
R17958 vdd.n1654 vdd.n1653 19.3944
R17959 vdd.n1938 vdd.n1937 19.3944
R17960 vdd.n1937 vdd.n1515 19.3944
R17961 vdd.n1932 vdd.n1931 19.3944
R17962 vdd.n1714 vdd.n1519 19.3944
R17963 vdd.n1714 vdd.n1521 19.3944
R17964 vdd.n1524 vdd.n1521 19.3944
R17965 vdd.n1707 vdd.n1524 19.3944
R17966 vdd.n1707 vdd.n1706 19.3944
R17967 vdd.n1706 vdd.n1705 19.3944
R17968 vdd.n1705 vdd.n1530 19.3944
R17969 vdd.n1700 vdd.n1530 19.3944
R17970 vdd.n1700 vdd.n1699 19.3944
R17971 vdd.n1699 vdd.n1698 19.3944
R17972 vdd.n1698 vdd.n1537 19.3944
R17973 vdd.n1693 vdd.n1537 19.3944
R17974 vdd.n1693 vdd.n1692 19.3944
R17975 vdd.n1428 vdd.n1193 19.3944
R17976 vdd.n1428 vdd.n1184 19.3944
R17977 vdd.n1441 vdd.n1184 19.3944
R17978 vdd.n1441 vdd.n1182 19.3944
R17979 vdd.n1445 vdd.n1182 19.3944
R17980 vdd.n1445 vdd.n1173 19.3944
R17981 vdd.n1458 vdd.n1173 19.3944
R17982 vdd.n1458 vdd.n1171 19.3944
R17983 vdd.n1463 vdd.n1171 19.3944
R17984 vdd.n1463 vdd.n1162 19.3944
R17985 vdd.n1475 vdd.n1162 19.3944
R17986 vdd.n1475 vdd.n890 19.3944
R17987 vdd.n1479 vdd.n890 19.3944
R17988 vdd.n1479 vdd.n880 19.3944
R17989 vdd.n1492 vdd.n880 19.3944
R17990 vdd.n1492 vdd.n878 19.3944
R17991 vdd.n1496 vdd.n878 19.3944
R17992 vdd.n1496 vdd.n868 19.3944
R17993 vdd.n1511 vdd.n868 19.3944
R17994 vdd.n1511 vdd.n866 19.3944
R17995 vdd.n1941 vdd.n866 19.3944
R17996 vdd.n2851 vdd.n477 19.3944
R17997 vdd.n2851 vdd.n475 19.3944
R17998 vdd.n2855 vdd.n475 19.3944
R17999 vdd.n2855 vdd.n465 19.3944
R18000 vdd.n2868 vdd.n465 19.3944
R18001 vdd.n2868 vdd.n463 19.3944
R18002 vdd.n2872 vdd.n463 19.3944
R18003 vdd.n2872 vdd.n453 19.3944
R18004 vdd.n2884 vdd.n453 19.3944
R18005 vdd.n2884 vdd.n451 19.3944
R18006 vdd.n2888 vdd.n451 19.3944
R18007 vdd.n2889 vdd.n2888 19.3944
R18008 vdd.n2890 vdd.n2889 19.3944
R18009 vdd.n2890 vdd.n449 19.3944
R18010 vdd.n2894 vdd.n449 19.3944
R18011 vdd.n2895 vdd.n2894 19.3944
R18012 vdd.n2896 vdd.n2895 19.3944
R18013 vdd.n2896 vdd.n446 19.3944
R18014 vdd.n2900 vdd.n446 19.3944
R18015 vdd.n2901 vdd.n2900 19.3944
R18016 vdd.n2902 vdd.n2901 19.3944
R18017 vdd.n2945 vdd.n404 19.3944
R18018 vdd.n2945 vdd.n410 19.3944
R18019 vdd.n2940 vdd.n410 19.3944
R18020 vdd.n2940 vdd.n2939 19.3944
R18021 vdd.n2939 vdd.n2938 19.3944
R18022 vdd.n2938 vdd.n417 19.3944
R18023 vdd.n2933 vdd.n417 19.3944
R18024 vdd.n2933 vdd.n2932 19.3944
R18025 vdd.n2932 vdd.n2931 19.3944
R18026 vdd.n2931 vdd.n424 19.3944
R18027 vdd.n2926 vdd.n424 19.3944
R18028 vdd.n2926 vdd.n2925 19.3944
R18029 vdd.n2925 vdd.n2924 19.3944
R18030 vdd.n2924 vdd.n431 19.3944
R18031 vdd.n2919 vdd.n431 19.3944
R18032 vdd.n2919 vdd.n2918 19.3944
R18033 vdd.n2918 vdd.n2917 19.3944
R18034 vdd.n2917 vdd.n438 19.3944
R18035 vdd.n2912 vdd.n438 19.3944
R18036 vdd.n2912 vdd.n2911 19.3944
R18037 vdd.n2984 vdd.n364 19.3944
R18038 vdd.n2984 vdd.n370 19.3944
R18039 vdd.n2979 vdd.n370 19.3944
R18040 vdd.n2979 vdd.n2978 19.3944
R18041 vdd.n2978 vdd.n2977 19.3944
R18042 vdd.n2977 vdd.n377 19.3944
R18043 vdd.n2972 vdd.n377 19.3944
R18044 vdd.n2972 vdd.n2971 19.3944
R18045 vdd.n2971 vdd.n2970 19.3944
R18046 vdd.n2970 vdd.n384 19.3944
R18047 vdd.n2965 vdd.n384 19.3944
R18048 vdd.n2965 vdd.n2964 19.3944
R18049 vdd.n2964 vdd.n2963 19.3944
R18050 vdd.n2963 vdd.n391 19.3944
R18051 vdd.n2958 vdd.n391 19.3944
R18052 vdd.n2958 vdd.n2957 19.3944
R18053 vdd.n2957 vdd.n2956 19.3944
R18054 vdd.n2956 vdd.n398 19.3944
R18055 vdd.n2951 vdd.n398 19.3944
R18056 vdd.n2951 vdd.n2950 19.3944
R18057 vdd.n3020 vdd.n3019 19.3944
R18058 vdd.n3019 vdd.n3018 19.3944
R18059 vdd.n3018 vdd.n336 19.3944
R18060 vdd.n337 vdd.n336 19.3944
R18061 vdd.n3011 vdd.n337 19.3944
R18062 vdd.n3011 vdd.n3010 19.3944
R18063 vdd.n3010 vdd.n3009 19.3944
R18064 vdd.n3009 vdd.n344 19.3944
R18065 vdd.n3004 vdd.n344 19.3944
R18066 vdd.n3004 vdd.n3003 19.3944
R18067 vdd.n3003 vdd.n3002 19.3944
R18068 vdd.n3002 vdd.n351 19.3944
R18069 vdd.n2997 vdd.n351 19.3944
R18070 vdd.n2997 vdd.n2996 19.3944
R18071 vdd.n2996 vdd.n2995 19.3944
R18072 vdd.n2995 vdd.n358 19.3944
R18073 vdd.n2990 vdd.n358 19.3944
R18074 vdd.n2990 vdd.n2989 19.3944
R18075 vdd.n2847 vdd.n480 19.3944
R18076 vdd.n2847 vdd.n471 19.3944
R18077 vdd.n2860 vdd.n471 19.3944
R18078 vdd.n2860 vdd.n469 19.3944
R18079 vdd.n2864 vdd.n469 19.3944
R18080 vdd.n2864 vdd.n460 19.3944
R18081 vdd.n2876 vdd.n460 19.3944
R18082 vdd.n2876 vdd.n458 19.3944
R18083 vdd.n2880 vdd.n458 19.3944
R18084 vdd.n2880 vdd.n300 19.3944
R18085 vdd.n3045 vdd.n300 19.3944
R18086 vdd.n3045 vdd.n301 19.3944
R18087 vdd.n3039 vdd.n301 19.3944
R18088 vdd.n3039 vdd.n3038 19.3944
R18089 vdd.n3038 vdd.n3037 19.3944
R18090 vdd.n3037 vdd.n313 19.3944
R18091 vdd.n3031 vdd.n313 19.3944
R18092 vdd.n3031 vdd.n3030 19.3944
R18093 vdd.n3030 vdd.n3029 19.3944
R18094 vdd.n3029 vdd.n324 19.3944
R18095 vdd.n3023 vdd.n324 19.3944
R18096 vdd.n2800 vdd.n536 19.3944
R18097 vdd.n2800 vdd.n2797 19.3944
R18098 vdd.n2797 vdd.n2794 19.3944
R18099 vdd.n2794 vdd.n2793 19.3944
R18100 vdd.n2793 vdd.n2790 19.3944
R18101 vdd.n2790 vdd.n2789 19.3944
R18102 vdd.n2789 vdd.n2786 19.3944
R18103 vdd.n2786 vdd.n2785 19.3944
R18104 vdd.n2785 vdd.n2782 19.3944
R18105 vdd.n2782 vdd.n2781 19.3944
R18106 vdd.n2781 vdd.n2778 19.3944
R18107 vdd.n2778 vdd.n2777 19.3944
R18108 vdd.n2777 vdd.n2774 19.3944
R18109 vdd.n2774 vdd.n2773 19.3944
R18110 vdd.n2773 vdd.n2770 19.3944
R18111 vdd.n2770 vdd.n2769 19.3944
R18112 vdd.n2769 vdd.n2766 19.3944
R18113 vdd.n2766 vdd.n2765 19.3944
R18114 vdd.n2765 vdd.n2762 19.3944
R18115 vdd.n2762 vdd.n2761 19.3944
R18116 vdd.n2843 vdd.n482 19.3944
R18117 vdd.n2838 vdd.n482 19.3944
R18118 vdd.n521 vdd.n518 19.3944
R18119 vdd.n2834 vdd.n2833 19.3944
R18120 vdd.n2833 vdd.n2830 19.3944
R18121 vdd.n2830 vdd.n2829 19.3944
R18122 vdd.n2829 vdd.n2826 19.3944
R18123 vdd.n2826 vdd.n2825 19.3944
R18124 vdd.n2825 vdd.n2822 19.3944
R18125 vdd.n2822 vdd.n2821 19.3944
R18126 vdd.n2821 vdd.n2818 19.3944
R18127 vdd.n2818 vdd.n2817 19.3944
R18128 vdd.n2817 vdd.n2814 19.3944
R18129 vdd.n2814 vdd.n2813 19.3944
R18130 vdd.n2813 vdd.n2810 19.3944
R18131 vdd.n2810 vdd.n2809 19.3944
R18132 vdd.n2754 vdd.n556 19.3944
R18133 vdd.n2754 vdd.n2751 19.3944
R18134 vdd.n2751 vdd.n2748 19.3944
R18135 vdd.n2748 vdd.n2747 19.3944
R18136 vdd.n2747 vdd.n2744 19.3944
R18137 vdd.n2744 vdd.n2743 19.3944
R18138 vdd.n2743 vdd.n2740 19.3944
R18139 vdd.n2740 vdd.n2739 19.3944
R18140 vdd.n2739 vdd.n2736 19.3944
R18141 vdd.n2736 vdd.n2735 19.3944
R18142 vdd.n2735 vdd.n2732 19.3944
R18143 vdd.n2732 vdd.n2731 19.3944
R18144 vdd.n2731 vdd.n2728 19.3944
R18145 vdd.n2728 vdd.n2727 19.3944
R18146 vdd.n2727 vdd.n2724 19.3944
R18147 vdd.n2724 vdd.n2723 19.3944
R18148 vdd.n2720 vdd.n2719 19.3944
R18149 vdd.n2716 vdd.n2715 19.3944
R18150 vdd.n1360 vdd.n1356 19.0066
R18151 vdd.n1652 vdd.n1583 19.0066
R18152 vdd.n2949 vdd.n404 19.0066
R18153 vdd.n2758 vdd.n556 19.0066
R18154 vdd.n1792 vdd.n1791 16.0975
R18155 vdd.n756 vdd.n755 16.0975
R18156 vdd.n1321 vdd.n1320 16.0975
R18157 vdd.n1359 vdd.n1358 16.0975
R18158 vdd.n1255 vdd.n1254 16.0975
R18159 vdd.n1948 vdd.n1947 16.0975
R18160 vdd.n1585 vdd.n1584 16.0975
R18161 vdd.n1545 vdd.n1544 16.0975
R18162 vdd.n1766 vdd.n1765 16.0975
R18163 vdd.n748 vdd.n747 16.0975
R18164 vdd.n2257 vdd.n2256 16.0975
R18165 vdd.n2909 vdd.n2908 16.0975
R18166 vdd.n406 vdd.n405 16.0975
R18167 vdd.n366 vdd.n365 16.0975
R18168 vdd.n558 vdd.n557 16.0975
R18169 vdd.n2805 vdd.n2804 16.0975
R18170 vdd.n623 vdd.n622 16.0975
R18171 vdd.n2254 vdd.n2253 16.0975
R18172 vdd.n2712 vdd.n2711 16.0975
R18173 vdd.n590 vdd.n589 16.0975
R18174 vdd.t192 vdd.n2218 15.4182
R18175 vdd.n2471 vdd.t98 15.4182
R18176 vdd.n1989 vdd.n839 14.5112
R18177 vdd.n2673 vdd.n484 14.5112
R18178 vdd.n28 vdd.n27 14.4007
R18179 vdd.n292 vdd.n257 13.1884
R18180 vdd.n245 vdd.n210 13.1884
R18181 vdd.n202 vdd.n167 13.1884
R18182 vdd.n155 vdd.n120 13.1884
R18183 vdd.n113 vdd.n78 13.1884
R18184 vdd.n66 vdd.n31 13.1884
R18185 vdd.n1107 vdd.n1072 13.1884
R18186 vdd.n1154 vdd.n1119 13.1884
R18187 vdd.n1017 vdd.n982 13.1884
R18188 vdd.n1064 vdd.n1029 13.1884
R18189 vdd.n928 vdd.n893 13.1884
R18190 vdd.n975 vdd.n940 13.1884
R18191 vdd.n1391 vdd.n1256 12.9944
R18192 vdd.n1395 vdd.n1256 12.9944
R18193 vdd.n1691 vdd.n1543 12.9944
R18194 vdd.n1692 vdd.n1691 12.9944
R18195 vdd.n2988 vdd.n364 12.9944
R18196 vdd.n2989 vdd.n2988 12.9944
R18197 vdd.n2806 vdd.n536 12.9944
R18198 vdd.n2809 vdd.n2806 12.9944
R18199 vdd.n293 vdd.n255 12.8005
R18200 vdd.n288 vdd.n259 12.8005
R18201 vdd.n246 vdd.n208 12.8005
R18202 vdd.n241 vdd.n212 12.8005
R18203 vdd.n203 vdd.n165 12.8005
R18204 vdd.n198 vdd.n169 12.8005
R18205 vdd.n156 vdd.n118 12.8005
R18206 vdd.n151 vdd.n122 12.8005
R18207 vdd.n114 vdd.n76 12.8005
R18208 vdd.n109 vdd.n80 12.8005
R18209 vdd.n67 vdd.n29 12.8005
R18210 vdd.n62 vdd.n33 12.8005
R18211 vdd.n1108 vdd.n1070 12.8005
R18212 vdd.n1103 vdd.n1074 12.8005
R18213 vdd.n1155 vdd.n1117 12.8005
R18214 vdd.n1150 vdd.n1121 12.8005
R18215 vdd.n1018 vdd.n980 12.8005
R18216 vdd.n1013 vdd.n984 12.8005
R18217 vdd.n1065 vdd.n1027 12.8005
R18218 vdd.n1060 vdd.n1031 12.8005
R18219 vdd.n929 vdd.n891 12.8005
R18220 vdd.n924 vdd.n895 12.8005
R18221 vdd.n976 vdd.n938 12.8005
R18222 vdd.n971 vdd.n942 12.8005
R18223 vdd.n287 vdd.n260 12.0247
R18224 vdd.n240 vdd.n213 12.0247
R18225 vdd.n197 vdd.n170 12.0247
R18226 vdd.n150 vdd.n123 12.0247
R18227 vdd.n108 vdd.n81 12.0247
R18228 vdd.n61 vdd.n34 12.0247
R18229 vdd.n1102 vdd.n1075 12.0247
R18230 vdd.n1149 vdd.n1122 12.0247
R18231 vdd.n1012 vdd.n985 12.0247
R18232 vdd.n1059 vdd.n1032 12.0247
R18233 vdd.n923 vdd.n896 12.0247
R18234 vdd.n970 vdd.n943 12.0247
R18235 vdd.n1430 vdd.n1186 11.337
R18236 vdd.n1439 vdd.n1186 11.337
R18237 vdd.n1439 vdd.n1438 11.337
R18238 vdd.n1447 vdd.n1180 11.337
R18239 vdd.n1456 vdd.n1455 11.337
R18240 vdd.n1473 vdd.n1164 11.337
R18241 vdd.n1481 vdd.n887 11.337
R18242 vdd.n1490 vdd.n1489 11.337
R18243 vdd.n1498 vdd.n870 11.337
R18244 vdd.n1509 vdd.n870 11.337
R18245 vdd.n1509 vdd.n1508 11.337
R18246 vdd.n2849 vdd.n473 11.337
R18247 vdd.n2858 vdd.n473 11.337
R18248 vdd.n2858 vdd.n2857 11.337
R18249 vdd.n2866 vdd.n467 11.337
R18250 vdd.n2882 vdd.n456 11.337
R18251 vdd.n3043 vdd.n304 11.337
R18252 vdd.n3041 vdd.n308 11.337
R18253 vdd.n3035 vdd.n3034 11.337
R18254 vdd.n3033 vdd.n318 11.337
R18255 vdd.n3027 vdd.n318 11.337
R18256 vdd.n3027 vdd.n3026 11.337
R18257 vdd.n284 vdd.n283 11.249
R18258 vdd.n237 vdd.n236 11.249
R18259 vdd.n194 vdd.n193 11.249
R18260 vdd.n147 vdd.n146 11.249
R18261 vdd.n105 vdd.n104 11.249
R18262 vdd.n58 vdd.n57 11.249
R18263 vdd.n1099 vdd.n1098 11.249
R18264 vdd.n1146 vdd.n1145 11.249
R18265 vdd.n1009 vdd.n1008 11.249
R18266 vdd.n1056 vdd.n1055 11.249
R18267 vdd.n920 vdd.n919 11.249
R18268 vdd.n967 vdd.n966 11.249
R18269 vdd.n2146 vdd.t194 11.1103
R18270 vdd.n2478 vdd.t5 11.1103
R18271 vdd.n1228 vdd.t26 10.7702
R18272 vdd.t37 vdd.n3025 10.7702
R18273 vdd.n269 vdd.n268 10.7238
R18274 vdd.n222 vdd.n221 10.7238
R18275 vdd.n179 vdd.n178 10.7238
R18276 vdd.n132 vdd.n131 10.7238
R18277 vdd.n90 vdd.n89 10.7238
R18278 vdd.n43 vdd.n42 10.7238
R18279 vdd.n1084 vdd.n1083 10.7238
R18280 vdd.n1131 vdd.n1130 10.7238
R18281 vdd.n994 vdd.n993 10.7238
R18282 vdd.n1041 vdd.n1040 10.7238
R18283 vdd.n905 vdd.n904 10.7238
R18284 vdd.n952 vdd.n951 10.7238
R18285 vdd.n1992 vdd.n1991 10.6151
R18286 vdd.n1993 vdd.n1992 10.6151
R18287 vdd.n1993 vdd.n825 10.6151
R18288 vdd.n2003 vdd.n825 10.6151
R18289 vdd.n2004 vdd.n2003 10.6151
R18290 vdd.n2005 vdd.n2004 10.6151
R18291 vdd.n2005 vdd.n812 10.6151
R18292 vdd.n2016 vdd.n812 10.6151
R18293 vdd.n2017 vdd.n2016 10.6151
R18294 vdd.n2018 vdd.n2017 10.6151
R18295 vdd.n2018 vdd.n800 10.6151
R18296 vdd.n2028 vdd.n800 10.6151
R18297 vdd.n2029 vdd.n2028 10.6151
R18298 vdd.n2030 vdd.n2029 10.6151
R18299 vdd.n2030 vdd.n788 10.6151
R18300 vdd.n2040 vdd.n788 10.6151
R18301 vdd.n2041 vdd.n2040 10.6151
R18302 vdd.n2042 vdd.n2041 10.6151
R18303 vdd.n2042 vdd.n777 10.6151
R18304 vdd.n2052 vdd.n777 10.6151
R18305 vdd.n2053 vdd.n2052 10.6151
R18306 vdd.n2054 vdd.n2053 10.6151
R18307 vdd.n2054 vdd.n764 10.6151
R18308 vdd.n2066 vdd.n764 10.6151
R18309 vdd.n2067 vdd.n2066 10.6151
R18310 vdd.n2069 vdd.n2067 10.6151
R18311 vdd.n2069 vdd.n2068 10.6151
R18312 vdd.n2068 vdd.n746 10.6151
R18313 vdd.n2216 vdd.n2215 10.6151
R18314 vdd.n2215 vdd.n2214 10.6151
R18315 vdd.n2214 vdd.n2211 10.6151
R18316 vdd.n2211 vdd.n2210 10.6151
R18317 vdd.n2210 vdd.n2207 10.6151
R18318 vdd.n2207 vdd.n2206 10.6151
R18319 vdd.n2206 vdd.n2203 10.6151
R18320 vdd.n2203 vdd.n2202 10.6151
R18321 vdd.n2202 vdd.n2199 10.6151
R18322 vdd.n2199 vdd.n2198 10.6151
R18323 vdd.n2198 vdd.n2195 10.6151
R18324 vdd.n2195 vdd.n2194 10.6151
R18325 vdd.n2194 vdd.n2191 10.6151
R18326 vdd.n2191 vdd.n2190 10.6151
R18327 vdd.n2190 vdd.n2187 10.6151
R18328 vdd.n2187 vdd.n2186 10.6151
R18329 vdd.n2186 vdd.n2183 10.6151
R18330 vdd.n2183 vdd.n2182 10.6151
R18331 vdd.n2182 vdd.n2179 10.6151
R18332 vdd.n2179 vdd.n2178 10.6151
R18333 vdd.n2178 vdd.n2175 10.6151
R18334 vdd.n2175 vdd.n2174 10.6151
R18335 vdd.n2174 vdd.n2171 10.6151
R18336 vdd.n2171 vdd.n2170 10.6151
R18337 vdd.n2170 vdd.n2167 10.6151
R18338 vdd.n2167 vdd.n2166 10.6151
R18339 vdd.n2166 vdd.n2163 10.6151
R18340 vdd.n2163 vdd.n2162 10.6151
R18341 vdd.n2162 vdd.n2159 10.6151
R18342 vdd.n2159 vdd.n2158 10.6151
R18343 vdd.n2158 vdd.n2155 10.6151
R18344 vdd.n2153 vdd.n2150 10.6151
R18345 vdd.n2150 vdd.n2149 10.6151
R18346 vdd.n1892 vdd.n1891 10.6151
R18347 vdd.n1891 vdd.n1889 10.6151
R18348 vdd.n1889 vdd.n1888 10.6151
R18349 vdd.n1888 vdd.n1886 10.6151
R18350 vdd.n1886 vdd.n1885 10.6151
R18351 vdd.n1885 vdd.n1883 10.6151
R18352 vdd.n1883 vdd.n1882 10.6151
R18353 vdd.n1882 vdd.n1880 10.6151
R18354 vdd.n1880 vdd.n1879 10.6151
R18355 vdd.n1879 vdd.n1877 10.6151
R18356 vdd.n1877 vdd.n1876 10.6151
R18357 vdd.n1876 vdd.n1874 10.6151
R18358 vdd.n1874 vdd.n1873 10.6151
R18359 vdd.n1873 vdd.n1788 10.6151
R18360 vdd.n1788 vdd.n1787 10.6151
R18361 vdd.n1787 vdd.n1785 10.6151
R18362 vdd.n1785 vdd.n1784 10.6151
R18363 vdd.n1784 vdd.n1782 10.6151
R18364 vdd.n1782 vdd.n1781 10.6151
R18365 vdd.n1781 vdd.n1779 10.6151
R18366 vdd.n1779 vdd.n1778 10.6151
R18367 vdd.n1778 vdd.n1776 10.6151
R18368 vdd.n1776 vdd.n1775 10.6151
R18369 vdd.n1775 vdd.n1773 10.6151
R18370 vdd.n1773 vdd.n1772 10.6151
R18371 vdd.n1772 vdd.n1769 10.6151
R18372 vdd.n1769 vdd.n1768 10.6151
R18373 vdd.n1768 vdd.n749 10.6151
R18374 vdd.n1726 vdd.n837 10.6151
R18375 vdd.n1727 vdd.n1726 10.6151
R18376 vdd.n1728 vdd.n1727 10.6151
R18377 vdd.n1728 vdd.n1722 10.6151
R18378 vdd.n1734 vdd.n1722 10.6151
R18379 vdd.n1735 vdd.n1734 10.6151
R18380 vdd.n1736 vdd.n1735 10.6151
R18381 vdd.n1736 vdd.n1720 10.6151
R18382 vdd.n1742 vdd.n1720 10.6151
R18383 vdd.n1743 vdd.n1742 10.6151
R18384 vdd.n1744 vdd.n1743 10.6151
R18385 vdd.n1744 vdd.n1718 10.6151
R18386 vdd.n1750 vdd.n1718 10.6151
R18387 vdd.n1751 vdd.n1750 10.6151
R18388 vdd.n1752 vdd.n1751 10.6151
R18389 vdd.n1752 vdd.n1716 10.6151
R18390 vdd.n1928 vdd.n1716 10.6151
R18391 vdd.n1928 vdd.n1927 10.6151
R18392 vdd.n1927 vdd.n1757 10.6151
R18393 vdd.n1921 vdd.n1757 10.6151
R18394 vdd.n1921 vdd.n1920 10.6151
R18395 vdd.n1920 vdd.n1919 10.6151
R18396 vdd.n1919 vdd.n1759 10.6151
R18397 vdd.n1913 vdd.n1759 10.6151
R18398 vdd.n1913 vdd.n1912 10.6151
R18399 vdd.n1912 vdd.n1911 10.6151
R18400 vdd.n1911 vdd.n1761 10.6151
R18401 vdd.n1905 vdd.n1761 10.6151
R18402 vdd.n1905 vdd.n1904 10.6151
R18403 vdd.n1904 vdd.n1903 10.6151
R18404 vdd.n1903 vdd.n1763 10.6151
R18405 vdd.n1897 vdd.n1896 10.6151
R18406 vdd.n1896 vdd.n1895 10.6151
R18407 vdd.n2401 vdd.n2400 10.6151
R18408 vdd.n2400 vdd.n2398 10.6151
R18409 vdd.n2398 vdd.n2397 10.6151
R18410 vdd.n2397 vdd.n2255 10.6151
R18411 vdd.n2344 vdd.n2255 10.6151
R18412 vdd.n2345 vdd.n2344 10.6151
R18413 vdd.n2347 vdd.n2345 10.6151
R18414 vdd.n2348 vdd.n2347 10.6151
R18415 vdd.n2350 vdd.n2348 10.6151
R18416 vdd.n2351 vdd.n2350 10.6151
R18417 vdd.n2353 vdd.n2351 10.6151
R18418 vdd.n2354 vdd.n2353 10.6151
R18419 vdd.n2356 vdd.n2354 10.6151
R18420 vdd.n2357 vdd.n2356 10.6151
R18421 vdd.n2372 vdd.n2357 10.6151
R18422 vdd.n2372 vdd.n2371 10.6151
R18423 vdd.n2371 vdd.n2370 10.6151
R18424 vdd.n2370 vdd.n2368 10.6151
R18425 vdd.n2368 vdd.n2367 10.6151
R18426 vdd.n2367 vdd.n2365 10.6151
R18427 vdd.n2365 vdd.n2364 10.6151
R18428 vdd.n2364 vdd.n2362 10.6151
R18429 vdd.n2362 vdd.n2361 10.6151
R18430 vdd.n2361 vdd.n2359 10.6151
R18431 vdd.n2359 vdd.n2358 10.6151
R18432 vdd.n2358 vdd.n626 10.6151
R18433 vdd.n2606 vdd.n626 10.6151
R18434 vdd.n2607 vdd.n2606 10.6151
R18435 vdd.n2468 vdd.n702 10.6151
R18436 vdd.n2468 vdd.n2467 10.6151
R18437 vdd.n2467 vdd.n2466 10.6151
R18438 vdd.n2466 vdd.n2464 10.6151
R18439 vdd.n2464 vdd.n2461 10.6151
R18440 vdd.n2461 vdd.n2460 10.6151
R18441 vdd.n2460 vdd.n2457 10.6151
R18442 vdd.n2457 vdd.n2456 10.6151
R18443 vdd.n2456 vdd.n2453 10.6151
R18444 vdd.n2453 vdd.n2452 10.6151
R18445 vdd.n2452 vdd.n2449 10.6151
R18446 vdd.n2449 vdd.n2448 10.6151
R18447 vdd.n2448 vdd.n2445 10.6151
R18448 vdd.n2445 vdd.n2444 10.6151
R18449 vdd.n2444 vdd.n2441 10.6151
R18450 vdd.n2441 vdd.n2440 10.6151
R18451 vdd.n2440 vdd.n2437 10.6151
R18452 vdd.n2437 vdd.n2436 10.6151
R18453 vdd.n2436 vdd.n2433 10.6151
R18454 vdd.n2433 vdd.n2432 10.6151
R18455 vdd.n2432 vdd.n2429 10.6151
R18456 vdd.n2429 vdd.n2428 10.6151
R18457 vdd.n2428 vdd.n2425 10.6151
R18458 vdd.n2425 vdd.n2424 10.6151
R18459 vdd.n2424 vdd.n2421 10.6151
R18460 vdd.n2421 vdd.n2420 10.6151
R18461 vdd.n2420 vdd.n2417 10.6151
R18462 vdd.n2417 vdd.n2416 10.6151
R18463 vdd.n2416 vdd.n2413 10.6151
R18464 vdd.n2413 vdd.n2412 10.6151
R18465 vdd.n2412 vdd.n2409 10.6151
R18466 vdd.n2407 vdd.n2404 10.6151
R18467 vdd.n2404 vdd.n2403 10.6151
R18468 vdd.n2481 vdd.n2480 10.6151
R18469 vdd.n2482 vdd.n2481 10.6151
R18470 vdd.n2482 vdd.n692 10.6151
R18471 vdd.n2492 vdd.n692 10.6151
R18472 vdd.n2493 vdd.n2492 10.6151
R18473 vdd.n2494 vdd.n2493 10.6151
R18474 vdd.n2494 vdd.n679 10.6151
R18475 vdd.n2504 vdd.n679 10.6151
R18476 vdd.n2505 vdd.n2504 10.6151
R18477 vdd.n2506 vdd.n2505 10.6151
R18478 vdd.n2506 vdd.n668 10.6151
R18479 vdd.n2516 vdd.n668 10.6151
R18480 vdd.n2517 vdd.n2516 10.6151
R18481 vdd.n2518 vdd.n2517 10.6151
R18482 vdd.n2518 vdd.n656 10.6151
R18483 vdd.n2528 vdd.n656 10.6151
R18484 vdd.n2529 vdd.n2528 10.6151
R18485 vdd.n2530 vdd.n2529 10.6151
R18486 vdd.n2530 vdd.n645 10.6151
R18487 vdd.n2542 vdd.n645 10.6151
R18488 vdd.n2543 vdd.n2542 10.6151
R18489 vdd.n2544 vdd.n2543 10.6151
R18490 vdd.n2544 vdd.n631 10.6151
R18491 vdd.n2599 vdd.n631 10.6151
R18492 vdd.n2600 vdd.n2599 10.6151
R18493 vdd.n2601 vdd.n2600 10.6151
R18494 vdd.n2601 vdd.n600 10.6151
R18495 vdd.n2671 vdd.n600 10.6151
R18496 vdd.n2670 vdd.n2669 10.6151
R18497 vdd.n2669 vdd.n601 10.6151
R18498 vdd.n602 vdd.n601 10.6151
R18499 vdd.n2662 vdd.n602 10.6151
R18500 vdd.n2662 vdd.n2661 10.6151
R18501 vdd.n2661 vdd.n2660 10.6151
R18502 vdd.n2660 vdd.n604 10.6151
R18503 vdd.n2655 vdd.n604 10.6151
R18504 vdd.n2655 vdd.n2654 10.6151
R18505 vdd.n2654 vdd.n2653 10.6151
R18506 vdd.n2653 vdd.n607 10.6151
R18507 vdd.n2648 vdd.n607 10.6151
R18508 vdd.n2648 vdd.n2647 10.6151
R18509 vdd.n2647 vdd.n2646 10.6151
R18510 vdd.n2646 vdd.n610 10.6151
R18511 vdd.n2641 vdd.n610 10.6151
R18512 vdd.n2641 vdd.n520 10.6151
R18513 vdd.n2637 vdd.n520 10.6151
R18514 vdd.n2637 vdd.n2636 10.6151
R18515 vdd.n2636 vdd.n2635 10.6151
R18516 vdd.n2635 vdd.n613 10.6151
R18517 vdd.n2630 vdd.n613 10.6151
R18518 vdd.n2630 vdd.n2629 10.6151
R18519 vdd.n2629 vdd.n2628 10.6151
R18520 vdd.n2628 vdd.n616 10.6151
R18521 vdd.n2623 vdd.n616 10.6151
R18522 vdd.n2623 vdd.n2622 10.6151
R18523 vdd.n2622 vdd.n2621 10.6151
R18524 vdd.n2621 vdd.n619 10.6151
R18525 vdd.n2616 vdd.n619 10.6151
R18526 vdd.n2616 vdd.n2615 10.6151
R18527 vdd.n2613 vdd.n624 10.6151
R18528 vdd.n2608 vdd.n624 10.6151
R18529 vdd.n2589 vdd.n2550 10.6151
R18530 vdd.n2584 vdd.n2550 10.6151
R18531 vdd.n2584 vdd.n2583 10.6151
R18532 vdd.n2583 vdd.n2582 10.6151
R18533 vdd.n2582 vdd.n2552 10.6151
R18534 vdd.n2577 vdd.n2552 10.6151
R18535 vdd.n2577 vdd.n2576 10.6151
R18536 vdd.n2576 vdd.n2575 10.6151
R18537 vdd.n2575 vdd.n2555 10.6151
R18538 vdd.n2570 vdd.n2555 10.6151
R18539 vdd.n2570 vdd.n2569 10.6151
R18540 vdd.n2569 vdd.n2568 10.6151
R18541 vdd.n2568 vdd.n2558 10.6151
R18542 vdd.n2563 vdd.n2558 10.6151
R18543 vdd.n2563 vdd.n2562 10.6151
R18544 vdd.n2562 vdd.n575 10.6151
R18545 vdd.n2706 vdd.n575 10.6151
R18546 vdd.n2706 vdd.n576 10.6151
R18547 vdd.n578 vdd.n576 10.6151
R18548 vdd.n2699 vdd.n578 10.6151
R18549 vdd.n2699 vdd.n2698 10.6151
R18550 vdd.n2698 vdd.n2697 10.6151
R18551 vdd.n2697 vdd.n580 10.6151
R18552 vdd.n2692 vdd.n580 10.6151
R18553 vdd.n2692 vdd.n2691 10.6151
R18554 vdd.n2691 vdd.n2690 10.6151
R18555 vdd.n2690 vdd.n583 10.6151
R18556 vdd.n2685 vdd.n583 10.6151
R18557 vdd.n2685 vdd.n2684 10.6151
R18558 vdd.n2684 vdd.n2683 10.6151
R18559 vdd.n2683 vdd.n586 10.6151
R18560 vdd.n2678 vdd.n2677 10.6151
R18561 vdd.n2677 vdd.n2676 10.6151
R18562 vdd.n2324 vdd.n2322 10.6151
R18563 vdd.n2325 vdd.n2324 10.6151
R18564 vdd.n2393 vdd.n2325 10.6151
R18565 vdd.n2393 vdd.n2392 10.6151
R18566 vdd.n2392 vdd.n2391 10.6151
R18567 vdd.n2391 vdd.n2389 10.6151
R18568 vdd.n2389 vdd.n2388 10.6151
R18569 vdd.n2388 vdd.n2386 10.6151
R18570 vdd.n2386 vdd.n2385 10.6151
R18571 vdd.n2385 vdd.n2383 10.6151
R18572 vdd.n2383 vdd.n2382 10.6151
R18573 vdd.n2382 vdd.n2380 10.6151
R18574 vdd.n2380 vdd.n2379 10.6151
R18575 vdd.n2379 vdd.n2377 10.6151
R18576 vdd.n2377 vdd.n2376 10.6151
R18577 vdd.n2376 vdd.n2342 10.6151
R18578 vdd.n2342 vdd.n2341 10.6151
R18579 vdd.n2341 vdd.n2339 10.6151
R18580 vdd.n2339 vdd.n2338 10.6151
R18581 vdd.n2338 vdd.n2336 10.6151
R18582 vdd.n2336 vdd.n2335 10.6151
R18583 vdd.n2335 vdd.n2333 10.6151
R18584 vdd.n2333 vdd.n2332 10.6151
R18585 vdd.n2332 vdd.n2330 10.6151
R18586 vdd.n2330 vdd.n2329 10.6151
R18587 vdd.n2329 vdd.n2327 10.6151
R18588 vdd.n2327 vdd.n2326 10.6151
R18589 vdd.n2326 vdd.n592 10.6151
R18590 vdd.n2475 vdd.n2474 10.6151
R18591 vdd.n2474 vdd.n707 10.6151
R18592 vdd.n2259 vdd.n707 10.6151
R18593 vdd.n2262 vdd.n2259 10.6151
R18594 vdd.n2263 vdd.n2262 10.6151
R18595 vdd.n2266 vdd.n2263 10.6151
R18596 vdd.n2267 vdd.n2266 10.6151
R18597 vdd.n2270 vdd.n2267 10.6151
R18598 vdd.n2271 vdd.n2270 10.6151
R18599 vdd.n2274 vdd.n2271 10.6151
R18600 vdd.n2275 vdd.n2274 10.6151
R18601 vdd.n2278 vdd.n2275 10.6151
R18602 vdd.n2279 vdd.n2278 10.6151
R18603 vdd.n2282 vdd.n2279 10.6151
R18604 vdd.n2283 vdd.n2282 10.6151
R18605 vdd.n2286 vdd.n2283 10.6151
R18606 vdd.n2287 vdd.n2286 10.6151
R18607 vdd.n2290 vdd.n2287 10.6151
R18608 vdd.n2291 vdd.n2290 10.6151
R18609 vdd.n2294 vdd.n2291 10.6151
R18610 vdd.n2295 vdd.n2294 10.6151
R18611 vdd.n2298 vdd.n2295 10.6151
R18612 vdd.n2299 vdd.n2298 10.6151
R18613 vdd.n2302 vdd.n2299 10.6151
R18614 vdd.n2303 vdd.n2302 10.6151
R18615 vdd.n2306 vdd.n2303 10.6151
R18616 vdd.n2307 vdd.n2306 10.6151
R18617 vdd.n2310 vdd.n2307 10.6151
R18618 vdd.n2311 vdd.n2310 10.6151
R18619 vdd.n2314 vdd.n2311 10.6151
R18620 vdd.n2315 vdd.n2314 10.6151
R18621 vdd.n2320 vdd.n2318 10.6151
R18622 vdd.n2321 vdd.n2320 10.6151
R18623 vdd.n2476 vdd.n697 10.6151
R18624 vdd.n2486 vdd.n697 10.6151
R18625 vdd.n2487 vdd.n2486 10.6151
R18626 vdd.n2488 vdd.n2487 10.6151
R18627 vdd.n2488 vdd.n685 10.6151
R18628 vdd.n2498 vdd.n685 10.6151
R18629 vdd.n2499 vdd.n2498 10.6151
R18630 vdd.n2500 vdd.n2499 10.6151
R18631 vdd.n2500 vdd.n674 10.6151
R18632 vdd.n2510 vdd.n674 10.6151
R18633 vdd.n2511 vdd.n2510 10.6151
R18634 vdd.n2512 vdd.n2511 10.6151
R18635 vdd.n2512 vdd.n662 10.6151
R18636 vdd.n2522 vdd.n662 10.6151
R18637 vdd.n2523 vdd.n2522 10.6151
R18638 vdd.n2524 vdd.n2523 10.6151
R18639 vdd.n2524 vdd.n651 10.6151
R18640 vdd.n2534 vdd.n651 10.6151
R18641 vdd.n2535 vdd.n2534 10.6151
R18642 vdd.n2538 vdd.n2535 10.6151
R18643 vdd.n2548 vdd.n639 10.6151
R18644 vdd.n2549 vdd.n2548 10.6151
R18645 vdd.n2595 vdd.n2549 10.6151
R18646 vdd.n2595 vdd.n2594 10.6151
R18647 vdd.n2594 vdd.n2593 10.6151
R18648 vdd.n2593 vdd.n2592 10.6151
R18649 vdd.n2592 vdd.n2590 10.6151
R18650 vdd.n1987 vdd.n831 10.6151
R18651 vdd.n1997 vdd.n831 10.6151
R18652 vdd.n1998 vdd.n1997 10.6151
R18653 vdd.n1999 vdd.n1998 10.6151
R18654 vdd.n1999 vdd.n818 10.6151
R18655 vdd.n2009 vdd.n818 10.6151
R18656 vdd.n2010 vdd.n2009 10.6151
R18657 vdd.n2012 vdd.n806 10.6151
R18658 vdd.n2022 vdd.n806 10.6151
R18659 vdd.n2023 vdd.n2022 10.6151
R18660 vdd.n2024 vdd.n2023 10.6151
R18661 vdd.n2024 vdd.n794 10.6151
R18662 vdd.n2034 vdd.n794 10.6151
R18663 vdd.n2035 vdd.n2034 10.6151
R18664 vdd.n2036 vdd.n2035 10.6151
R18665 vdd.n2036 vdd.n783 10.6151
R18666 vdd.n2046 vdd.n783 10.6151
R18667 vdd.n2047 vdd.n2046 10.6151
R18668 vdd.n2048 vdd.n2047 10.6151
R18669 vdd.n2048 vdd.n771 10.6151
R18670 vdd.n2058 vdd.n771 10.6151
R18671 vdd.n2059 vdd.n2058 10.6151
R18672 vdd.n2062 vdd.n2059 10.6151
R18673 vdd.n2062 vdd.n2061 10.6151
R18674 vdd.n2061 vdd.n2060 10.6151
R18675 vdd.n2060 vdd.n754 10.6151
R18676 vdd.n2144 vdd.n754 10.6151
R18677 vdd.n2143 vdd.n2142 10.6151
R18678 vdd.n2142 vdd.n2139 10.6151
R18679 vdd.n2139 vdd.n2138 10.6151
R18680 vdd.n2138 vdd.n2135 10.6151
R18681 vdd.n2135 vdd.n2134 10.6151
R18682 vdd.n2134 vdd.n2131 10.6151
R18683 vdd.n2131 vdd.n2130 10.6151
R18684 vdd.n2130 vdd.n2127 10.6151
R18685 vdd.n2127 vdd.n2126 10.6151
R18686 vdd.n2126 vdd.n2123 10.6151
R18687 vdd.n2123 vdd.n2122 10.6151
R18688 vdd.n2122 vdd.n2119 10.6151
R18689 vdd.n2119 vdd.n2118 10.6151
R18690 vdd.n2118 vdd.n2115 10.6151
R18691 vdd.n2115 vdd.n2114 10.6151
R18692 vdd.n2114 vdd.n2111 10.6151
R18693 vdd.n2111 vdd.n2110 10.6151
R18694 vdd.n2110 vdd.n2107 10.6151
R18695 vdd.n2107 vdd.n2106 10.6151
R18696 vdd.n2106 vdd.n2103 10.6151
R18697 vdd.n2103 vdd.n2102 10.6151
R18698 vdd.n2102 vdd.n2099 10.6151
R18699 vdd.n2099 vdd.n2098 10.6151
R18700 vdd.n2098 vdd.n2095 10.6151
R18701 vdd.n2095 vdd.n2094 10.6151
R18702 vdd.n2094 vdd.n2091 10.6151
R18703 vdd.n2091 vdd.n2090 10.6151
R18704 vdd.n2090 vdd.n2087 10.6151
R18705 vdd.n2087 vdd.n2086 10.6151
R18706 vdd.n2086 vdd.n2083 10.6151
R18707 vdd.n2083 vdd.n2082 10.6151
R18708 vdd.n2079 vdd.n2078 10.6151
R18709 vdd.n2078 vdd.n2076 10.6151
R18710 vdd.n1835 vdd.n1833 10.6151
R18711 vdd.n1836 vdd.n1835 10.6151
R18712 vdd.n1838 vdd.n1836 10.6151
R18713 vdd.n1839 vdd.n1838 10.6151
R18714 vdd.n1841 vdd.n1839 10.6151
R18715 vdd.n1842 vdd.n1841 10.6151
R18716 vdd.n1844 vdd.n1842 10.6151
R18717 vdd.n1845 vdd.n1844 10.6151
R18718 vdd.n1847 vdd.n1845 10.6151
R18719 vdd.n1848 vdd.n1847 10.6151
R18720 vdd.n1850 vdd.n1848 10.6151
R18721 vdd.n1851 vdd.n1850 10.6151
R18722 vdd.n1869 vdd.n1851 10.6151
R18723 vdd.n1869 vdd.n1868 10.6151
R18724 vdd.n1868 vdd.n1867 10.6151
R18725 vdd.n1867 vdd.n1865 10.6151
R18726 vdd.n1865 vdd.n1864 10.6151
R18727 vdd.n1864 vdd.n1862 10.6151
R18728 vdd.n1862 vdd.n1861 10.6151
R18729 vdd.n1861 vdd.n1859 10.6151
R18730 vdd.n1859 vdd.n1858 10.6151
R18731 vdd.n1858 vdd.n1856 10.6151
R18732 vdd.n1856 vdd.n1855 10.6151
R18733 vdd.n1855 vdd.n1853 10.6151
R18734 vdd.n1853 vdd.n1852 10.6151
R18735 vdd.n1852 vdd.n758 10.6151
R18736 vdd.n2074 vdd.n758 10.6151
R18737 vdd.n2075 vdd.n2074 10.6151
R18738 vdd.n1986 vdd.n1985 10.6151
R18739 vdd.n1985 vdd.n843 10.6151
R18740 vdd.n1979 vdd.n843 10.6151
R18741 vdd.n1979 vdd.n1978 10.6151
R18742 vdd.n1978 vdd.n1977 10.6151
R18743 vdd.n1977 vdd.n845 10.6151
R18744 vdd.n1971 vdd.n845 10.6151
R18745 vdd.n1971 vdd.n1970 10.6151
R18746 vdd.n1970 vdd.n1969 10.6151
R18747 vdd.n1969 vdd.n847 10.6151
R18748 vdd.n1963 vdd.n847 10.6151
R18749 vdd.n1963 vdd.n1962 10.6151
R18750 vdd.n1962 vdd.n1961 10.6151
R18751 vdd.n1961 vdd.n849 10.6151
R18752 vdd.n1955 vdd.n849 10.6151
R18753 vdd.n1955 vdd.n1954 10.6151
R18754 vdd.n1954 vdd.n1953 10.6151
R18755 vdd.n1953 vdd.n853 10.6151
R18756 vdd.n1801 vdd.n853 10.6151
R18757 vdd.n1802 vdd.n1801 10.6151
R18758 vdd.n1802 vdd.n1797 10.6151
R18759 vdd.n1808 vdd.n1797 10.6151
R18760 vdd.n1809 vdd.n1808 10.6151
R18761 vdd.n1810 vdd.n1809 10.6151
R18762 vdd.n1810 vdd.n1795 10.6151
R18763 vdd.n1816 vdd.n1795 10.6151
R18764 vdd.n1817 vdd.n1816 10.6151
R18765 vdd.n1818 vdd.n1817 10.6151
R18766 vdd.n1818 vdd.n1793 10.6151
R18767 vdd.n1824 vdd.n1793 10.6151
R18768 vdd.n1825 vdd.n1824 10.6151
R18769 vdd.n1827 vdd.n1789 10.6151
R18770 vdd.n1832 vdd.n1789 10.6151
R18771 vdd.n280 vdd.n262 10.4732
R18772 vdd.n233 vdd.n215 10.4732
R18773 vdd.n190 vdd.n172 10.4732
R18774 vdd.n143 vdd.n125 10.4732
R18775 vdd.n101 vdd.n83 10.4732
R18776 vdd.n54 vdd.n36 10.4732
R18777 vdd.n1095 vdd.n1077 10.4732
R18778 vdd.n1142 vdd.n1124 10.4732
R18779 vdd.n1005 vdd.n987 10.4732
R18780 vdd.n1052 vdd.n1034 10.4732
R18781 vdd.n916 vdd.n898 10.4732
R18782 vdd.n963 vdd.n945 10.4732
R18783 vdd.t120 vdd.n888 10.3167
R18784 vdd.n2874 vdd.t140 10.3167
R18785 vdd.n1465 vdd.t116 10.09
R18786 vdd.n3042 vdd.t153 10.09
R18787 vdd.n279 vdd.n264 9.69747
R18788 vdd.n232 vdd.n217 9.69747
R18789 vdd.n189 vdd.n174 9.69747
R18790 vdd.n142 vdd.n127 9.69747
R18791 vdd.n100 vdd.n85 9.69747
R18792 vdd.n53 vdd.n38 9.69747
R18793 vdd.n1094 vdd.n1079 9.69747
R18794 vdd.n1141 vdd.n1126 9.69747
R18795 vdd.n1004 vdd.n989 9.69747
R18796 vdd.n1051 vdd.n1036 9.69747
R18797 vdd.n915 vdd.n900 9.69747
R18798 vdd.n962 vdd.n947 9.69747
R18799 vdd.n1929 vdd.n1928 9.67831
R18800 vdd.n2836 vdd.n520 9.67831
R18801 vdd.n2707 vdd.n2706 9.67831
R18802 vdd.n1953 vdd.n1952 9.67831
R18803 vdd.n295 vdd.n294 9.45567
R18804 vdd.n248 vdd.n247 9.45567
R18805 vdd.n205 vdd.n204 9.45567
R18806 vdd.n158 vdd.n157 9.45567
R18807 vdd.n116 vdd.n115 9.45567
R18808 vdd.n69 vdd.n68 9.45567
R18809 vdd.n1110 vdd.n1109 9.45567
R18810 vdd.n1157 vdd.n1156 9.45567
R18811 vdd.n1020 vdd.n1019 9.45567
R18812 vdd.n1067 vdd.n1066 9.45567
R18813 vdd.n931 vdd.n930 9.45567
R18814 vdd.n978 vdd.n977 9.45567
R18815 vdd.n1689 vdd.n1543 9.3005
R18816 vdd.n1688 vdd.n1687 9.3005
R18817 vdd.n1549 vdd.n1548 9.3005
R18818 vdd.n1682 vdd.n1553 9.3005
R18819 vdd.n1681 vdd.n1554 9.3005
R18820 vdd.n1680 vdd.n1555 9.3005
R18821 vdd.n1559 vdd.n1556 9.3005
R18822 vdd.n1675 vdd.n1560 9.3005
R18823 vdd.n1674 vdd.n1561 9.3005
R18824 vdd.n1673 vdd.n1562 9.3005
R18825 vdd.n1566 vdd.n1563 9.3005
R18826 vdd.n1668 vdd.n1567 9.3005
R18827 vdd.n1667 vdd.n1568 9.3005
R18828 vdd.n1666 vdd.n1569 9.3005
R18829 vdd.n1573 vdd.n1570 9.3005
R18830 vdd.n1661 vdd.n1574 9.3005
R18831 vdd.n1660 vdd.n1575 9.3005
R18832 vdd.n1659 vdd.n1576 9.3005
R18833 vdd.n1580 vdd.n1577 9.3005
R18834 vdd.n1654 vdd.n1581 9.3005
R18835 vdd.n1653 vdd.n1582 9.3005
R18836 vdd.n1652 vdd.n1651 9.3005
R18837 vdd.n1650 vdd.n1583 9.3005
R18838 vdd.n1649 vdd.n1648 9.3005
R18839 vdd.n1589 vdd.n1588 9.3005
R18840 vdd.n1643 vdd.n1593 9.3005
R18841 vdd.n1642 vdd.n1594 9.3005
R18842 vdd.n1641 vdd.n1595 9.3005
R18843 vdd.n1599 vdd.n1596 9.3005
R18844 vdd.n1636 vdd.n1600 9.3005
R18845 vdd.n1635 vdd.n1601 9.3005
R18846 vdd.n1634 vdd.n1602 9.3005
R18847 vdd.n1606 vdd.n1603 9.3005
R18848 vdd.n1629 vdd.n1607 9.3005
R18849 vdd.n1628 vdd.n1608 9.3005
R18850 vdd.n1627 vdd.n1609 9.3005
R18851 vdd.n1611 vdd.n1610 9.3005
R18852 vdd.n1622 vdd.n854 9.3005
R18853 vdd.n1691 vdd.n1690 9.3005
R18854 vdd.n1715 vdd.n1714 9.3005
R18855 vdd.n1521 vdd.n1520 9.3005
R18856 vdd.n1526 vdd.n1524 9.3005
R18857 vdd.n1707 vdd.n1527 9.3005
R18858 vdd.n1706 vdd.n1528 9.3005
R18859 vdd.n1705 vdd.n1529 9.3005
R18860 vdd.n1533 vdd.n1530 9.3005
R18861 vdd.n1700 vdd.n1534 9.3005
R18862 vdd.n1699 vdd.n1535 9.3005
R18863 vdd.n1698 vdd.n1536 9.3005
R18864 vdd.n1540 vdd.n1537 9.3005
R18865 vdd.n1693 vdd.n1541 9.3005
R18866 vdd.n1692 vdd.n1542 9.3005
R18867 vdd.n1937 vdd.n1514 9.3005
R18868 vdd.n1939 vdd.n1938 9.3005
R18869 vdd.n1476 vdd.n1475 9.3005
R18870 vdd.n1477 vdd.n890 9.3005
R18871 vdd.n1479 vdd.n1478 9.3005
R18872 vdd.n880 vdd.n879 9.3005
R18873 vdd.n1493 vdd.n1492 9.3005
R18874 vdd.n1494 vdd.n878 9.3005
R18875 vdd.n1496 vdd.n1495 9.3005
R18876 vdd.n868 vdd.n867 9.3005
R18877 vdd.n1512 vdd.n1511 9.3005
R18878 vdd.n1513 vdd.n866 9.3005
R18879 vdd.n1941 vdd.n1940 9.3005
R18880 vdd.n271 vdd.n270 9.3005
R18881 vdd.n266 vdd.n265 9.3005
R18882 vdd.n277 vdd.n276 9.3005
R18883 vdd.n279 vdd.n278 9.3005
R18884 vdd.n262 vdd.n261 9.3005
R18885 vdd.n285 vdd.n284 9.3005
R18886 vdd.n287 vdd.n286 9.3005
R18887 vdd.n259 vdd.n256 9.3005
R18888 vdd.n294 vdd.n293 9.3005
R18889 vdd.n224 vdd.n223 9.3005
R18890 vdd.n219 vdd.n218 9.3005
R18891 vdd.n230 vdd.n229 9.3005
R18892 vdd.n232 vdd.n231 9.3005
R18893 vdd.n215 vdd.n214 9.3005
R18894 vdd.n238 vdd.n237 9.3005
R18895 vdd.n240 vdd.n239 9.3005
R18896 vdd.n212 vdd.n209 9.3005
R18897 vdd.n247 vdd.n246 9.3005
R18898 vdd.n181 vdd.n180 9.3005
R18899 vdd.n176 vdd.n175 9.3005
R18900 vdd.n187 vdd.n186 9.3005
R18901 vdd.n189 vdd.n188 9.3005
R18902 vdd.n172 vdd.n171 9.3005
R18903 vdd.n195 vdd.n194 9.3005
R18904 vdd.n197 vdd.n196 9.3005
R18905 vdd.n169 vdd.n166 9.3005
R18906 vdd.n204 vdd.n203 9.3005
R18907 vdd.n134 vdd.n133 9.3005
R18908 vdd.n129 vdd.n128 9.3005
R18909 vdd.n140 vdd.n139 9.3005
R18910 vdd.n142 vdd.n141 9.3005
R18911 vdd.n125 vdd.n124 9.3005
R18912 vdd.n148 vdd.n147 9.3005
R18913 vdd.n150 vdd.n149 9.3005
R18914 vdd.n122 vdd.n119 9.3005
R18915 vdd.n157 vdd.n156 9.3005
R18916 vdd.n92 vdd.n91 9.3005
R18917 vdd.n87 vdd.n86 9.3005
R18918 vdd.n98 vdd.n97 9.3005
R18919 vdd.n100 vdd.n99 9.3005
R18920 vdd.n83 vdd.n82 9.3005
R18921 vdd.n106 vdd.n105 9.3005
R18922 vdd.n108 vdd.n107 9.3005
R18923 vdd.n80 vdd.n77 9.3005
R18924 vdd.n115 vdd.n114 9.3005
R18925 vdd.n45 vdd.n44 9.3005
R18926 vdd.n40 vdd.n39 9.3005
R18927 vdd.n51 vdd.n50 9.3005
R18928 vdd.n53 vdd.n52 9.3005
R18929 vdd.n36 vdd.n35 9.3005
R18930 vdd.n59 vdd.n58 9.3005
R18931 vdd.n61 vdd.n60 9.3005
R18932 vdd.n33 vdd.n30 9.3005
R18933 vdd.n68 vdd.n67 9.3005
R18934 vdd.n2758 vdd.n2757 9.3005
R18935 vdd.n2761 vdd.n555 9.3005
R18936 vdd.n2762 vdd.n554 9.3005
R18937 vdd.n2765 vdd.n553 9.3005
R18938 vdd.n2766 vdd.n552 9.3005
R18939 vdd.n2769 vdd.n551 9.3005
R18940 vdd.n2770 vdd.n550 9.3005
R18941 vdd.n2773 vdd.n549 9.3005
R18942 vdd.n2774 vdd.n548 9.3005
R18943 vdd.n2777 vdd.n547 9.3005
R18944 vdd.n2778 vdd.n546 9.3005
R18945 vdd.n2781 vdd.n545 9.3005
R18946 vdd.n2782 vdd.n544 9.3005
R18947 vdd.n2785 vdd.n543 9.3005
R18948 vdd.n2786 vdd.n542 9.3005
R18949 vdd.n2789 vdd.n541 9.3005
R18950 vdd.n2790 vdd.n540 9.3005
R18951 vdd.n2793 vdd.n539 9.3005
R18952 vdd.n2794 vdd.n538 9.3005
R18953 vdd.n2797 vdd.n537 9.3005
R18954 vdd.n2801 vdd.n2800 9.3005
R18955 vdd.n2802 vdd.n536 9.3005
R18956 vdd.n2806 vdd.n2803 9.3005
R18957 vdd.n2809 vdd.n535 9.3005
R18958 vdd.n2810 vdd.n534 9.3005
R18959 vdd.n2813 vdd.n533 9.3005
R18960 vdd.n2814 vdd.n532 9.3005
R18961 vdd.n2817 vdd.n531 9.3005
R18962 vdd.n2818 vdd.n530 9.3005
R18963 vdd.n2821 vdd.n529 9.3005
R18964 vdd.n2822 vdd.n528 9.3005
R18965 vdd.n2825 vdd.n527 9.3005
R18966 vdd.n2826 vdd.n526 9.3005
R18967 vdd.n2829 vdd.n525 9.3005
R18968 vdd.n2830 vdd.n524 9.3005
R18969 vdd.n2833 vdd.n519 9.3005
R18970 vdd.n482 vdd.n481 9.3005
R18971 vdd.n2844 vdd.n2843 9.3005
R18972 vdd.n2847 vdd.n2846 9.3005
R18973 vdd.n471 vdd.n470 9.3005
R18974 vdd.n2861 vdd.n2860 9.3005
R18975 vdd.n2862 vdd.n469 9.3005
R18976 vdd.n2864 vdd.n2863 9.3005
R18977 vdd.n460 vdd.n459 9.3005
R18978 vdd.n2877 vdd.n2876 9.3005
R18979 vdd.n2878 vdd.n458 9.3005
R18980 vdd.n2880 vdd.n2879 9.3005
R18981 vdd.n300 vdd.n298 9.3005
R18982 vdd.n2845 vdd.n480 9.3005
R18983 vdd.n3046 vdd.n3045 9.3005
R18984 vdd.n301 vdd.n299 9.3005
R18985 vdd.n3039 vdd.n310 9.3005
R18986 vdd.n3038 vdd.n311 9.3005
R18987 vdd.n3037 vdd.n312 9.3005
R18988 vdd.n320 vdd.n313 9.3005
R18989 vdd.n3031 vdd.n321 9.3005
R18990 vdd.n3030 vdd.n322 9.3005
R18991 vdd.n3029 vdd.n323 9.3005
R18992 vdd.n331 vdd.n324 9.3005
R18993 vdd.n3023 vdd.n3022 9.3005
R18994 vdd.n3019 vdd.n332 9.3005
R18995 vdd.n3018 vdd.n335 9.3005
R18996 vdd.n339 vdd.n336 9.3005
R18997 vdd.n340 vdd.n337 9.3005
R18998 vdd.n3011 vdd.n341 9.3005
R18999 vdd.n3010 vdd.n342 9.3005
R19000 vdd.n3009 vdd.n343 9.3005
R19001 vdd.n347 vdd.n344 9.3005
R19002 vdd.n3004 vdd.n348 9.3005
R19003 vdd.n3003 vdd.n349 9.3005
R19004 vdd.n3002 vdd.n350 9.3005
R19005 vdd.n354 vdd.n351 9.3005
R19006 vdd.n2997 vdd.n355 9.3005
R19007 vdd.n2996 vdd.n356 9.3005
R19008 vdd.n2995 vdd.n357 9.3005
R19009 vdd.n361 vdd.n358 9.3005
R19010 vdd.n2990 vdd.n362 9.3005
R19011 vdd.n2989 vdd.n363 9.3005
R19012 vdd.n2988 vdd.n2987 9.3005
R19013 vdd.n2986 vdd.n364 9.3005
R19014 vdd.n2985 vdd.n2984 9.3005
R19015 vdd.n370 vdd.n369 9.3005
R19016 vdd.n2979 vdd.n374 9.3005
R19017 vdd.n2978 vdd.n375 9.3005
R19018 vdd.n2977 vdd.n376 9.3005
R19019 vdd.n380 vdd.n377 9.3005
R19020 vdd.n2972 vdd.n381 9.3005
R19021 vdd.n2971 vdd.n382 9.3005
R19022 vdd.n2970 vdd.n383 9.3005
R19023 vdd.n387 vdd.n384 9.3005
R19024 vdd.n2965 vdd.n388 9.3005
R19025 vdd.n2964 vdd.n389 9.3005
R19026 vdd.n2963 vdd.n390 9.3005
R19027 vdd.n394 vdd.n391 9.3005
R19028 vdd.n2958 vdd.n395 9.3005
R19029 vdd.n2957 vdd.n396 9.3005
R19030 vdd.n2956 vdd.n397 9.3005
R19031 vdd.n401 vdd.n398 9.3005
R19032 vdd.n2951 vdd.n402 9.3005
R19033 vdd.n2950 vdd.n403 9.3005
R19034 vdd.n2949 vdd.n2948 9.3005
R19035 vdd.n2947 vdd.n404 9.3005
R19036 vdd.n2946 vdd.n2945 9.3005
R19037 vdd.n410 vdd.n409 9.3005
R19038 vdd.n2940 vdd.n414 9.3005
R19039 vdd.n2939 vdd.n415 9.3005
R19040 vdd.n2938 vdd.n416 9.3005
R19041 vdd.n420 vdd.n417 9.3005
R19042 vdd.n2933 vdd.n421 9.3005
R19043 vdd.n2932 vdd.n422 9.3005
R19044 vdd.n2931 vdd.n423 9.3005
R19045 vdd.n427 vdd.n424 9.3005
R19046 vdd.n2926 vdd.n428 9.3005
R19047 vdd.n2925 vdd.n429 9.3005
R19048 vdd.n2924 vdd.n430 9.3005
R19049 vdd.n434 vdd.n431 9.3005
R19050 vdd.n2919 vdd.n435 9.3005
R19051 vdd.n2918 vdd.n436 9.3005
R19052 vdd.n2917 vdd.n437 9.3005
R19053 vdd.n441 vdd.n438 9.3005
R19054 vdd.n2912 vdd.n442 9.3005
R19055 vdd.n2911 vdd.n443 9.3005
R19056 vdd.n2907 vdd.n2904 9.3005
R19057 vdd.n3021 vdd.n3020 9.3005
R19058 vdd.n2852 vdd.n2851 9.3005
R19059 vdd.n2853 vdd.n475 9.3005
R19060 vdd.n2855 vdd.n2854 9.3005
R19061 vdd.n465 vdd.n464 9.3005
R19062 vdd.n2869 vdd.n2868 9.3005
R19063 vdd.n2870 vdd.n463 9.3005
R19064 vdd.n2872 vdd.n2871 9.3005
R19065 vdd.n453 vdd.n452 9.3005
R19066 vdd.n2885 vdd.n2884 9.3005
R19067 vdd.n2886 vdd.n451 9.3005
R19068 vdd.n2888 vdd.n2887 9.3005
R19069 vdd.n2889 vdd.n450 9.3005
R19070 vdd.n2891 vdd.n2890 9.3005
R19071 vdd.n2892 vdd.n449 9.3005
R19072 vdd.n2894 vdd.n2893 9.3005
R19073 vdd.n2895 vdd.n447 9.3005
R19074 vdd.n2897 vdd.n2896 9.3005
R19075 vdd.n2898 vdd.n446 9.3005
R19076 vdd.n2900 vdd.n2899 9.3005
R19077 vdd.n2901 vdd.n444 9.3005
R19078 vdd.n2903 vdd.n2902 9.3005
R19079 vdd.n477 vdd.n476 9.3005
R19080 vdd.n2710 vdd.n2709 9.3005
R19081 vdd.n2715 vdd.n2708 9.3005
R19082 vdd.n2724 vdd.n572 9.3005
R19083 vdd.n2727 vdd.n571 9.3005
R19084 vdd.n2728 vdd.n570 9.3005
R19085 vdd.n2731 vdd.n569 9.3005
R19086 vdd.n2732 vdd.n568 9.3005
R19087 vdd.n2735 vdd.n567 9.3005
R19088 vdd.n2736 vdd.n566 9.3005
R19089 vdd.n2739 vdd.n565 9.3005
R19090 vdd.n2740 vdd.n564 9.3005
R19091 vdd.n2743 vdd.n563 9.3005
R19092 vdd.n2744 vdd.n562 9.3005
R19093 vdd.n2747 vdd.n561 9.3005
R19094 vdd.n2748 vdd.n560 9.3005
R19095 vdd.n2751 vdd.n559 9.3005
R19096 vdd.n2755 vdd.n2754 9.3005
R19097 vdd.n2756 vdd.n556 9.3005
R19098 vdd.n1951 vdd.n1950 9.3005
R19099 vdd.n1946 vdd.n857 9.3005
R19100 vdd.n1433 vdd.n1432 9.3005
R19101 vdd.n1434 vdd.n1188 9.3005
R19102 vdd.n1436 vdd.n1435 9.3005
R19103 vdd.n1178 vdd.n1177 9.3005
R19104 vdd.n1450 vdd.n1449 9.3005
R19105 vdd.n1451 vdd.n1176 9.3005
R19106 vdd.n1453 vdd.n1452 9.3005
R19107 vdd.n1168 vdd.n1167 9.3005
R19108 vdd.n1468 vdd.n1467 9.3005
R19109 vdd.n1469 vdd.n1166 9.3005
R19110 vdd.n1471 vdd.n1470 9.3005
R19111 vdd.n885 vdd.n884 9.3005
R19112 vdd.n1484 vdd.n1483 9.3005
R19113 vdd.n1485 vdd.n883 9.3005
R19114 vdd.n1487 vdd.n1486 9.3005
R19115 vdd.n875 vdd.n874 9.3005
R19116 vdd.n1501 vdd.n1500 9.3005
R19117 vdd.n1502 vdd.n872 9.3005
R19118 vdd.n1506 vdd.n1505 9.3005
R19119 vdd.n1504 vdd.n873 9.3005
R19120 vdd.n1503 vdd.n862 9.3005
R19121 vdd.n1190 vdd.n1189 9.3005
R19122 vdd.n1326 vdd.n1325 9.3005
R19123 vdd.n1327 vdd.n1316 9.3005
R19124 vdd.n1329 vdd.n1328 9.3005
R19125 vdd.n1330 vdd.n1315 9.3005
R19126 vdd.n1332 vdd.n1331 9.3005
R19127 vdd.n1333 vdd.n1310 9.3005
R19128 vdd.n1335 vdd.n1334 9.3005
R19129 vdd.n1336 vdd.n1309 9.3005
R19130 vdd.n1338 vdd.n1337 9.3005
R19131 vdd.n1339 vdd.n1304 9.3005
R19132 vdd.n1341 vdd.n1340 9.3005
R19133 vdd.n1342 vdd.n1303 9.3005
R19134 vdd.n1344 vdd.n1343 9.3005
R19135 vdd.n1345 vdd.n1298 9.3005
R19136 vdd.n1347 vdd.n1346 9.3005
R19137 vdd.n1348 vdd.n1297 9.3005
R19138 vdd.n1350 vdd.n1349 9.3005
R19139 vdd.n1351 vdd.n1292 9.3005
R19140 vdd.n1353 vdd.n1352 9.3005
R19141 vdd.n1354 vdd.n1291 9.3005
R19142 vdd.n1356 vdd.n1355 9.3005
R19143 vdd.n1360 vdd.n1287 9.3005
R19144 vdd.n1362 vdd.n1361 9.3005
R19145 vdd.n1363 vdd.n1286 9.3005
R19146 vdd.n1365 vdd.n1364 9.3005
R19147 vdd.n1366 vdd.n1281 9.3005
R19148 vdd.n1368 vdd.n1367 9.3005
R19149 vdd.n1369 vdd.n1280 9.3005
R19150 vdd.n1371 vdd.n1370 9.3005
R19151 vdd.n1372 vdd.n1275 9.3005
R19152 vdd.n1374 vdd.n1373 9.3005
R19153 vdd.n1375 vdd.n1274 9.3005
R19154 vdd.n1377 vdd.n1376 9.3005
R19155 vdd.n1378 vdd.n1269 9.3005
R19156 vdd.n1380 vdd.n1379 9.3005
R19157 vdd.n1381 vdd.n1268 9.3005
R19158 vdd.n1383 vdd.n1382 9.3005
R19159 vdd.n1384 vdd.n1263 9.3005
R19160 vdd.n1386 vdd.n1385 9.3005
R19161 vdd.n1387 vdd.n1262 9.3005
R19162 vdd.n1389 vdd.n1388 9.3005
R19163 vdd.n1390 vdd.n1257 9.3005
R19164 vdd.n1392 vdd.n1391 9.3005
R19165 vdd.n1393 vdd.n1256 9.3005
R19166 vdd.n1395 vdd.n1394 9.3005
R19167 vdd.n1396 vdd.n1249 9.3005
R19168 vdd.n1398 vdd.n1397 9.3005
R19169 vdd.n1399 vdd.n1248 9.3005
R19170 vdd.n1401 vdd.n1400 9.3005
R19171 vdd.n1402 vdd.n1243 9.3005
R19172 vdd.n1404 vdd.n1403 9.3005
R19173 vdd.n1405 vdd.n1242 9.3005
R19174 vdd.n1407 vdd.n1406 9.3005
R19175 vdd.n1408 vdd.n1237 9.3005
R19176 vdd.n1410 vdd.n1409 9.3005
R19177 vdd.n1411 vdd.n1236 9.3005
R19178 vdd.n1413 vdd.n1412 9.3005
R19179 vdd.n1414 vdd.n1231 9.3005
R19180 vdd.n1416 vdd.n1415 9.3005
R19181 vdd.n1417 vdd.n1230 9.3005
R19182 vdd.n1419 vdd.n1418 9.3005
R19183 vdd.n1195 vdd.n1194 9.3005
R19184 vdd.n1425 vdd.n1424 9.3005
R19185 vdd.n1324 vdd.n1323 9.3005
R19186 vdd.n1428 vdd.n1427 9.3005
R19187 vdd.n1184 vdd.n1183 9.3005
R19188 vdd.n1442 vdd.n1441 9.3005
R19189 vdd.n1443 vdd.n1182 9.3005
R19190 vdd.n1445 vdd.n1444 9.3005
R19191 vdd.n1173 vdd.n1172 9.3005
R19192 vdd.n1459 vdd.n1458 9.3005
R19193 vdd.n1460 vdd.n1171 9.3005
R19194 vdd.n1463 vdd.n1462 9.3005
R19195 vdd.n1461 vdd.n1162 9.3005
R19196 vdd.n1426 vdd.n1193 9.3005
R19197 vdd.n1086 vdd.n1085 9.3005
R19198 vdd.n1081 vdd.n1080 9.3005
R19199 vdd.n1092 vdd.n1091 9.3005
R19200 vdd.n1094 vdd.n1093 9.3005
R19201 vdd.n1077 vdd.n1076 9.3005
R19202 vdd.n1100 vdd.n1099 9.3005
R19203 vdd.n1102 vdd.n1101 9.3005
R19204 vdd.n1074 vdd.n1071 9.3005
R19205 vdd.n1109 vdd.n1108 9.3005
R19206 vdd.n1133 vdd.n1132 9.3005
R19207 vdd.n1128 vdd.n1127 9.3005
R19208 vdd.n1139 vdd.n1138 9.3005
R19209 vdd.n1141 vdd.n1140 9.3005
R19210 vdd.n1124 vdd.n1123 9.3005
R19211 vdd.n1147 vdd.n1146 9.3005
R19212 vdd.n1149 vdd.n1148 9.3005
R19213 vdd.n1121 vdd.n1118 9.3005
R19214 vdd.n1156 vdd.n1155 9.3005
R19215 vdd.n996 vdd.n995 9.3005
R19216 vdd.n991 vdd.n990 9.3005
R19217 vdd.n1002 vdd.n1001 9.3005
R19218 vdd.n1004 vdd.n1003 9.3005
R19219 vdd.n987 vdd.n986 9.3005
R19220 vdd.n1010 vdd.n1009 9.3005
R19221 vdd.n1012 vdd.n1011 9.3005
R19222 vdd.n984 vdd.n981 9.3005
R19223 vdd.n1019 vdd.n1018 9.3005
R19224 vdd.n1043 vdd.n1042 9.3005
R19225 vdd.n1038 vdd.n1037 9.3005
R19226 vdd.n1049 vdd.n1048 9.3005
R19227 vdd.n1051 vdd.n1050 9.3005
R19228 vdd.n1034 vdd.n1033 9.3005
R19229 vdd.n1057 vdd.n1056 9.3005
R19230 vdd.n1059 vdd.n1058 9.3005
R19231 vdd.n1031 vdd.n1028 9.3005
R19232 vdd.n1066 vdd.n1065 9.3005
R19233 vdd.n907 vdd.n906 9.3005
R19234 vdd.n902 vdd.n901 9.3005
R19235 vdd.n913 vdd.n912 9.3005
R19236 vdd.n915 vdd.n914 9.3005
R19237 vdd.n898 vdd.n897 9.3005
R19238 vdd.n921 vdd.n920 9.3005
R19239 vdd.n923 vdd.n922 9.3005
R19240 vdd.n895 vdd.n892 9.3005
R19241 vdd.n930 vdd.n929 9.3005
R19242 vdd.n954 vdd.n953 9.3005
R19243 vdd.n949 vdd.n948 9.3005
R19244 vdd.n960 vdd.n959 9.3005
R19245 vdd.n962 vdd.n961 9.3005
R19246 vdd.n945 vdd.n944 9.3005
R19247 vdd.n968 vdd.n967 9.3005
R19248 vdd.n970 vdd.n969 9.3005
R19249 vdd.n942 vdd.n939 9.3005
R19250 vdd.n977 vdd.n976 9.3005
R19251 vdd.n1438 vdd.t149 8.95635
R19252 vdd.t131 vdd.n3033 8.95635
R19253 vdd.n276 vdd.n275 8.92171
R19254 vdd.n229 vdd.n228 8.92171
R19255 vdd.n186 vdd.n185 8.92171
R19256 vdd.n139 vdd.n138 8.92171
R19257 vdd.n97 vdd.n96 8.92171
R19258 vdd.n50 vdd.n49 8.92171
R19259 vdd.n1091 vdd.n1090 8.92171
R19260 vdd.n1138 vdd.n1137 8.92171
R19261 vdd.n1001 vdd.n1000 8.92171
R19262 vdd.n1048 vdd.n1047 8.92171
R19263 vdd.n912 vdd.n911 8.92171
R19264 vdd.n959 vdd.n958 8.92171
R19265 vdd.n207 vdd.n117 8.81535
R19266 vdd.n1069 vdd.n979 8.81535
R19267 vdd.n1465 vdd.t127 8.72962
R19268 vdd.t129 vdd.n3042 8.72962
R19269 vdd.n888 vdd.t165 8.50289
R19270 vdd.n1943 vdd.t22 8.50289
R19271 vdd.n516 vdd.t15 8.50289
R19272 vdd.n2874 vdd.t143 8.50289
R19273 vdd.n28 vdd.n14 8.42249
R19274 vdd.n3048 vdd.n3047 8.16225
R19275 vdd.n1161 vdd.n1160 8.16225
R19276 vdd.n272 vdd.n266 8.14595
R19277 vdd.n225 vdd.n219 8.14595
R19278 vdd.n182 vdd.n176 8.14595
R19279 vdd.n135 vdd.n129 8.14595
R19280 vdd.n93 vdd.n87 8.14595
R19281 vdd.n46 vdd.n40 8.14595
R19282 vdd.n1087 vdd.n1081 8.14595
R19283 vdd.n1134 vdd.n1128 8.14595
R19284 vdd.n997 vdd.n991 8.14595
R19285 vdd.n1044 vdd.n1038 8.14595
R19286 vdd.n908 vdd.n902 8.14595
R19287 vdd.n955 vdd.n949 8.14595
R19288 vdd.n2537 vdd.n639 8.11757
R19289 vdd.n2011 vdd.n2010 8.11757
R19290 vdd.n1989 vdd.n833 7.70933
R19291 vdd.n1995 vdd.n833 7.70933
R19292 vdd.n2001 vdd.n827 7.70933
R19293 vdd.n2001 vdd.n820 7.70933
R19294 vdd.n2007 vdd.n820 7.70933
R19295 vdd.n2007 vdd.n823 7.70933
R19296 vdd.n2014 vdd.n808 7.70933
R19297 vdd.n2020 vdd.n808 7.70933
R19298 vdd.n2026 vdd.n802 7.70933
R19299 vdd.n2032 vdd.n798 7.70933
R19300 vdd.n2038 vdd.n792 7.70933
R19301 vdd.n2050 vdd.n779 7.70933
R19302 vdd.n2056 vdd.n773 7.70933
R19303 vdd.n2056 vdd.n766 7.70933
R19304 vdd.n2064 vdd.n766 7.70933
R19305 vdd.n2071 vdd.t91 7.70933
R19306 vdd.n2146 vdd.t91 7.70933
R19307 vdd.n2478 vdd.t3 7.70933
R19308 vdd.n2484 vdd.t3 7.70933
R19309 vdd.n2490 vdd.n687 7.70933
R19310 vdd.n2496 vdd.n687 7.70933
R19311 vdd.n2496 vdd.n690 7.70933
R19312 vdd.n2502 vdd.n683 7.70933
R19313 vdd.n2514 vdd.n670 7.70933
R19314 vdd.n2520 vdd.n664 7.70933
R19315 vdd.n2526 vdd.n660 7.70933
R19316 vdd.n2532 vdd.n647 7.70933
R19317 vdd.n2540 vdd.n647 7.70933
R19318 vdd.n2546 vdd.n641 7.70933
R19319 vdd.n2546 vdd.n633 7.70933
R19320 vdd.n2597 vdd.n633 7.70933
R19321 vdd.n2597 vdd.n636 7.70933
R19322 vdd.n2603 vdd.n595 7.70933
R19323 vdd.n2673 vdd.n595 7.70933
R19324 vdd.n271 vdd.n268 7.3702
R19325 vdd.n224 vdd.n221 7.3702
R19326 vdd.n181 vdd.n178 7.3702
R19327 vdd.n134 vdd.n131 7.3702
R19328 vdd.n92 vdd.n89 7.3702
R19329 vdd.n45 vdd.n42 7.3702
R19330 vdd.n1086 vdd.n1083 7.3702
R19331 vdd.n1133 vdd.n1130 7.3702
R19332 vdd.n996 vdd.n993 7.3702
R19333 vdd.n1043 vdd.n1040 7.3702
R19334 vdd.n907 vdd.n904 7.3702
R19335 vdd.n954 vdd.n951 7.3702
R19336 vdd.n1361 vdd.n1360 6.98232
R19337 vdd.n1653 vdd.n1652 6.98232
R19338 vdd.n2950 vdd.n2949 6.98232
R19339 vdd.n2761 vdd.n2758 6.98232
R19340 vdd.n1498 vdd.t112 6.68904
R19341 vdd.n2857 vdd.t114 6.68904
R19342 vdd.t151 vdd.n887 6.46231
R19343 vdd.n2882 vdd.t118 6.46231
R19344 vdd.n1456 vdd.t133 6.23558
R19345 vdd.t122 vdd.n308 6.23558
R19346 vdd.n3048 vdd.n297 6.22547
R19347 vdd.n1160 vdd.n1159 6.22547
R19348 vdd.n2026 vdd.t109 6.00885
R19349 vdd.n2526 vdd.t90 6.00885
R19350 vdd.n823 vdd.t66 5.89549
R19351 vdd.t30 vdd.n641 5.89549
R19352 vdd.n272 vdd.n271 5.81868
R19353 vdd.n225 vdd.n224 5.81868
R19354 vdd.n182 vdd.n181 5.81868
R19355 vdd.n135 vdd.n134 5.81868
R19356 vdd.n93 vdd.n92 5.81868
R19357 vdd.n46 vdd.n45 5.81868
R19358 vdd.n1087 vdd.n1086 5.81868
R19359 vdd.n1134 vdd.n1133 5.81868
R19360 vdd.n997 vdd.n996 5.81868
R19361 vdd.n1044 vdd.n1043 5.81868
R19362 vdd.n908 vdd.n907 5.81868
R19363 vdd.n955 vdd.n954 5.81868
R19364 vdd.t62 vdd.n827 5.78212
R19365 vdd.n1770 vdd.t47 5.78212
R19366 vdd.n2395 vdd.t55 5.78212
R19367 vdd.n636 vdd.t51 5.78212
R19368 vdd.n2154 vdd.n2153 5.77611
R19369 vdd.n1897 vdd.n1767 5.77611
R19370 vdd.n2408 vdd.n2407 5.77611
R19371 vdd.n2614 vdd.n2613 5.77611
R19372 vdd.n2678 vdd.n591 5.77611
R19373 vdd.n2318 vdd.n2258 5.77611
R19374 vdd.n2079 vdd.n757 5.77611
R19375 vdd.n1827 vdd.n1826 5.77611
R19376 vdd.n1323 vdd.n1322 5.62474
R19377 vdd.n1949 vdd.n1946 5.62474
R19378 vdd.n2910 vdd.n2907 5.62474
R19379 vdd.n2713 vdd.n2710 5.62474
R19380 vdd.t93 vdd.n779 5.44203
R19381 vdd.n683 vdd.t196 5.44203
R19382 vdd.n1180 vdd.t133 5.10193
R19383 vdd.t104 vdd.n802 5.10193
R19384 vdd.n792 vdd.t2 5.10193
R19385 vdd.t10 vdd.n670 5.10193
R19386 vdd.n660 vdd.t103 5.10193
R19387 vdd.n3035 vdd.t122 5.10193
R19388 vdd.n275 vdd.n266 5.04292
R19389 vdd.n228 vdd.n219 5.04292
R19390 vdd.n185 vdd.n176 5.04292
R19391 vdd.n138 vdd.n129 5.04292
R19392 vdd.n96 vdd.n87 5.04292
R19393 vdd.n49 vdd.n40 5.04292
R19394 vdd.n1090 vdd.n1081 5.04292
R19395 vdd.n1137 vdd.n1128 5.04292
R19396 vdd.n1000 vdd.n991 5.04292
R19397 vdd.n1047 vdd.n1038 5.04292
R19398 vdd.n911 vdd.n902 5.04292
R19399 vdd.n958 vdd.n949 5.04292
R19400 vdd.n1473 vdd.t151 4.8752
R19401 vdd.t7 vdd.t101 4.8752
R19402 vdd.t110 vdd.t198 4.8752
R19403 vdd.t0 vdd.t13 4.8752
R19404 vdd.t95 vdd.t111 4.8752
R19405 vdd.t118 vdd.n304 4.8752
R19406 vdd.n2155 vdd.n2154 4.83952
R19407 vdd.n1767 vdd.n1763 4.83952
R19408 vdd.n2409 vdd.n2408 4.83952
R19409 vdd.n2615 vdd.n2614 4.83952
R19410 vdd.n591 vdd.n586 4.83952
R19411 vdd.n2315 vdd.n2258 4.83952
R19412 vdd.n2082 vdd.n757 4.83952
R19413 vdd.n1826 vdd.n1825 4.83952
R19414 vdd.n1621 vdd.n855 4.74817
R19415 vdd.n1616 vdd.n856 4.74817
R19416 vdd.n1518 vdd.n1515 4.74817
R19417 vdd.n1930 vdd.n1519 4.74817
R19418 vdd.n1932 vdd.n1518 4.74817
R19419 vdd.n1931 vdd.n1930 4.74817
R19420 vdd.n2838 vdd.n2837 4.74817
R19421 vdd.n2835 vdd.n2834 4.74817
R19422 vdd.n2835 vdd.n521 4.74817
R19423 vdd.n2837 vdd.n518 4.74817
R19424 vdd.n2720 vdd.n573 4.74817
R19425 vdd.n2716 vdd.n574 4.74817
R19426 vdd.n2719 vdd.n574 4.74817
R19427 vdd.n2723 vdd.n573 4.74817
R19428 vdd.n1617 vdd.n855 4.74817
R19429 vdd.n858 vdd.n856 4.74817
R19430 vdd.n297 vdd.n296 4.7074
R19431 vdd.n207 vdd.n206 4.7074
R19432 vdd.n1159 vdd.n1158 4.7074
R19433 vdd.n1069 vdd.n1068 4.7074
R19434 vdd.n1489 vdd.t112 4.64847
R19435 vdd.n2866 vdd.t114 4.64847
R19436 vdd.n2032 vdd.t8 4.53511
R19437 vdd.n2520 vdd.t107 4.53511
R19438 vdd.n2064 vdd.t105 4.30838
R19439 vdd.n2490 vdd.t11 4.30838
R19440 vdd.n276 vdd.n264 4.26717
R19441 vdd.n229 vdd.n217 4.26717
R19442 vdd.n186 vdd.n174 4.26717
R19443 vdd.n139 vdd.n127 4.26717
R19444 vdd.n97 vdd.n85 4.26717
R19445 vdd.n50 vdd.n38 4.26717
R19446 vdd.n1091 vdd.n1079 4.26717
R19447 vdd.n1138 vdd.n1126 4.26717
R19448 vdd.n1001 vdd.n989 4.26717
R19449 vdd.n1048 vdd.n1036 4.26717
R19450 vdd.n912 vdd.n900 4.26717
R19451 vdd.n959 vdd.n947 4.26717
R19452 vdd.n297 vdd.n207 4.10845
R19453 vdd.n1159 vdd.n1069 4.10845
R19454 vdd.n253 vdd.t159 4.06363
R19455 vdd.n253 vdd.t123 4.06363
R19456 vdd.n251 vdd.t125 4.06363
R19457 vdd.n251 vdd.t146 4.06363
R19458 vdd.n249 vdd.t148 4.06363
R19459 vdd.n249 vdd.t164 4.06363
R19460 vdd.n163 vdd.t154 4.06363
R19461 vdd.n163 vdd.t175 4.06363
R19462 vdd.n161 vdd.t119 4.06363
R19463 vdd.n161 vdd.t138 4.06363
R19464 vdd.n159 vdd.t144 4.06363
R19465 vdd.n159 vdd.t155 4.06363
R19466 vdd.n74 vdd.t160 4.06363
R19467 vdd.n74 vdd.t135 4.06363
R19468 vdd.n72 vdd.t174 4.06363
R19469 vdd.n72 vdd.t130 4.06363
R19470 vdd.n70 vdd.t167 4.06363
R19471 vdd.n70 vdd.t141 4.06363
R19472 vdd.n1111 vdd.t126 4.06363
R19473 vdd.n1111 vdd.t170 4.06363
R19474 vdd.n1113 vdd.t169 4.06363
R19475 vdd.n1113 vdd.t158 4.06363
R19476 vdd.n1115 vdd.t145 4.06363
R19477 vdd.n1115 vdd.t124 4.06363
R19478 vdd.n1021 vdd.t121 4.06363
R19479 vdd.n1021 vdd.t166 4.06363
R19480 vdd.n1023 vdd.t161 4.06363
R19481 vdd.n1023 vdd.t152 4.06363
R19482 vdd.n1025 vdd.t137 4.06363
R19483 vdd.n1025 vdd.t117 4.06363
R19484 vdd.n932 vdd.t139 4.06363
R19485 vdd.n932 vdd.t168 4.06363
R19486 vdd.n934 vdd.t128 4.06363
R19487 vdd.n934 vdd.t156 4.06363
R19488 vdd.n936 vdd.t134 4.06363
R19489 vdd.n936 vdd.t162 4.06363
R19490 vdd.n26 vdd.t183 3.9605
R19491 vdd.n26 vdd.t185 3.9605
R19492 vdd.n23 vdd.t184 3.9605
R19493 vdd.n23 vdd.t180 3.9605
R19494 vdd.n21 vdd.t190 3.9605
R19495 vdd.n21 vdd.t186 3.9605
R19496 vdd.n20 vdd.t176 3.9605
R19497 vdd.n20 vdd.t181 3.9605
R19498 vdd.n15 vdd.t177 3.9605
R19499 vdd.n15 vdd.t187 3.9605
R19500 vdd.n16 vdd.t188 3.9605
R19501 vdd.n16 vdd.t182 3.9605
R19502 vdd.n18 vdd.t179 3.9605
R19503 vdd.n18 vdd.t189 3.9605
R19504 vdd.n25 vdd.t178 3.9605
R19505 vdd.n25 vdd.t191 3.9605
R19506 vdd.n7 vdd.t96 3.61217
R19507 vdd.n7 vdd.t108 3.61217
R19508 vdd.n8 vdd.t1 3.61217
R19509 vdd.n8 vdd.t197 3.61217
R19510 vdd.n10 vdd.t4 3.61217
R19511 vdd.n10 vdd.t12 3.61217
R19512 vdd.n12 vdd.t99 3.61217
R19513 vdd.n12 vdd.t6 3.61217
R19514 vdd.n5 vdd.t195 3.61217
R19515 vdd.n5 vdd.t193 3.61217
R19516 vdd.n3 vdd.t106 3.61217
R19517 vdd.n3 vdd.t92 3.61217
R19518 vdd.n1 vdd.t94 3.61217
R19519 vdd.n1 vdd.t199 3.61217
R19520 vdd.n0 vdd.t9 3.61217
R19521 vdd.n0 vdd.t102 3.61217
R19522 vdd.n280 vdd.n279 3.49141
R19523 vdd.n233 vdd.n232 3.49141
R19524 vdd.n190 vdd.n189 3.49141
R19525 vdd.n143 vdd.n142 3.49141
R19526 vdd.n101 vdd.n100 3.49141
R19527 vdd.n54 vdd.n53 3.49141
R19528 vdd.n1095 vdd.n1094 3.49141
R19529 vdd.n1142 vdd.n1141 3.49141
R19530 vdd.n1005 vdd.n1004 3.49141
R19531 vdd.n1052 vdd.n1051 3.49141
R19532 vdd.n916 vdd.n915 3.49141
R19533 vdd.n963 vdd.n962 3.49141
R19534 vdd.n1770 vdd.t105 3.40145
R19535 vdd.n2218 vdd.t194 3.40145
R19536 vdd.n2471 vdd.t5 3.40145
R19537 vdd.n2395 vdd.t11 3.40145
R19538 vdd.n1871 vdd.t8 3.17472
R19539 vdd.n2374 vdd.t107 3.17472
R19540 vdd.n1490 vdd.t165 2.83463
R19541 vdd.n1508 vdd.t22 2.83463
R19542 vdd.n2849 vdd.t15 2.83463
R19543 vdd.n467 vdd.t143 2.83463
R19544 vdd.n283 vdd.n262 2.71565
R19545 vdd.n236 vdd.n215 2.71565
R19546 vdd.n193 vdd.n172 2.71565
R19547 vdd.n146 vdd.n125 2.71565
R19548 vdd.n104 vdd.n83 2.71565
R19549 vdd.n57 vdd.n36 2.71565
R19550 vdd.n1098 vdd.n1077 2.71565
R19551 vdd.n1145 vdd.n1124 2.71565
R19552 vdd.n1008 vdd.n987 2.71565
R19553 vdd.n1055 vdd.n1034 2.71565
R19554 vdd.n919 vdd.n898 2.71565
R19555 vdd.n966 vdd.n945 2.71565
R19556 vdd.t127 vdd.n1164 2.6079
R19557 vdd.n2020 vdd.t104 2.6079
R19558 vdd.n2044 vdd.t2 2.6079
R19559 vdd.n2508 vdd.t10 2.6079
R19560 vdd.n2532 vdd.t103 2.6079
R19561 vdd.n3043 vdd.t129 2.6079
R19562 vdd.n2538 vdd.n2537 2.49806
R19563 vdd.n2012 vdd.n2011 2.49806
R19564 vdd.n270 vdd.n269 2.4129
R19565 vdd.n223 vdd.n222 2.4129
R19566 vdd.n180 vdd.n179 2.4129
R19567 vdd.n133 vdd.n132 2.4129
R19568 vdd.n91 vdd.n90 2.4129
R19569 vdd.n44 vdd.n43 2.4129
R19570 vdd.n1085 vdd.n1084 2.4129
R19571 vdd.n1132 vdd.n1131 2.4129
R19572 vdd.n995 vdd.n994 2.4129
R19573 vdd.n1042 vdd.n1041 2.4129
R19574 vdd.n906 vdd.n905 2.4129
R19575 vdd.n953 vdd.n952 2.4129
R19576 vdd.n1447 vdd.t149 2.38117
R19577 vdd.n3034 vdd.t131 2.38117
R19578 vdd.n1929 vdd.n1518 2.27742
R19579 vdd.n1930 vdd.n1929 2.27742
R19580 vdd.n2836 vdd.n2835 2.27742
R19581 vdd.n2837 vdd.n2836 2.27742
R19582 vdd.n2707 vdd.n574 2.27742
R19583 vdd.n2707 vdd.n573 2.27742
R19584 vdd.n1952 vdd.n855 2.27742
R19585 vdd.n1952 vdd.n856 2.27742
R19586 vdd.n2044 vdd.t93 2.2678
R19587 vdd.n2508 vdd.t196 2.2678
R19588 vdd.t198 vdd.n773 2.04107
R19589 vdd.n690 vdd.t0 2.04107
R19590 vdd.n284 vdd.n260 1.93989
R19591 vdd.n237 vdd.n213 1.93989
R19592 vdd.n194 vdd.n170 1.93989
R19593 vdd.n147 vdd.n123 1.93989
R19594 vdd.n105 vdd.n81 1.93989
R19595 vdd.n58 vdd.n34 1.93989
R19596 vdd.n1099 vdd.n1075 1.93989
R19597 vdd.n1146 vdd.n1122 1.93989
R19598 vdd.n1009 vdd.n985 1.93989
R19599 vdd.n1056 vdd.n1032 1.93989
R19600 vdd.n920 vdd.n896 1.93989
R19601 vdd.n967 vdd.n943 1.93989
R19602 vdd.n1995 vdd.t62 1.92771
R19603 vdd.n2071 vdd.t47 1.92771
R19604 vdd.n2484 vdd.t55 1.92771
R19605 vdd.n2603 vdd.t51 1.92771
R19606 vdd.n1871 vdd.t109 1.70098
R19607 vdd.n798 vdd.t7 1.70098
R19608 vdd.t111 vdd.n664 1.70098
R19609 vdd.n2374 vdd.t90 1.70098
R19610 vdd.n1455 vdd.t116 1.24752
R19611 vdd.t153 vdd.n3041 1.24752
R19612 vdd.n295 vdd.n255 1.16414
R19613 vdd.n288 vdd.n287 1.16414
R19614 vdd.n248 vdd.n208 1.16414
R19615 vdd.n241 vdd.n240 1.16414
R19616 vdd.n205 vdd.n165 1.16414
R19617 vdd.n198 vdd.n197 1.16414
R19618 vdd.n158 vdd.n118 1.16414
R19619 vdd.n151 vdd.n150 1.16414
R19620 vdd.n116 vdd.n76 1.16414
R19621 vdd.n109 vdd.n108 1.16414
R19622 vdd.n69 vdd.n29 1.16414
R19623 vdd.n62 vdd.n61 1.16414
R19624 vdd.n1110 vdd.n1070 1.16414
R19625 vdd.n1103 vdd.n1102 1.16414
R19626 vdd.n1157 vdd.n1117 1.16414
R19627 vdd.n1150 vdd.n1149 1.16414
R19628 vdd.n1020 vdd.n980 1.16414
R19629 vdd.n1013 vdd.n1012 1.16414
R19630 vdd.n1067 vdd.n1027 1.16414
R19631 vdd.n1060 vdd.n1059 1.16414
R19632 vdd.n931 vdd.n891 1.16414
R19633 vdd.n924 vdd.n923 1.16414
R19634 vdd.n978 vdd.n938 1.16414
R19635 vdd.n971 vdd.n970 1.16414
R19636 vdd.n2038 vdd.t101 1.13415
R19637 vdd.n2514 vdd.t95 1.13415
R19638 vdd.n1481 vdd.t120 1.02079
R19639 vdd.t66 vdd.t97 1.02079
R19640 vdd.t100 vdd.t30 1.02079
R19641 vdd.t140 vdd.n456 1.02079
R19642 vdd.n1326 vdd.n1322 0.970197
R19643 vdd.n1950 vdd.n1949 0.970197
R19644 vdd.n2911 vdd.n2910 0.970197
R19645 vdd.n2715 vdd.n2713 0.970197
R19646 vdd.n2014 vdd.t97 0.794056
R19647 vdd.n2050 vdd.t110 0.794056
R19648 vdd.n2502 vdd.t13 0.794056
R19649 vdd.n2540 vdd.t100 0.794056
R19650 vdd.n1160 vdd.n28 0.74827
R19651 vdd vdd.n3048 0.740437
R19652 vdd.n1430 vdd.t26 0.567326
R19653 vdd.n3026 vdd.t37 0.567326
R19654 vdd.n1940 vdd.n1939 0.537085
R19655 vdd.n2845 vdd.n2844 0.537085
R19656 vdd.n3022 vdd.n3021 0.537085
R19657 vdd.n2904 vdd.n2903 0.537085
R19658 vdd.n2709 vdd.n476 0.537085
R19659 vdd.n1503 vdd.n857 0.537085
R19660 vdd.n1324 vdd.n1189 0.537085
R19661 vdd.n1426 vdd.n1425 0.537085
R19662 vdd.n4 vdd.n2 0.459552
R19663 vdd.n11 vdd.n9 0.459552
R19664 vdd.n293 vdd.n292 0.388379
R19665 vdd.n259 vdd.n257 0.388379
R19666 vdd.n246 vdd.n245 0.388379
R19667 vdd.n212 vdd.n210 0.388379
R19668 vdd.n203 vdd.n202 0.388379
R19669 vdd.n169 vdd.n167 0.388379
R19670 vdd.n156 vdd.n155 0.388379
R19671 vdd.n122 vdd.n120 0.388379
R19672 vdd.n114 vdd.n113 0.388379
R19673 vdd.n80 vdd.n78 0.388379
R19674 vdd.n67 vdd.n66 0.388379
R19675 vdd.n33 vdd.n31 0.388379
R19676 vdd.n1108 vdd.n1107 0.388379
R19677 vdd.n1074 vdd.n1072 0.388379
R19678 vdd.n1155 vdd.n1154 0.388379
R19679 vdd.n1121 vdd.n1119 0.388379
R19680 vdd.n1018 vdd.n1017 0.388379
R19681 vdd.n984 vdd.n982 0.388379
R19682 vdd.n1065 vdd.n1064 0.388379
R19683 vdd.n1031 vdd.n1029 0.388379
R19684 vdd.n929 vdd.n928 0.388379
R19685 vdd.n895 vdd.n893 0.388379
R19686 vdd.n976 vdd.n975 0.388379
R19687 vdd.n942 vdd.n940 0.388379
R19688 vdd.n19 vdd.n17 0.387128
R19689 vdd.n24 vdd.n22 0.387128
R19690 vdd.n6 vdd.n4 0.358259
R19691 vdd.n13 vdd.n11 0.358259
R19692 vdd.n252 vdd.n250 0.358259
R19693 vdd.n254 vdd.n252 0.358259
R19694 vdd.n296 vdd.n254 0.358259
R19695 vdd.n162 vdd.n160 0.358259
R19696 vdd.n164 vdd.n162 0.358259
R19697 vdd.n206 vdd.n164 0.358259
R19698 vdd.n73 vdd.n71 0.358259
R19699 vdd.n75 vdd.n73 0.358259
R19700 vdd.n117 vdd.n75 0.358259
R19701 vdd.n1158 vdd.n1116 0.358259
R19702 vdd.n1116 vdd.n1114 0.358259
R19703 vdd.n1114 vdd.n1112 0.358259
R19704 vdd.n1068 vdd.n1026 0.358259
R19705 vdd.n1026 vdd.n1024 0.358259
R19706 vdd.n1024 vdd.n1022 0.358259
R19707 vdd.n979 vdd.n937 0.358259
R19708 vdd.n937 vdd.n935 0.358259
R19709 vdd.n935 vdd.n933 0.358259
R19710 vdd.n14 vdd.n6 0.334552
R19711 vdd.n14 vdd.n13 0.334552
R19712 vdd.n27 vdd.n19 0.21707
R19713 vdd.n27 vdd.n24 0.21707
R19714 vdd.n294 vdd.n256 0.155672
R19715 vdd.n286 vdd.n256 0.155672
R19716 vdd.n286 vdd.n285 0.155672
R19717 vdd.n285 vdd.n261 0.155672
R19718 vdd.n278 vdd.n261 0.155672
R19719 vdd.n278 vdd.n277 0.155672
R19720 vdd.n277 vdd.n265 0.155672
R19721 vdd.n270 vdd.n265 0.155672
R19722 vdd.n247 vdd.n209 0.155672
R19723 vdd.n239 vdd.n209 0.155672
R19724 vdd.n239 vdd.n238 0.155672
R19725 vdd.n238 vdd.n214 0.155672
R19726 vdd.n231 vdd.n214 0.155672
R19727 vdd.n231 vdd.n230 0.155672
R19728 vdd.n230 vdd.n218 0.155672
R19729 vdd.n223 vdd.n218 0.155672
R19730 vdd.n204 vdd.n166 0.155672
R19731 vdd.n196 vdd.n166 0.155672
R19732 vdd.n196 vdd.n195 0.155672
R19733 vdd.n195 vdd.n171 0.155672
R19734 vdd.n188 vdd.n171 0.155672
R19735 vdd.n188 vdd.n187 0.155672
R19736 vdd.n187 vdd.n175 0.155672
R19737 vdd.n180 vdd.n175 0.155672
R19738 vdd.n157 vdd.n119 0.155672
R19739 vdd.n149 vdd.n119 0.155672
R19740 vdd.n149 vdd.n148 0.155672
R19741 vdd.n148 vdd.n124 0.155672
R19742 vdd.n141 vdd.n124 0.155672
R19743 vdd.n141 vdd.n140 0.155672
R19744 vdd.n140 vdd.n128 0.155672
R19745 vdd.n133 vdd.n128 0.155672
R19746 vdd.n115 vdd.n77 0.155672
R19747 vdd.n107 vdd.n77 0.155672
R19748 vdd.n107 vdd.n106 0.155672
R19749 vdd.n106 vdd.n82 0.155672
R19750 vdd.n99 vdd.n82 0.155672
R19751 vdd.n99 vdd.n98 0.155672
R19752 vdd.n98 vdd.n86 0.155672
R19753 vdd.n91 vdd.n86 0.155672
R19754 vdd.n68 vdd.n30 0.155672
R19755 vdd.n60 vdd.n30 0.155672
R19756 vdd.n60 vdd.n59 0.155672
R19757 vdd.n59 vdd.n35 0.155672
R19758 vdd.n52 vdd.n35 0.155672
R19759 vdd.n52 vdd.n51 0.155672
R19760 vdd.n51 vdd.n39 0.155672
R19761 vdd.n44 vdd.n39 0.155672
R19762 vdd.n1109 vdd.n1071 0.155672
R19763 vdd.n1101 vdd.n1071 0.155672
R19764 vdd.n1101 vdd.n1100 0.155672
R19765 vdd.n1100 vdd.n1076 0.155672
R19766 vdd.n1093 vdd.n1076 0.155672
R19767 vdd.n1093 vdd.n1092 0.155672
R19768 vdd.n1092 vdd.n1080 0.155672
R19769 vdd.n1085 vdd.n1080 0.155672
R19770 vdd.n1156 vdd.n1118 0.155672
R19771 vdd.n1148 vdd.n1118 0.155672
R19772 vdd.n1148 vdd.n1147 0.155672
R19773 vdd.n1147 vdd.n1123 0.155672
R19774 vdd.n1140 vdd.n1123 0.155672
R19775 vdd.n1140 vdd.n1139 0.155672
R19776 vdd.n1139 vdd.n1127 0.155672
R19777 vdd.n1132 vdd.n1127 0.155672
R19778 vdd.n1019 vdd.n981 0.155672
R19779 vdd.n1011 vdd.n981 0.155672
R19780 vdd.n1011 vdd.n1010 0.155672
R19781 vdd.n1010 vdd.n986 0.155672
R19782 vdd.n1003 vdd.n986 0.155672
R19783 vdd.n1003 vdd.n1002 0.155672
R19784 vdd.n1002 vdd.n990 0.155672
R19785 vdd.n995 vdd.n990 0.155672
R19786 vdd.n1066 vdd.n1028 0.155672
R19787 vdd.n1058 vdd.n1028 0.155672
R19788 vdd.n1058 vdd.n1057 0.155672
R19789 vdd.n1057 vdd.n1033 0.155672
R19790 vdd.n1050 vdd.n1033 0.155672
R19791 vdd.n1050 vdd.n1049 0.155672
R19792 vdd.n1049 vdd.n1037 0.155672
R19793 vdd.n1042 vdd.n1037 0.155672
R19794 vdd.n930 vdd.n892 0.155672
R19795 vdd.n922 vdd.n892 0.155672
R19796 vdd.n922 vdd.n921 0.155672
R19797 vdd.n921 vdd.n897 0.155672
R19798 vdd.n914 vdd.n897 0.155672
R19799 vdd.n914 vdd.n913 0.155672
R19800 vdd.n913 vdd.n901 0.155672
R19801 vdd.n906 vdd.n901 0.155672
R19802 vdd.n977 vdd.n939 0.155672
R19803 vdd.n969 vdd.n939 0.155672
R19804 vdd.n969 vdd.n968 0.155672
R19805 vdd.n968 vdd.n944 0.155672
R19806 vdd.n961 vdd.n944 0.155672
R19807 vdd.n961 vdd.n960 0.155672
R19808 vdd.n960 vdd.n948 0.155672
R19809 vdd.n953 vdd.n948 0.155672
R19810 vdd.n1715 vdd.n1520 0.152939
R19811 vdd.n1526 vdd.n1520 0.152939
R19812 vdd.n1527 vdd.n1526 0.152939
R19813 vdd.n1528 vdd.n1527 0.152939
R19814 vdd.n1529 vdd.n1528 0.152939
R19815 vdd.n1533 vdd.n1529 0.152939
R19816 vdd.n1534 vdd.n1533 0.152939
R19817 vdd.n1535 vdd.n1534 0.152939
R19818 vdd.n1536 vdd.n1535 0.152939
R19819 vdd.n1540 vdd.n1536 0.152939
R19820 vdd.n1541 vdd.n1540 0.152939
R19821 vdd.n1542 vdd.n1541 0.152939
R19822 vdd.n1690 vdd.n1542 0.152939
R19823 vdd.n1690 vdd.n1689 0.152939
R19824 vdd.n1689 vdd.n1688 0.152939
R19825 vdd.n1688 vdd.n1548 0.152939
R19826 vdd.n1553 vdd.n1548 0.152939
R19827 vdd.n1554 vdd.n1553 0.152939
R19828 vdd.n1555 vdd.n1554 0.152939
R19829 vdd.n1559 vdd.n1555 0.152939
R19830 vdd.n1560 vdd.n1559 0.152939
R19831 vdd.n1561 vdd.n1560 0.152939
R19832 vdd.n1562 vdd.n1561 0.152939
R19833 vdd.n1566 vdd.n1562 0.152939
R19834 vdd.n1567 vdd.n1566 0.152939
R19835 vdd.n1568 vdd.n1567 0.152939
R19836 vdd.n1569 vdd.n1568 0.152939
R19837 vdd.n1573 vdd.n1569 0.152939
R19838 vdd.n1574 vdd.n1573 0.152939
R19839 vdd.n1575 vdd.n1574 0.152939
R19840 vdd.n1576 vdd.n1575 0.152939
R19841 vdd.n1580 vdd.n1576 0.152939
R19842 vdd.n1581 vdd.n1580 0.152939
R19843 vdd.n1582 vdd.n1581 0.152939
R19844 vdd.n1651 vdd.n1582 0.152939
R19845 vdd.n1651 vdd.n1650 0.152939
R19846 vdd.n1650 vdd.n1649 0.152939
R19847 vdd.n1649 vdd.n1588 0.152939
R19848 vdd.n1593 vdd.n1588 0.152939
R19849 vdd.n1594 vdd.n1593 0.152939
R19850 vdd.n1595 vdd.n1594 0.152939
R19851 vdd.n1599 vdd.n1595 0.152939
R19852 vdd.n1600 vdd.n1599 0.152939
R19853 vdd.n1601 vdd.n1600 0.152939
R19854 vdd.n1602 vdd.n1601 0.152939
R19855 vdd.n1606 vdd.n1602 0.152939
R19856 vdd.n1607 vdd.n1606 0.152939
R19857 vdd.n1608 vdd.n1607 0.152939
R19858 vdd.n1609 vdd.n1608 0.152939
R19859 vdd.n1610 vdd.n1609 0.152939
R19860 vdd.n1610 vdd.n854 0.152939
R19861 vdd.n1939 vdd.n1514 0.152939
R19862 vdd.n1477 vdd.n1476 0.152939
R19863 vdd.n1478 vdd.n1477 0.152939
R19864 vdd.n1478 vdd.n879 0.152939
R19865 vdd.n1493 vdd.n879 0.152939
R19866 vdd.n1494 vdd.n1493 0.152939
R19867 vdd.n1495 vdd.n1494 0.152939
R19868 vdd.n1495 vdd.n867 0.152939
R19869 vdd.n1512 vdd.n867 0.152939
R19870 vdd.n1513 vdd.n1512 0.152939
R19871 vdd.n1940 vdd.n1513 0.152939
R19872 vdd.n524 vdd.n519 0.152939
R19873 vdd.n525 vdd.n524 0.152939
R19874 vdd.n526 vdd.n525 0.152939
R19875 vdd.n527 vdd.n526 0.152939
R19876 vdd.n528 vdd.n527 0.152939
R19877 vdd.n529 vdd.n528 0.152939
R19878 vdd.n530 vdd.n529 0.152939
R19879 vdd.n531 vdd.n530 0.152939
R19880 vdd.n532 vdd.n531 0.152939
R19881 vdd.n533 vdd.n532 0.152939
R19882 vdd.n534 vdd.n533 0.152939
R19883 vdd.n535 vdd.n534 0.152939
R19884 vdd.n2803 vdd.n535 0.152939
R19885 vdd.n2803 vdd.n2802 0.152939
R19886 vdd.n2802 vdd.n2801 0.152939
R19887 vdd.n2801 vdd.n537 0.152939
R19888 vdd.n538 vdd.n537 0.152939
R19889 vdd.n539 vdd.n538 0.152939
R19890 vdd.n540 vdd.n539 0.152939
R19891 vdd.n541 vdd.n540 0.152939
R19892 vdd.n542 vdd.n541 0.152939
R19893 vdd.n543 vdd.n542 0.152939
R19894 vdd.n544 vdd.n543 0.152939
R19895 vdd.n545 vdd.n544 0.152939
R19896 vdd.n546 vdd.n545 0.152939
R19897 vdd.n547 vdd.n546 0.152939
R19898 vdd.n548 vdd.n547 0.152939
R19899 vdd.n549 vdd.n548 0.152939
R19900 vdd.n550 vdd.n549 0.152939
R19901 vdd.n551 vdd.n550 0.152939
R19902 vdd.n552 vdd.n551 0.152939
R19903 vdd.n553 vdd.n552 0.152939
R19904 vdd.n554 vdd.n553 0.152939
R19905 vdd.n555 vdd.n554 0.152939
R19906 vdd.n2757 vdd.n555 0.152939
R19907 vdd.n2757 vdd.n2756 0.152939
R19908 vdd.n2756 vdd.n2755 0.152939
R19909 vdd.n2755 vdd.n559 0.152939
R19910 vdd.n560 vdd.n559 0.152939
R19911 vdd.n561 vdd.n560 0.152939
R19912 vdd.n562 vdd.n561 0.152939
R19913 vdd.n563 vdd.n562 0.152939
R19914 vdd.n564 vdd.n563 0.152939
R19915 vdd.n565 vdd.n564 0.152939
R19916 vdd.n566 vdd.n565 0.152939
R19917 vdd.n567 vdd.n566 0.152939
R19918 vdd.n568 vdd.n567 0.152939
R19919 vdd.n569 vdd.n568 0.152939
R19920 vdd.n570 vdd.n569 0.152939
R19921 vdd.n571 vdd.n570 0.152939
R19922 vdd.n572 vdd.n571 0.152939
R19923 vdd.n2844 vdd.n481 0.152939
R19924 vdd.n2846 vdd.n2845 0.152939
R19925 vdd.n2846 vdd.n470 0.152939
R19926 vdd.n2861 vdd.n470 0.152939
R19927 vdd.n2862 vdd.n2861 0.152939
R19928 vdd.n2863 vdd.n2862 0.152939
R19929 vdd.n2863 vdd.n459 0.152939
R19930 vdd.n2877 vdd.n459 0.152939
R19931 vdd.n2878 vdd.n2877 0.152939
R19932 vdd.n2879 vdd.n2878 0.152939
R19933 vdd.n2879 vdd.n298 0.152939
R19934 vdd.n3046 vdd.n299 0.152939
R19935 vdd.n310 vdd.n299 0.152939
R19936 vdd.n311 vdd.n310 0.152939
R19937 vdd.n312 vdd.n311 0.152939
R19938 vdd.n320 vdd.n312 0.152939
R19939 vdd.n321 vdd.n320 0.152939
R19940 vdd.n322 vdd.n321 0.152939
R19941 vdd.n323 vdd.n322 0.152939
R19942 vdd.n331 vdd.n323 0.152939
R19943 vdd.n3022 vdd.n331 0.152939
R19944 vdd.n3021 vdd.n332 0.152939
R19945 vdd.n335 vdd.n332 0.152939
R19946 vdd.n339 vdd.n335 0.152939
R19947 vdd.n340 vdd.n339 0.152939
R19948 vdd.n341 vdd.n340 0.152939
R19949 vdd.n342 vdd.n341 0.152939
R19950 vdd.n343 vdd.n342 0.152939
R19951 vdd.n347 vdd.n343 0.152939
R19952 vdd.n348 vdd.n347 0.152939
R19953 vdd.n349 vdd.n348 0.152939
R19954 vdd.n350 vdd.n349 0.152939
R19955 vdd.n354 vdd.n350 0.152939
R19956 vdd.n355 vdd.n354 0.152939
R19957 vdd.n356 vdd.n355 0.152939
R19958 vdd.n357 vdd.n356 0.152939
R19959 vdd.n361 vdd.n357 0.152939
R19960 vdd.n362 vdd.n361 0.152939
R19961 vdd.n363 vdd.n362 0.152939
R19962 vdd.n2987 vdd.n363 0.152939
R19963 vdd.n2987 vdd.n2986 0.152939
R19964 vdd.n2986 vdd.n2985 0.152939
R19965 vdd.n2985 vdd.n369 0.152939
R19966 vdd.n374 vdd.n369 0.152939
R19967 vdd.n375 vdd.n374 0.152939
R19968 vdd.n376 vdd.n375 0.152939
R19969 vdd.n380 vdd.n376 0.152939
R19970 vdd.n381 vdd.n380 0.152939
R19971 vdd.n382 vdd.n381 0.152939
R19972 vdd.n383 vdd.n382 0.152939
R19973 vdd.n387 vdd.n383 0.152939
R19974 vdd.n388 vdd.n387 0.152939
R19975 vdd.n389 vdd.n388 0.152939
R19976 vdd.n390 vdd.n389 0.152939
R19977 vdd.n394 vdd.n390 0.152939
R19978 vdd.n395 vdd.n394 0.152939
R19979 vdd.n396 vdd.n395 0.152939
R19980 vdd.n397 vdd.n396 0.152939
R19981 vdd.n401 vdd.n397 0.152939
R19982 vdd.n402 vdd.n401 0.152939
R19983 vdd.n403 vdd.n402 0.152939
R19984 vdd.n2948 vdd.n403 0.152939
R19985 vdd.n2948 vdd.n2947 0.152939
R19986 vdd.n2947 vdd.n2946 0.152939
R19987 vdd.n2946 vdd.n409 0.152939
R19988 vdd.n414 vdd.n409 0.152939
R19989 vdd.n415 vdd.n414 0.152939
R19990 vdd.n416 vdd.n415 0.152939
R19991 vdd.n420 vdd.n416 0.152939
R19992 vdd.n421 vdd.n420 0.152939
R19993 vdd.n422 vdd.n421 0.152939
R19994 vdd.n423 vdd.n422 0.152939
R19995 vdd.n427 vdd.n423 0.152939
R19996 vdd.n428 vdd.n427 0.152939
R19997 vdd.n429 vdd.n428 0.152939
R19998 vdd.n430 vdd.n429 0.152939
R19999 vdd.n434 vdd.n430 0.152939
R20000 vdd.n435 vdd.n434 0.152939
R20001 vdd.n436 vdd.n435 0.152939
R20002 vdd.n437 vdd.n436 0.152939
R20003 vdd.n441 vdd.n437 0.152939
R20004 vdd.n442 vdd.n441 0.152939
R20005 vdd.n443 vdd.n442 0.152939
R20006 vdd.n2904 vdd.n443 0.152939
R20007 vdd.n2852 vdd.n476 0.152939
R20008 vdd.n2853 vdd.n2852 0.152939
R20009 vdd.n2854 vdd.n2853 0.152939
R20010 vdd.n2854 vdd.n464 0.152939
R20011 vdd.n2869 vdd.n464 0.152939
R20012 vdd.n2870 vdd.n2869 0.152939
R20013 vdd.n2871 vdd.n2870 0.152939
R20014 vdd.n2871 vdd.n452 0.152939
R20015 vdd.n2885 vdd.n452 0.152939
R20016 vdd.n2886 vdd.n2885 0.152939
R20017 vdd.n2887 vdd.n2886 0.152939
R20018 vdd.n2887 vdd.n450 0.152939
R20019 vdd.n2891 vdd.n450 0.152939
R20020 vdd.n2892 vdd.n2891 0.152939
R20021 vdd.n2893 vdd.n2892 0.152939
R20022 vdd.n2893 vdd.n447 0.152939
R20023 vdd.n2897 vdd.n447 0.152939
R20024 vdd.n2898 vdd.n2897 0.152939
R20025 vdd.n2899 vdd.n2898 0.152939
R20026 vdd.n2899 vdd.n444 0.152939
R20027 vdd.n2903 vdd.n444 0.152939
R20028 vdd.n2709 vdd.n2708 0.152939
R20029 vdd.n1951 vdd.n857 0.152939
R20030 vdd.n1433 vdd.n1189 0.152939
R20031 vdd.n1434 vdd.n1433 0.152939
R20032 vdd.n1435 vdd.n1434 0.152939
R20033 vdd.n1435 vdd.n1177 0.152939
R20034 vdd.n1450 vdd.n1177 0.152939
R20035 vdd.n1451 vdd.n1450 0.152939
R20036 vdd.n1452 vdd.n1451 0.152939
R20037 vdd.n1452 vdd.n1167 0.152939
R20038 vdd.n1468 vdd.n1167 0.152939
R20039 vdd.n1469 vdd.n1468 0.152939
R20040 vdd.n1470 vdd.n1469 0.152939
R20041 vdd.n1470 vdd.n884 0.152939
R20042 vdd.n1484 vdd.n884 0.152939
R20043 vdd.n1485 vdd.n1484 0.152939
R20044 vdd.n1486 vdd.n1485 0.152939
R20045 vdd.n1486 vdd.n874 0.152939
R20046 vdd.n1501 vdd.n874 0.152939
R20047 vdd.n1502 vdd.n1501 0.152939
R20048 vdd.n1505 vdd.n1502 0.152939
R20049 vdd.n1505 vdd.n1504 0.152939
R20050 vdd.n1504 vdd.n1503 0.152939
R20051 vdd.n1425 vdd.n1194 0.152939
R20052 vdd.n1418 vdd.n1194 0.152939
R20053 vdd.n1418 vdd.n1417 0.152939
R20054 vdd.n1417 vdd.n1416 0.152939
R20055 vdd.n1416 vdd.n1231 0.152939
R20056 vdd.n1412 vdd.n1231 0.152939
R20057 vdd.n1412 vdd.n1411 0.152939
R20058 vdd.n1411 vdd.n1410 0.152939
R20059 vdd.n1410 vdd.n1237 0.152939
R20060 vdd.n1406 vdd.n1237 0.152939
R20061 vdd.n1406 vdd.n1405 0.152939
R20062 vdd.n1405 vdd.n1404 0.152939
R20063 vdd.n1404 vdd.n1243 0.152939
R20064 vdd.n1400 vdd.n1243 0.152939
R20065 vdd.n1400 vdd.n1399 0.152939
R20066 vdd.n1399 vdd.n1398 0.152939
R20067 vdd.n1398 vdd.n1249 0.152939
R20068 vdd.n1394 vdd.n1249 0.152939
R20069 vdd.n1394 vdd.n1393 0.152939
R20070 vdd.n1393 vdd.n1392 0.152939
R20071 vdd.n1392 vdd.n1257 0.152939
R20072 vdd.n1388 vdd.n1257 0.152939
R20073 vdd.n1388 vdd.n1387 0.152939
R20074 vdd.n1387 vdd.n1386 0.152939
R20075 vdd.n1386 vdd.n1263 0.152939
R20076 vdd.n1382 vdd.n1263 0.152939
R20077 vdd.n1382 vdd.n1381 0.152939
R20078 vdd.n1381 vdd.n1380 0.152939
R20079 vdd.n1380 vdd.n1269 0.152939
R20080 vdd.n1376 vdd.n1269 0.152939
R20081 vdd.n1376 vdd.n1375 0.152939
R20082 vdd.n1375 vdd.n1374 0.152939
R20083 vdd.n1374 vdd.n1275 0.152939
R20084 vdd.n1370 vdd.n1275 0.152939
R20085 vdd.n1370 vdd.n1369 0.152939
R20086 vdd.n1369 vdd.n1368 0.152939
R20087 vdd.n1368 vdd.n1281 0.152939
R20088 vdd.n1364 vdd.n1281 0.152939
R20089 vdd.n1364 vdd.n1363 0.152939
R20090 vdd.n1363 vdd.n1362 0.152939
R20091 vdd.n1362 vdd.n1287 0.152939
R20092 vdd.n1355 vdd.n1287 0.152939
R20093 vdd.n1355 vdd.n1354 0.152939
R20094 vdd.n1354 vdd.n1353 0.152939
R20095 vdd.n1353 vdd.n1292 0.152939
R20096 vdd.n1349 vdd.n1292 0.152939
R20097 vdd.n1349 vdd.n1348 0.152939
R20098 vdd.n1348 vdd.n1347 0.152939
R20099 vdd.n1347 vdd.n1298 0.152939
R20100 vdd.n1343 vdd.n1298 0.152939
R20101 vdd.n1343 vdd.n1342 0.152939
R20102 vdd.n1342 vdd.n1341 0.152939
R20103 vdd.n1341 vdd.n1304 0.152939
R20104 vdd.n1337 vdd.n1304 0.152939
R20105 vdd.n1337 vdd.n1336 0.152939
R20106 vdd.n1336 vdd.n1335 0.152939
R20107 vdd.n1335 vdd.n1310 0.152939
R20108 vdd.n1331 vdd.n1310 0.152939
R20109 vdd.n1331 vdd.n1330 0.152939
R20110 vdd.n1330 vdd.n1329 0.152939
R20111 vdd.n1329 vdd.n1316 0.152939
R20112 vdd.n1325 vdd.n1316 0.152939
R20113 vdd.n1325 vdd.n1324 0.152939
R20114 vdd.n1427 vdd.n1426 0.152939
R20115 vdd.n1427 vdd.n1183 0.152939
R20116 vdd.n1442 vdd.n1183 0.152939
R20117 vdd.n1443 vdd.n1442 0.152939
R20118 vdd.n1444 vdd.n1443 0.152939
R20119 vdd.n1444 vdd.n1172 0.152939
R20120 vdd.n1459 vdd.n1172 0.152939
R20121 vdd.n1460 vdd.n1459 0.152939
R20122 vdd.n1462 vdd.n1460 0.152939
R20123 vdd.n1462 vdd.n1461 0.152939
R20124 vdd.n1929 vdd.n1514 0.110256
R20125 vdd.n2836 vdd.n481 0.110256
R20126 vdd.n2708 vdd.n2707 0.110256
R20127 vdd.n1952 vdd.n1951 0.110256
R20128 vdd.n1476 vdd.n1161 0.0695946
R20129 vdd.n3047 vdd.n298 0.0695946
R20130 vdd.n3047 vdd.n3046 0.0695946
R20131 vdd.n1461 vdd.n1161 0.0695946
R20132 vdd.n1929 vdd.n1715 0.0431829
R20133 vdd.n1952 vdd.n854 0.0431829
R20134 vdd.n2836 vdd.n519 0.0431829
R20135 vdd.n2707 vdd.n572 0.0431829
R20136 vdd vdd.n28 0.00833333
R20137 a_n2848_n452.n3 a_n2848_n452.t75 539.01
R20138 a_n2848_n452.n57 a_n2848_n452.t58 512.366
R20139 a_n2848_n452.n56 a_n2848_n452.t62 512.366
R20140 a_n2848_n452.n54 a_n2848_n452.t52 512.366
R20141 a_n2848_n452.n55 a_n2848_n452.t67 512.366
R20142 a_n2848_n452.n45 a_n2848_n452.t37 533.058
R20143 a_n2848_n452.n58 a_n2848_n452.t21 512.366
R20144 a_n2848_n452.n59 a_n2848_n452.t29 512.366
R20145 a_n2848_n452.n50 a_n2848_n452.t33 512.366
R20146 a_n2848_n452.n80 a_n2848_n452.t31 512.366
R20147 a_n2848_n452.n78 a_n2848_n452.t35 512.366
R20148 a_n2848_n452.n17 a_n2848_n452.t19 539.01
R20149 a_n2848_n452.n102 a_n2848_n452.t39 512.366
R20150 a_n2848_n452.n103 a_n2848_n452.t25 512.366
R20151 a_n2848_n452.n52 a_n2848_n452.t23 512.366
R20152 a_n2848_n452.n104 a_n2848_n452.t17 512.366
R20153 a_n2848_n452.n21 a_n2848_n452.t70 539.01
R20154 a_n2848_n452.n99 a_n2848_n452.t71 512.366
R20155 a_n2848_n452.n100 a_n2848_n452.t50 512.366
R20156 a_n2848_n452.n53 a_n2848_n452.t56 512.366
R20157 a_n2848_n452.n101 a_n2848_n452.t65 512.366
R20158 a_n2848_n452.n91 a_n2848_n452.t64 512.366
R20159 a_n2848_n452.n90 a_n2848_n452.t55 512.366
R20160 a_n2848_n452.n89 a_n2848_n452.t49 512.366
R20161 a_n2848_n452.n93 a_n2848_n452.t72 512.366
R20162 a_n2848_n452.n92 a_n2848_n452.t61 512.366
R20163 a_n2848_n452.n88 a_n2848_n452.t60 512.366
R20164 a_n2848_n452.n95 a_n2848_n452.t68 512.366
R20165 a_n2848_n452.n94 a_n2848_n452.t53 512.366
R20166 a_n2848_n452.n87 a_n2848_n452.t54 512.366
R20167 a_n2848_n452.n97 a_n2848_n452.t57 512.366
R20168 a_n2848_n452.n96 a_n2848_n452.t66 512.366
R20169 a_n2848_n452.n86 a_n2848_n452.t48 512.366
R20170 a_n2848_n452.n48 a_n2848_n452.n1 70.3058
R20171 a_n2848_n452.n49 a_n2848_n452.n5 70.1674
R20172 a_n2848_n452.n14 a_n2848_n452.n34 70.3058
R20173 a_n2848_n452.n18 a_n2848_n452.n31 70.3058
R20174 a_n2848_n452.n30 a_n2848_n452.n19 70.1674
R20175 a_n2848_n452.n30 a_n2848_n452.n53 20.9683
R20176 a_n2848_n452.n19 a_n2848_n452.n29 75.0448
R20177 a_n2848_n452.n100 a_n2848_n452.n29 11.2134
R20178 a_n2848_n452.n20 a_n2848_n452.n21 44.8194
R20179 a_n2848_n452.n33 a_n2848_n452.n15 70.1674
R20180 a_n2848_n452.n33 a_n2848_n452.n52 20.9683
R20181 a_n2848_n452.n15 a_n2848_n452.n32 75.0448
R20182 a_n2848_n452.n103 a_n2848_n452.n32 11.2134
R20183 a_n2848_n452.n16 a_n2848_n452.n17 44.8194
R20184 a_n2848_n452.n6 a_n2848_n452.n43 70.1674
R20185 a_n2848_n452.n8 a_n2848_n452.n40 70.1674
R20186 a_n2848_n452.n10 a_n2848_n452.n38 70.1674
R20187 a_n2848_n452.n12 a_n2848_n452.n36 70.1674
R20188 a_n2848_n452.n36 a_n2848_n452.n86 20.9683
R20189 a_n2848_n452.n35 a_n2848_n452.n13 75.0448
R20190 a_n2848_n452.n96 a_n2848_n452.n35 11.2134
R20191 a_n2848_n452.n13 a_n2848_n452.n97 161.3
R20192 a_n2848_n452.n38 a_n2848_n452.n87 20.9683
R20193 a_n2848_n452.n37 a_n2848_n452.n11 75.0448
R20194 a_n2848_n452.n94 a_n2848_n452.n37 11.2134
R20195 a_n2848_n452.n11 a_n2848_n452.n95 161.3
R20196 a_n2848_n452.n40 a_n2848_n452.n88 20.9683
R20197 a_n2848_n452.n39 a_n2848_n452.n9 75.0448
R20198 a_n2848_n452.n92 a_n2848_n452.n39 11.2134
R20199 a_n2848_n452.n9 a_n2848_n452.n93 161.3
R20200 a_n2848_n452.n43 a_n2848_n452.n89 20.9683
R20201 a_n2848_n452.n41 a_n2848_n452.n7 75.0448
R20202 a_n2848_n452.n90 a_n2848_n452.n41 11.2134
R20203 a_n2848_n452.n7 a_n2848_n452.n91 161.3
R20204 a_n2848_n452.n79 a_n2848_n452.n5 161.3
R20205 a_n2848_n452.n81 a_n2848_n452.n80 161.3
R20206 a_n2848_n452.n49 a_n2848_n452.n50 20.9683
R20207 a_n2848_n452.n4 a_n2848_n452.n45 70.3058
R20208 a_n2848_n452.n44 a_n2848_n452.n5 70.1674
R20209 a_n2848_n452.n59 a_n2848_n452.n44 20.9683
R20210 a_n2848_n452.n5 a_n2848_n452.n60 161.3
R20211 a_n2848_n452.n2 a_n2848_n452.n47 70.1674
R20212 a_n2848_n452.n47 a_n2848_n452.n54 20.9683
R20213 a_n2848_n452.n46 a_n2848_n452.n2 75.0448
R20214 a_n2848_n452.n56 a_n2848_n452.n46 11.2134
R20215 a_n2848_n452.n0 a_n2848_n452.n3 44.8194
R20216 a_n2848_n452.n76 a_n2848_n452.n74 81.4626
R20217 a_n2848_n452.n67 a_n2848_n452.n65 81.4626
R20218 a_n2848_n452.n63 a_n2848_n452.n61 81.4626
R20219 a_n2848_n452.n76 a_n2848_n452.n75 80.9324
R20220 a_n2848_n452.n28 a_n2848_n452.n77 80.9324
R20221 a_n2848_n452.n27 a_n2848_n452.n73 80.9324
R20222 a_n2848_n452.n72 a_n2848_n452.n71 80.9324
R20223 a_n2848_n452.n70 a_n2848_n452.n69 80.9324
R20224 a_n2848_n452.n67 a_n2848_n452.n66 80.9324
R20225 a_n2848_n452.n26 a_n2848_n452.n68 80.9324
R20226 a_n2848_n452.n25 a_n2848_n452.n64 80.9324
R20227 a_n2848_n452.n63 a_n2848_n452.n62 80.9324
R20228 a_n2848_n452.n23 a_n2848_n452.t20 74.6477
R20229 a_n2848_n452.n22 a_n2848_n452.t38 74.6477
R20230 a_n2848_n452.n84 a_n2848_n452.t32 74.2899
R20231 a_n2848_n452.n24 a_n2848_n452.t28 74.2897
R20232 a_n2848_n452.n23 a_n2848_n452.n51 70.6783
R20233 a_n2848_n452.n22 a_n2848_n452.n82 70.6783
R20234 a_n2848_n452.n22 a_n2848_n452.n83 70.6783
R20235 a_n2848_n452.n106 a_n2848_n452.n24 70.6782
R20236 a_n2848_n452.n57 a_n2848_n452.n56 48.2005
R20237 a_n2848_n452.n55 a_n2848_n452.n47 20.9683
R20238 a_n2848_n452.n44 a_n2848_n452.n58 20.9683
R20239 a_n2848_n452.n78 a_n2848_n452.n49 20.9683
R20240 a_n2848_n452.n103 a_n2848_n452.n102 48.2005
R20241 a_n2848_n452.n104 a_n2848_n452.n33 20.9683
R20242 a_n2848_n452.n100 a_n2848_n452.n99 48.2005
R20243 a_n2848_n452.n101 a_n2848_n452.n30 20.9683
R20244 a_n2848_n452.n91 a_n2848_n452.n90 48.2005
R20245 a_n2848_n452.t69 a_n2848_n452.n43 533.335
R20246 a_n2848_n452.n93 a_n2848_n452.n92 48.2005
R20247 a_n2848_n452.t74 a_n2848_n452.n40 533.335
R20248 a_n2848_n452.n95 a_n2848_n452.n94 48.2005
R20249 a_n2848_n452.t63 a_n2848_n452.n38 533.335
R20250 a_n2848_n452.n97 a_n2848_n452.n96 48.2005
R20251 a_n2848_n452.t59 a_n2848_n452.n36 533.335
R20252 a_n2848_n452.n48 a_n2848_n452.t73 533.058
R20253 a_n2848_n452.n80 a_n2848_n452.n79 47.4702
R20254 a_n2848_n452.t27 a_n2848_n452.n34 533.058
R20255 a_n2848_n452.t51 a_n2848_n452.n31 533.058
R20256 a_n2848_n452.n70 a_n2848_n452.n26 33.585
R20257 a_n2848_n452.n46 a_n2848_n452.n54 35.3134
R20258 a_n2848_n452.n60 a_n2848_n452.n50 24.1005
R20259 a_n2848_n452.n60 a_n2848_n452.n59 24.1005
R20260 a_n2848_n452.n52 a_n2848_n452.n32 35.3134
R20261 a_n2848_n452.n53 a_n2848_n452.n29 35.3134
R20262 a_n2848_n452.n41 a_n2848_n452.n89 35.3134
R20263 a_n2848_n452.n39 a_n2848_n452.n88 35.3134
R20264 a_n2848_n452.n37 a_n2848_n452.n87 35.3134
R20265 a_n2848_n452.n35 a_n2848_n452.n86 35.3134
R20266 a_n2848_n452.n5 a_n2848_n452.n28 23.891
R20267 a_n2848_n452.n20 a_n2848_n452.n98 12.046
R20268 a_n2848_n452.n1 a_n2848_n452.n42 11.8414
R20269 a_n2848_n452.n85 a_n2848_n452.n81 10.5365
R20270 a_n2848_n452.n24 a_n2848_n452.n105 9.50122
R20271 a_n2848_n452.n6 a_n2848_n452.n42 7.47588
R20272 a_n2848_n452.n98 a_n2848_n452.n13 7.47588
R20273 a_n2848_n452.n105 a_n2848_n452.n14 6.70126
R20274 a_n2848_n452.n85 a_n2848_n452.n84 5.65783
R20275 a_n2848_n452.n105 a_n2848_n452.n42 5.3452
R20276 a_n2848_n452.n16 a_n2848_n452.n18 3.95126
R20277 a_n2848_n452.n4 a_n2848_n452.n0 3.95126
R20278 a_n2848_n452.n51 a_n2848_n452.t40 3.61217
R20279 a_n2848_n452.n51 a_n2848_n452.t26 3.61217
R20280 a_n2848_n452.n82 a_n2848_n452.t30 3.61217
R20281 a_n2848_n452.n82 a_n2848_n452.t22 3.61217
R20282 a_n2848_n452.n83 a_n2848_n452.t36 3.61217
R20283 a_n2848_n452.n83 a_n2848_n452.t34 3.61217
R20284 a_n2848_n452.n106 a_n2848_n452.t24 3.61217
R20285 a_n2848_n452.t18 a_n2848_n452.n106 3.61217
R20286 a_n2848_n452.n74 a_n2848_n452.t46 2.82907
R20287 a_n2848_n452.n74 a_n2848_n452.t43 2.82907
R20288 a_n2848_n452.n75 a_n2848_n452.t16 2.82907
R20289 a_n2848_n452.n75 a_n2848_n452.t13 2.82907
R20290 a_n2848_n452.n77 a_n2848_n452.t14 2.82907
R20291 a_n2848_n452.n77 a_n2848_n452.t8 2.82907
R20292 a_n2848_n452.n73 a_n2848_n452.t47 2.82907
R20293 a_n2848_n452.n73 a_n2848_n452.t11 2.82907
R20294 a_n2848_n452.n71 a_n2848_n452.t6 2.82907
R20295 a_n2848_n452.n71 a_n2848_n452.t0 2.82907
R20296 a_n2848_n452.n69 a_n2848_n452.t44 2.82907
R20297 a_n2848_n452.n69 a_n2848_n452.t10 2.82907
R20298 a_n2848_n452.n65 a_n2848_n452.t5 2.82907
R20299 a_n2848_n452.n65 a_n2848_n452.t1 2.82907
R20300 a_n2848_n452.n66 a_n2848_n452.t42 2.82907
R20301 a_n2848_n452.n66 a_n2848_n452.t7 2.82907
R20302 a_n2848_n452.n68 a_n2848_n452.t2 2.82907
R20303 a_n2848_n452.n68 a_n2848_n452.t15 2.82907
R20304 a_n2848_n452.n64 a_n2848_n452.t12 2.82907
R20305 a_n2848_n452.n64 a_n2848_n452.t41 2.82907
R20306 a_n2848_n452.n62 a_n2848_n452.t4 2.82907
R20307 a_n2848_n452.n62 a_n2848_n452.t45 2.82907
R20308 a_n2848_n452.n61 a_n2848_n452.t9 2.82907
R20309 a_n2848_n452.n61 a_n2848_n452.t3 2.82907
R20310 a_n2848_n452.n98 a_n2848_n452.n85 1.30542
R20311 a_n2848_n452.n10 a_n2848_n452.n9 1.04595
R20312 a_n2848_n452.n3 a_n2848_n452.n57 13.657
R20313 a_n2848_n452.n55 a_n2848_n452.n48 21.4216
R20314 a_n2848_n452.n58 a_n2848_n452.n45 21.4216
R20315 a_n2848_n452.n79 a_n2848_n452.n78 0.730803
R20316 a_n2848_n452.n102 a_n2848_n452.n17 13.657
R20317 a_n2848_n452.n34 a_n2848_n452.n104 21.4216
R20318 a_n2848_n452.n99 a_n2848_n452.n21 13.657
R20319 a_n2848_n452.n31 a_n2848_n452.n101 21.4216
R20320 a_n2848_n452.n20 a_n2848_n452.n19 0.758076
R20321 a_n2848_n452.n19 a_n2848_n452.n18 0.758076
R20322 a_n2848_n452.n16 a_n2848_n452.n15 0.758076
R20323 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R20324 a_n2848_n452.n13 a_n2848_n452.n12 0.758076
R20325 a_n2848_n452.n11 a_n2848_n452.n10 0.758076
R20326 a_n2848_n452.n9 a_n2848_n452.n8 0.758076
R20327 a_n2848_n452.n7 a_n2848_n452.n6 0.758076
R20328 a_n2848_n452.n5 a_n2848_n452.n4 0.758076
R20329 a_n2848_n452.n2 a_n2848_n452.n0 0.758076
R20330 a_n2848_n452.n2 a_n2848_n452.n1 0.758076
R20331 a_n2848_n452.n81 a_n2848_n452.n5 0.720197
R20332 a_n2848_n452.n24 a_n2848_n452.n23 0.716017
R20333 a_n2848_n452.n84 a_n2848_n452.n22 0.716017
R20334 a_n2848_n452.n12 a_n2848_n452.n11 0.67853
R20335 a_n2848_n452.n8 a_n2848_n452.n7 0.67853
R20336 a_n2848_n452.n25 a_n2848_n452.n63 0.530672
R20337 a_n2848_n452.n26 a_n2848_n452.n67 0.530672
R20338 a_n2848_n452.n72 a_n2848_n452.n70 0.530672
R20339 a_n2848_n452.n27 a_n2848_n452.n72 0.530672
R20340 a_n2848_n452.n28 a_n2848_n452.n76 0.530672
R20341 a_n2848_n452.n28 a_n2848_n452.n27 0.530672
R20342 a_n2848_n452.n26 a_n2848_n452.n25 0.530672
R20343 a_n1986_8322.n6 a_n1986_8322.t6 74.6477
R20344 a_n1986_8322.n1 a_n1986_8322.t13 74.6477
R20345 a_n1986_8322.t22 a_n1986_8322.n18 74.6476
R20346 a_n1986_8322.n14 a_n1986_8322.t15 74.2899
R20347 a_n1986_8322.n7 a_n1986_8322.t4 74.2899
R20348 a_n1986_8322.n8 a_n1986_8322.t7 74.2899
R20349 a_n1986_8322.n11 a_n1986_8322.t8 74.2899
R20350 a_n1986_8322.n4 a_n1986_8322.t12 74.2899
R20351 a_n1986_8322.n18 a_n1986_8322.n17 70.6783
R20352 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R20353 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R20354 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R20355 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R20356 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R20357 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R20358 a_n1986_8322.n13 a_n1986_8322.t2 9.7972
R20359 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R20360 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R20361 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R20362 a_n1986_8322.n17 a_n1986_8322.t20 3.61217
R20363 a_n1986_8322.n17 a_n1986_8322.t17 3.61217
R20364 a_n1986_8322.n15 a_n1986_8322.t14 3.61217
R20365 a_n1986_8322.n15 a_n1986_8322.t23 3.61217
R20366 a_n1986_8322.n5 a_n1986_8322.t10 3.61217
R20367 a_n1986_8322.n5 a_n1986_8322.t9 3.61217
R20368 a_n1986_8322.n9 a_n1986_8322.t5 3.61217
R20369 a_n1986_8322.n9 a_n1986_8322.t11 3.61217
R20370 a_n1986_8322.n0 a_n1986_8322.t21 3.61217
R20371 a_n1986_8322.n0 a_n1986_8322.t16 3.61217
R20372 a_n1986_8322.n2 a_n1986_8322.t19 3.61217
R20373 a_n1986_8322.n2 a_n1986_8322.t18 3.61217
R20374 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R20375 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R20376 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R20377 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R20378 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R20379 a_n1986_8322.n16 a_n1986_8322.n14 0.358259
R20380 a_n1986_8322.n18 a_n1986_8322.n16 0.358259
R20381 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R20382 a_n1986_8322.t3 a_n1986_8322.t0 0.0788333
R20383 a_n1986_8322.t1 a_n1986_8322.t3 0.0631667
R20384 a_n1986_8322.t2 a_n1986_8322.t1 0.0471944
R20385 a_n1986_8322.t2 a_n1986_8322.t0 0.0453889
R20386 a_n1808_13878.n16 a_n1808_13878.n0 98.9633
R20387 a_n1808_13878.n3 a_n1808_13878.n1 98.7517
R20388 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R20389 a_n1808_13878.n3 a_n1808_13878.n2 98.6055
R20390 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R20391 a_n1808_13878.n15 a_n1808_13878.n14 98.6054
R20392 a_n1808_13878.n7 a_n1808_13878.t1 74.6477
R20393 a_n1808_13878.n12 a_n1808_13878.t2 74.2899
R20394 a_n1808_13878.n9 a_n1808_13878.t3 74.2899
R20395 a_n1808_13878.n8 a_n1808_13878.t0 74.2899
R20396 a_n1808_13878.n11 a_n1808_13878.n10 70.6783
R20397 a_n1808_13878.n7 a_n1808_13878.n6 70.6783
R20398 a_n1808_13878.n13 a_n1808_13878.n5 13.5694
R20399 a_n1808_13878.n15 a_n1808_13878.n13 11.5762
R20400 a_n1808_13878.n13 a_n1808_13878.n12 6.2408
R20401 a_n1808_13878.n14 a_n1808_13878.t15 3.61217
R20402 a_n1808_13878.n14 a_n1808_13878.t16 3.61217
R20403 a_n1808_13878.n0 a_n1808_13878.t13 3.61217
R20404 a_n1808_13878.n0 a_n1808_13878.t17 3.61217
R20405 a_n1808_13878.n10 a_n1808_13878.t6 3.61217
R20406 a_n1808_13878.n10 a_n1808_13878.t7 3.61217
R20407 a_n1808_13878.n6 a_n1808_13878.t4 3.61217
R20408 a_n1808_13878.n6 a_n1808_13878.t5 3.61217
R20409 a_n1808_13878.n4 a_n1808_13878.t12 3.61217
R20410 a_n1808_13878.n4 a_n1808_13878.t19 3.61217
R20411 a_n1808_13878.n2 a_n1808_13878.t14 3.61217
R20412 a_n1808_13878.n2 a_n1808_13878.t9 3.61217
R20413 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R20414 a_n1808_13878.n1 a_n1808_13878.t10 3.61217
R20415 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R20416 a_n1808_13878.n17 a_n1808_13878.t11 3.61217
R20417 a_n1808_13878.n8 a_n1808_13878.n7 0.358259
R20418 a_n1808_13878.n11 a_n1808_13878.n9 0.358259
R20419 a_n1808_13878.n12 a_n1808_13878.n11 0.358259
R20420 a_n1808_13878.n16 a_n1808_13878.n15 0.358259
R20421 a_n1808_13878.n5 a_n1808_13878.n3 0.146627
R20422 a_n1808_13878.n9 a_n1808_13878.n8 0.101793
R20423 plus.n76 plus.t11 250.337
R20424 plus.n15 plus.t14 250.337
R20425 plus.n124 plus.t1 243.97
R20426 plus.n120 plus.t24 231.093
R20427 plus.n59 plus.t20 231.093
R20428 plus.n124 plus.n123 223.454
R20429 plus.n126 plus.n125 223.454
R20430 plus.n77 plus.t5 187.445
R20431 plus.n74 plus.t22 187.445
R20432 plus.n72 plus.t21 187.445
R20433 plus.n89 plus.t16 187.445
R20434 plus.n95 plus.t17 187.445
R20435 plus.n68 plus.t13 187.445
R20436 plus.n66 plus.t15 187.445
R20437 plus.n107 plus.t10 187.445
R20438 plus.n113 plus.t26 187.445
R20439 plus.n62 plus.t28 187.445
R20440 plus.n1 plus.t23 187.445
R20441 plus.n52 plus.t6 187.445
R20442 plus.n46 plus.t12 187.445
R20443 plus.n5 plus.t8 187.445
R20444 plus.n7 plus.t7 187.445
R20445 plus.n34 plus.t19 187.445
R20446 plus.n28 plus.t18 187.445
R20447 plus.n11 plus.t27 187.445
R20448 plus.n13 plus.t25 187.445
R20449 plus.n16 plus.t9 187.445
R20450 plus.n121 plus.n120 161.3
R20451 plus.n119 plus.n61 161.3
R20452 plus.n118 plus.n117 161.3
R20453 plus.n116 plus.n115 161.3
R20454 plus.n114 plus.n63 161.3
R20455 plus.n112 plus.n111 161.3
R20456 plus.n110 plus.n64 161.3
R20457 plus.n109 plus.n108 161.3
R20458 plus.n106 plus.n65 161.3
R20459 plus.n105 plus.n104 161.3
R20460 plus.n103 plus.n102 161.3
R20461 plus.n101 plus.n67 161.3
R20462 plus.n100 plus.n99 161.3
R20463 plus.n98 plus.n97 161.3
R20464 plus.n96 plus.n69 161.3
R20465 plus.n94 plus.n93 161.3
R20466 plus.n92 plus.n70 161.3
R20467 plus.n91 plus.n90 161.3
R20468 plus.n88 plus.n71 161.3
R20469 plus.n87 plus.n86 161.3
R20470 plus.n85 plus.n84 161.3
R20471 plus.n83 plus.n73 161.3
R20472 plus.n82 plus.n81 161.3
R20473 plus.n80 plus.n79 161.3
R20474 plus.n78 plus.n75 161.3
R20475 plus.n17 plus.n14 161.3
R20476 plus.n19 plus.n18 161.3
R20477 plus.n21 plus.n20 161.3
R20478 plus.n22 plus.n12 161.3
R20479 plus.n24 plus.n23 161.3
R20480 plus.n26 plus.n25 161.3
R20481 plus.n27 plus.n10 161.3
R20482 plus.n30 plus.n29 161.3
R20483 plus.n31 plus.n9 161.3
R20484 plus.n33 plus.n32 161.3
R20485 plus.n35 plus.n8 161.3
R20486 plus.n37 plus.n36 161.3
R20487 plus.n39 plus.n38 161.3
R20488 plus.n40 plus.n6 161.3
R20489 plus.n42 plus.n41 161.3
R20490 plus.n44 plus.n43 161.3
R20491 plus.n45 plus.n4 161.3
R20492 plus.n48 plus.n47 161.3
R20493 plus.n49 plus.n3 161.3
R20494 plus.n51 plus.n50 161.3
R20495 plus.n53 plus.n2 161.3
R20496 plus.n55 plus.n54 161.3
R20497 plus.n57 plus.n56 161.3
R20498 plus.n58 plus.n0 161.3
R20499 plus.n60 plus.n59 161.3
R20500 plus.n88 plus.n87 56.5617
R20501 plus.n97 plus.n96 56.5617
R20502 plus.n106 plus.n105 56.5617
R20503 plus.n45 plus.n44 56.5617
R20504 plus.n36 plus.n35 56.5617
R20505 plus.n27 plus.n26 56.5617
R20506 plus.n79 plus.n78 56.5617
R20507 plus.n115 plus.n114 56.5617
R20508 plus.n54 plus.n53 56.5617
R20509 plus.n18 plus.n17 56.5617
R20510 plus.n119 plus.n118 50.2647
R20511 plus.n58 plus.n57 50.2647
R20512 plus.n84 plus.n83 46.3896
R20513 plus.n108 plus.n64 46.3896
R20514 plus.n47 plus.n3 46.3896
R20515 plus.n23 plus.n22 46.3896
R20516 plus.n76 plus.n75 43.1929
R20517 plus.n15 plus.n14 43.1929
R20518 plus.n94 plus.n70 42.5146
R20519 plus.n101 plus.n100 42.5146
R20520 plus.n40 plus.n39 42.5146
R20521 plus.n33 plus.n9 42.5146
R20522 plus.n77 plus.n76 40.6041
R20523 plus.n16 plus.n15 40.6041
R20524 plus.n90 plus.n70 38.6395
R20525 plus.n102 plus.n101 38.6395
R20526 plus.n41 plus.n40 38.6395
R20527 plus.n29 plus.n9 38.6395
R20528 plus.n122 plus.n121 35.2031
R20529 plus.n83 plus.n82 34.7644
R20530 plus.n112 plus.n64 34.7644
R20531 plus.n51 plus.n3 34.7644
R20532 plus.n22 plus.n21 34.7644
R20533 plus.n79 plus.n74 21.8872
R20534 plus.n114 plus.n113 21.8872
R20535 plus.n53 plus.n52 21.8872
R20536 plus.n18 plus.n13 21.8872
R20537 plus.n89 plus.n88 19.9199
R20538 plus.n105 plus.n66 19.9199
R20539 plus.n44 plus.n5 19.9199
R20540 plus.n28 plus.n27 19.9199
R20541 plus.n123 plus.t2 19.8005
R20542 plus.n123 plus.t4 19.8005
R20543 plus.n125 plus.t3 19.8005
R20544 plus.n125 plus.t0 19.8005
R20545 plus.n96 plus.n95 17.9525
R20546 plus.n97 plus.n68 17.9525
R20547 plus.n36 plus.n7 17.9525
R20548 plus.n35 plus.n34 17.9525
R20549 plus.n87 plus.n72 15.9852
R20550 plus.n107 plus.n106 15.9852
R20551 plus.n46 plus.n45 15.9852
R20552 plus.n26 plus.n11 15.9852
R20553 plus plus.n127 14.4034
R20554 plus.n78 plus.n77 14.0178
R20555 plus.n115 plus.n62 14.0178
R20556 plus.n54 plus.n1 14.0178
R20557 plus.n17 plus.n16 14.0178
R20558 plus.n122 plus.n60 11.9342
R20559 plus.n118 plus.n62 10.575
R20560 plus.n57 plus.n1 10.575
R20561 plus.n120 plus.n119 9.49444
R20562 plus.n59 plus.n58 9.49444
R20563 plus.n84 plus.n72 8.60764
R20564 plus.n108 plus.n107 8.60764
R20565 plus.n47 plus.n46 8.60764
R20566 plus.n23 plus.n11 8.60764
R20567 plus.n95 plus.n94 6.6403
R20568 plus.n100 plus.n68 6.6403
R20569 plus.n39 plus.n7 6.6403
R20570 plus.n34 plus.n33 6.6403
R20571 plus.n127 plus.n126 5.40567
R20572 plus.n90 plus.n89 4.67295
R20573 plus.n102 plus.n66 4.67295
R20574 plus.n41 plus.n5 4.67295
R20575 plus.n29 plus.n28 4.67295
R20576 plus.n82 plus.n74 2.7056
R20577 plus.n113 plus.n112 2.7056
R20578 plus.n52 plus.n51 2.7056
R20579 plus.n21 plus.n13 2.7056
R20580 plus.n127 plus.n122 1.188
R20581 plus.n126 plus.n124 0.716017
R20582 plus.n80 plus.n75 0.189894
R20583 plus.n81 plus.n80 0.189894
R20584 plus.n81 plus.n73 0.189894
R20585 plus.n85 plus.n73 0.189894
R20586 plus.n86 plus.n85 0.189894
R20587 plus.n86 plus.n71 0.189894
R20588 plus.n91 plus.n71 0.189894
R20589 plus.n92 plus.n91 0.189894
R20590 plus.n93 plus.n92 0.189894
R20591 plus.n93 plus.n69 0.189894
R20592 plus.n98 plus.n69 0.189894
R20593 plus.n99 plus.n98 0.189894
R20594 plus.n99 plus.n67 0.189894
R20595 plus.n103 plus.n67 0.189894
R20596 plus.n104 plus.n103 0.189894
R20597 plus.n104 plus.n65 0.189894
R20598 plus.n109 plus.n65 0.189894
R20599 plus.n110 plus.n109 0.189894
R20600 plus.n111 plus.n110 0.189894
R20601 plus.n111 plus.n63 0.189894
R20602 plus.n116 plus.n63 0.189894
R20603 plus.n117 plus.n116 0.189894
R20604 plus.n117 plus.n61 0.189894
R20605 plus.n121 plus.n61 0.189894
R20606 plus.n60 plus.n0 0.189894
R20607 plus.n56 plus.n0 0.189894
R20608 plus.n56 plus.n55 0.189894
R20609 plus.n55 plus.n2 0.189894
R20610 plus.n50 plus.n2 0.189894
R20611 plus.n50 plus.n49 0.189894
R20612 plus.n49 plus.n48 0.189894
R20613 plus.n48 plus.n4 0.189894
R20614 plus.n43 plus.n4 0.189894
R20615 plus.n43 plus.n42 0.189894
R20616 plus.n42 plus.n6 0.189894
R20617 plus.n38 plus.n6 0.189894
R20618 plus.n38 plus.n37 0.189894
R20619 plus.n37 plus.n8 0.189894
R20620 plus.n32 plus.n8 0.189894
R20621 plus.n32 plus.n31 0.189894
R20622 plus.n31 plus.n30 0.189894
R20623 plus.n30 plus.n10 0.189894
R20624 plus.n25 plus.n10 0.189894
R20625 plus.n25 plus.n24 0.189894
R20626 plus.n24 plus.n12 0.189894
R20627 plus.n20 plus.n12 0.189894
R20628 plus.n20 plus.n19 0.189894
R20629 plus.n19 plus.n14 0.189894
R20630 a_n3106_n452.n1 a_n3106_n452.t33 214.321
R20631 a_n3106_n452.n14 a_n3106_n452.t54 214.321
R20632 a_n3106_n452.n15 a_n3106_n452.t52 214.321
R20633 a_n3106_n452.n16 a_n3106_n452.t40 214.321
R20634 a_n3106_n452.n17 a_n3106_n452.t41 214.321
R20635 a_n3106_n452.n18 a_n3106_n452.t55 214.321
R20636 a_n3106_n452.n19 a_n3106_n452.t0 214.321
R20637 a_n3106_n452.n20 a_n3106_n452.t53 214.321
R20638 a_n3106_n452.n0 a_n3106_n452.t19 55.8337
R20639 a_n3106_n452.n2 a_n3106_n452.t47 55.8337
R20640 a_n3106_n452.n13 a_n3106_n452.t48 55.8337
R20641 a_n3106_n452.n47 a_n3106_n452.t6 55.8335
R20642 a_n3106_n452.n45 a_n3106_n452.t26 55.8335
R20643 a_n3106_n452.n34 a_n3106_n452.t35 55.8335
R20644 a_n3106_n452.n33 a_n3106_n452.t16 55.8335
R20645 a_n3106_n452.n22 a_n3106_n452.t10 55.8335
R20646 a_n3106_n452.n49 a_n3106_n452.n48 53.0052
R20647 a_n3106_n452.n51 a_n3106_n452.n50 53.0052
R20648 a_n3106_n452.n53 a_n3106_n452.n52 53.0052
R20649 a_n3106_n452.n55 a_n3106_n452.n54 53.0052
R20650 a_n3106_n452.n4 a_n3106_n452.n3 53.0052
R20651 a_n3106_n452.n6 a_n3106_n452.n5 53.0052
R20652 a_n3106_n452.n8 a_n3106_n452.n7 53.0052
R20653 a_n3106_n452.n10 a_n3106_n452.n9 53.0052
R20654 a_n3106_n452.n12 a_n3106_n452.n11 53.0052
R20655 a_n3106_n452.n44 a_n3106_n452.n43 53.0051
R20656 a_n3106_n452.n42 a_n3106_n452.n41 53.0051
R20657 a_n3106_n452.n40 a_n3106_n452.n39 53.0051
R20658 a_n3106_n452.n38 a_n3106_n452.n37 53.0051
R20659 a_n3106_n452.n36 a_n3106_n452.n35 53.0051
R20660 a_n3106_n452.n32 a_n3106_n452.n31 53.0051
R20661 a_n3106_n452.n30 a_n3106_n452.n29 53.0051
R20662 a_n3106_n452.n28 a_n3106_n452.n27 53.0051
R20663 a_n3106_n452.n26 a_n3106_n452.n25 53.0051
R20664 a_n3106_n452.n24 a_n3106_n452.n23 53.0051
R20665 a_n3106_n452.n57 a_n3106_n452.n56 53.0051
R20666 a_n3106_n452.n21 a_n3106_n452.n13 12.2417
R20667 a_n3106_n452.n47 a_n3106_n452.n46 12.2417
R20668 a_n3106_n452.n22 a_n3106_n452.n21 5.16214
R20669 a_n3106_n452.n46 a_n3106_n452.n45 5.16214
R20670 a_n3106_n452.n48 a_n3106_n452.t4 2.82907
R20671 a_n3106_n452.n48 a_n3106_n452.t2 2.82907
R20672 a_n3106_n452.n50 a_n3106_n452.t15 2.82907
R20673 a_n3106_n452.n50 a_n3106_n452.t20 2.82907
R20674 a_n3106_n452.n52 a_n3106_n452.t13 2.82907
R20675 a_n3106_n452.n52 a_n3106_n452.t17 2.82907
R20676 a_n3106_n452.n54 a_n3106_n452.t9 2.82907
R20677 a_n3106_n452.n54 a_n3106_n452.t14 2.82907
R20678 a_n3106_n452.n3 a_n3106_n452.t39 2.82907
R20679 a_n3106_n452.n3 a_n3106_n452.t50 2.82907
R20680 a_n3106_n452.n5 a_n3106_n452.t34 2.82907
R20681 a_n3106_n452.n5 a_n3106_n452.t44 2.82907
R20682 a_n3106_n452.n7 a_n3106_n452.t37 2.82907
R20683 a_n3106_n452.n7 a_n3106_n452.t42 2.82907
R20684 a_n3106_n452.n9 a_n3106_n452.t1 2.82907
R20685 a_n3106_n452.n9 a_n3106_n452.t51 2.82907
R20686 a_n3106_n452.n11 a_n3106_n452.t36 2.82907
R20687 a_n3106_n452.n11 a_n3106_n452.t31 2.82907
R20688 a_n3106_n452.n43 a_n3106_n452.t32 2.82907
R20689 a_n3106_n452.n43 a_n3106_n452.t30 2.82907
R20690 a_n3106_n452.n41 a_n3106_n452.t43 2.82907
R20691 a_n3106_n452.n41 a_n3106_n452.t46 2.82907
R20692 a_n3106_n452.n39 a_n3106_n452.t45 2.82907
R20693 a_n3106_n452.n39 a_n3106_n452.t27 2.82907
R20694 a_n3106_n452.n37 a_n3106_n452.t49 2.82907
R20695 a_n3106_n452.n37 a_n3106_n452.t38 2.82907
R20696 a_n3106_n452.n35 a_n3106_n452.t28 2.82907
R20697 a_n3106_n452.n35 a_n3106_n452.t29 2.82907
R20698 a_n3106_n452.n31 a_n3106_n452.t5 2.82907
R20699 a_n3106_n452.n31 a_n3106_n452.t21 2.82907
R20700 a_n3106_n452.n29 a_n3106_n452.t12 2.82907
R20701 a_n3106_n452.n29 a_n3106_n452.t3 2.82907
R20702 a_n3106_n452.n27 a_n3106_n452.t23 2.82907
R20703 a_n3106_n452.n27 a_n3106_n452.t11 2.82907
R20704 a_n3106_n452.n25 a_n3106_n452.t18 2.82907
R20705 a_n3106_n452.n25 a_n3106_n452.t22 2.82907
R20706 a_n3106_n452.n23 a_n3106_n452.t7 2.82907
R20707 a_n3106_n452.n23 a_n3106_n452.t24 2.82907
R20708 a_n3106_n452.t25 a_n3106_n452.n57 2.82907
R20709 a_n3106_n452.n57 a_n3106_n452.t8 2.82907
R20710 a_n3106_n452.n46 a_n3106_n452.n1 2.54197
R20711 a_n3106_n452.n21 a_n3106_n452.n20 2.0129
R20712 a_n3106_n452.n20 a_n3106_n452.n19 0.672012
R20713 a_n3106_n452.n19 a_n3106_n452.n18 0.672012
R20714 a_n3106_n452.n18 a_n3106_n452.n17 0.672012
R20715 a_n3106_n452.n17 a_n3106_n452.n16 0.672012
R20716 a_n3106_n452.n16 a_n3106_n452.n15 0.672012
R20717 a_n3106_n452.n15 a_n3106_n452.n14 0.672012
R20718 a_n3106_n452.n14 a_n3106_n452.n1 0.672012
R20719 a_n3106_n452.n24 a_n3106_n452.n22 0.530672
R20720 a_n3106_n452.n26 a_n3106_n452.n24 0.530672
R20721 a_n3106_n452.n28 a_n3106_n452.n26 0.530672
R20722 a_n3106_n452.n30 a_n3106_n452.n28 0.530672
R20723 a_n3106_n452.n32 a_n3106_n452.n30 0.530672
R20724 a_n3106_n452.n33 a_n3106_n452.n32 0.530672
R20725 a_n3106_n452.n36 a_n3106_n452.n34 0.530672
R20726 a_n3106_n452.n38 a_n3106_n452.n36 0.530672
R20727 a_n3106_n452.n40 a_n3106_n452.n38 0.530672
R20728 a_n3106_n452.n42 a_n3106_n452.n40 0.530672
R20729 a_n3106_n452.n44 a_n3106_n452.n42 0.530672
R20730 a_n3106_n452.n45 a_n3106_n452.n44 0.530672
R20731 a_n3106_n452.n13 a_n3106_n452.n12 0.530672
R20732 a_n3106_n452.n12 a_n3106_n452.n10 0.530672
R20733 a_n3106_n452.n10 a_n3106_n452.n8 0.530672
R20734 a_n3106_n452.n8 a_n3106_n452.n6 0.530672
R20735 a_n3106_n452.n6 a_n3106_n452.n4 0.530672
R20736 a_n3106_n452.n4 a_n3106_n452.n2 0.530672
R20737 a_n3106_n452.n56 a_n3106_n452.n0 0.530672
R20738 a_n3106_n452.n56 a_n3106_n452.n55 0.530672
R20739 a_n3106_n452.n55 a_n3106_n452.n53 0.530672
R20740 a_n3106_n452.n53 a_n3106_n452.n51 0.530672
R20741 a_n3106_n452.n51 a_n3106_n452.n49 0.530672
R20742 a_n3106_n452.n49 a_n3106_n452.n47 0.530672
R20743 a_n3106_n452.n34 a_n3106_n452.n33 0.235414
R20744 a_n3106_n452.n2 a_n3106_n452.n0 0.235414
R20745 outputibias.n27 outputibias.n1 289.615
R20746 outputibias.n58 outputibias.n32 289.615
R20747 outputibias.n90 outputibias.n64 289.615
R20748 outputibias.n122 outputibias.n96 289.615
R20749 outputibias.n28 outputibias.n27 185
R20750 outputibias.n26 outputibias.n25 185
R20751 outputibias.n5 outputibias.n4 185
R20752 outputibias.n20 outputibias.n19 185
R20753 outputibias.n18 outputibias.n17 185
R20754 outputibias.n9 outputibias.n8 185
R20755 outputibias.n12 outputibias.n11 185
R20756 outputibias.n59 outputibias.n58 185
R20757 outputibias.n57 outputibias.n56 185
R20758 outputibias.n36 outputibias.n35 185
R20759 outputibias.n51 outputibias.n50 185
R20760 outputibias.n49 outputibias.n48 185
R20761 outputibias.n40 outputibias.n39 185
R20762 outputibias.n43 outputibias.n42 185
R20763 outputibias.n91 outputibias.n90 185
R20764 outputibias.n89 outputibias.n88 185
R20765 outputibias.n68 outputibias.n67 185
R20766 outputibias.n83 outputibias.n82 185
R20767 outputibias.n81 outputibias.n80 185
R20768 outputibias.n72 outputibias.n71 185
R20769 outputibias.n75 outputibias.n74 185
R20770 outputibias.n123 outputibias.n122 185
R20771 outputibias.n121 outputibias.n120 185
R20772 outputibias.n100 outputibias.n99 185
R20773 outputibias.n115 outputibias.n114 185
R20774 outputibias.n113 outputibias.n112 185
R20775 outputibias.n104 outputibias.n103 185
R20776 outputibias.n107 outputibias.n106 185
R20777 outputibias.n0 outputibias.t9 178.945
R20778 outputibias.n133 outputibias.t8 177.018
R20779 outputibias.n132 outputibias.t11 177.018
R20780 outputibias.n0 outputibias.t10 177.018
R20781 outputibias.t5 outputibias.n10 147.661
R20782 outputibias.t7 outputibias.n41 147.661
R20783 outputibias.t1 outputibias.n73 147.661
R20784 outputibias.t3 outputibias.n105 147.661
R20785 outputibias.n128 outputibias.t4 132.363
R20786 outputibias.n128 outputibias.t6 130.436
R20787 outputibias.n129 outputibias.t0 130.436
R20788 outputibias.n130 outputibias.t2 130.436
R20789 outputibias.n27 outputibias.n26 104.615
R20790 outputibias.n26 outputibias.n4 104.615
R20791 outputibias.n19 outputibias.n4 104.615
R20792 outputibias.n19 outputibias.n18 104.615
R20793 outputibias.n18 outputibias.n8 104.615
R20794 outputibias.n11 outputibias.n8 104.615
R20795 outputibias.n58 outputibias.n57 104.615
R20796 outputibias.n57 outputibias.n35 104.615
R20797 outputibias.n50 outputibias.n35 104.615
R20798 outputibias.n50 outputibias.n49 104.615
R20799 outputibias.n49 outputibias.n39 104.615
R20800 outputibias.n42 outputibias.n39 104.615
R20801 outputibias.n90 outputibias.n89 104.615
R20802 outputibias.n89 outputibias.n67 104.615
R20803 outputibias.n82 outputibias.n67 104.615
R20804 outputibias.n82 outputibias.n81 104.615
R20805 outputibias.n81 outputibias.n71 104.615
R20806 outputibias.n74 outputibias.n71 104.615
R20807 outputibias.n122 outputibias.n121 104.615
R20808 outputibias.n121 outputibias.n99 104.615
R20809 outputibias.n114 outputibias.n99 104.615
R20810 outputibias.n114 outputibias.n113 104.615
R20811 outputibias.n113 outputibias.n103 104.615
R20812 outputibias.n106 outputibias.n103 104.615
R20813 outputibias.n63 outputibias.n31 95.6354
R20814 outputibias.n63 outputibias.n62 94.6732
R20815 outputibias.n95 outputibias.n94 94.6732
R20816 outputibias.n127 outputibias.n126 94.6732
R20817 outputibias.n11 outputibias.t5 52.3082
R20818 outputibias.n42 outputibias.t7 52.3082
R20819 outputibias.n74 outputibias.t1 52.3082
R20820 outputibias.n106 outputibias.t3 52.3082
R20821 outputibias.n12 outputibias.n10 15.6674
R20822 outputibias.n43 outputibias.n41 15.6674
R20823 outputibias.n75 outputibias.n73 15.6674
R20824 outputibias.n107 outputibias.n105 15.6674
R20825 outputibias.n13 outputibias.n9 12.8005
R20826 outputibias.n44 outputibias.n40 12.8005
R20827 outputibias.n76 outputibias.n72 12.8005
R20828 outputibias.n108 outputibias.n104 12.8005
R20829 outputibias.n17 outputibias.n16 12.0247
R20830 outputibias.n48 outputibias.n47 12.0247
R20831 outputibias.n80 outputibias.n79 12.0247
R20832 outputibias.n112 outputibias.n111 12.0247
R20833 outputibias.n20 outputibias.n7 11.249
R20834 outputibias.n51 outputibias.n38 11.249
R20835 outputibias.n83 outputibias.n70 11.249
R20836 outputibias.n115 outputibias.n102 11.249
R20837 outputibias.n21 outputibias.n5 10.4732
R20838 outputibias.n52 outputibias.n36 10.4732
R20839 outputibias.n84 outputibias.n68 10.4732
R20840 outputibias.n116 outputibias.n100 10.4732
R20841 outputibias.n25 outputibias.n24 9.69747
R20842 outputibias.n56 outputibias.n55 9.69747
R20843 outputibias.n88 outputibias.n87 9.69747
R20844 outputibias.n120 outputibias.n119 9.69747
R20845 outputibias.n31 outputibias.n30 9.45567
R20846 outputibias.n62 outputibias.n61 9.45567
R20847 outputibias.n94 outputibias.n93 9.45567
R20848 outputibias.n126 outputibias.n125 9.45567
R20849 outputibias.n30 outputibias.n29 9.3005
R20850 outputibias.n3 outputibias.n2 9.3005
R20851 outputibias.n24 outputibias.n23 9.3005
R20852 outputibias.n22 outputibias.n21 9.3005
R20853 outputibias.n7 outputibias.n6 9.3005
R20854 outputibias.n16 outputibias.n15 9.3005
R20855 outputibias.n14 outputibias.n13 9.3005
R20856 outputibias.n61 outputibias.n60 9.3005
R20857 outputibias.n34 outputibias.n33 9.3005
R20858 outputibias.n55 outputibias.n54 9.3005
R20859 outputibias.n53 outputibias.n52 9.3005
R20860 outputibias.n38 outputibias.n37 9.3005
R20861 outputibias.n47 outputibias.n46 9.3005
R20862 outputibias.n45 outputibias.n44 9.3005
R20863 outputibias.n93 outputibias.n92 9.3005
R20864 outputibias.n66 outputibias.n65 9.3005
R20865 outputibias.n87 outputibias.n86 9.3005
R20866 outputibias.n85 outputibias.n84 9.3005
R20867 outputibias.n70 outputibias.n69 9.3005
R20868 outputibias.n79 outputibias.n78 9.3005
R20869 outputibias.n77 outputibias.n76 9.3005
R20870 outputibias.n125 outputibias.n124 9.3005
R20871 outputibias.n98 outputibias.n97 9.3005
R20872 outputibias.n119 outputibias.n118 9.3005
R20873 outputibias.n117 outputibias.n116 9.3005
R20874 outputibias.n102 outputibias.n101 9.3005
R20875 outputibias.n111 outputibias.n110 9.3005
R20876 outputibias.n109 outputibias.n108 9.3005
R20877 outputibias.n28 outputibias.n3 8.92171
R20878 outputibias.n59 outputibias.n34 8.92171
R20879 outputibias.n91 outputibias.n66 8.92171
R20880 outputibias.n123 outputibias.n98 8.92171
R20881 outputibias.n29 outputibias.n1 8.14595
R20882 outputibias.n60 outputibias.n32 8.14595
R20883 outputibias.n92 outputibias.n64 8.14595
R20884 outputibias.n124 outputibias.n96 8.14595
R20885 outputibias.n31 outputibias.n1 5.81868
R20886 outputibias.n62 outputibias.n32 5.81868
R20887 outputibias.n94 outputibias.n64 5.81868
R20888 outputibias.n126 outputibias.n96 5.81868
R20889 outputibias.n131 outputibias.n130 5.20947
R20890 outputibias.n29 outputibias.n28 5.04292
R20891 outputibias.n60 outputibias.n59 5.04292
R20892 outputibias.n92 outputibias.n91 5.04292
R20893 outputibias.n124 outputibias.n123 5.04292
R20894 outputibias.n131 outputibias.n127 4.42209
R20895 outputibias.n14 outputibias.n10 4.38594
R20896 outputibias.n45 outputibias.n41 4.38594
R20897 outputibias.n77 outputibias.n73 4.38594
R20898 outputibias.n109 outputibias.n105 4.38594
R20899 outputibias.n132 outputibias.n131 4.28454
R20900 outputibias.n25 outputibias.n3 4.26717
R20901 outputibias.n56 outputibias.n34 4.26717
R20902 outputibias.n88 outputibias.n66 4.26717
R20903 outputibias.n120 outputibias.n98 4.26717
R20904 outputibias.n24 outputibias.n5 3.49141
R20905 outputibias.n55 outputibias.n36 3.49141
R20906 outputibias.n87 outputibias.n68 3.49141
R20907 outputibias.n119 outputibias.n100 3.49141
R20908 outputibias.n21 outputibias.n20 2.71565
R20909 outputibias.n52 outputibias.n51 2.71565
R20910 outputibias.n84 outputibias.n83 2.71565
R20911 outputibias.n116 outputibias.n115 2.71565
R20912 outputibias.n17 outputibias.n7 1.93989
R20913 outputibias.n48 outputibias.n38 1.93989
R20914 outputibias.n80 outputibias.n70 1.93989
R20915 outputibias.n112 outputibias.n102 1.93989
R20916 outputibias.n130 outputibias.n129 1.9266
R20917 outputibias.n129 outputibias.n128 1.9266
R20918 outputibias.n133 outputibias.n132 1.92658
R20919 outputibias.n134 outputibias.n133 1.29913
R20920 outputibias.n16 outputibias.n9 1.16414
R20921 outputibias.n47 outputibias.n40 1.16414
R20922 outputibias.n79 outputibias.n72 1.16414
R20923 outputibias.n111 outputibias.n104 1.16414
R20924 outputibias.n127 outputibias.n95 0.962709
R20925 outputibias.n95 outputibias.n63 0.962709
R20926 outputibias.n13 outputibias.n12 0.388379
R20927 outputibias.n44 outputibias.n43 0.388379
R20928 outputibias.n76 outputibias.n75 0.388379
R20929 outputibias.n108 outputibias.n107 0.388379
R20930 outputibias.n134 outputibias.n0 0.337251
R20931 outputibias outputibias.n134 0.302375
R20932 outputibias.n30 outputibias.n2 0.155672
R20933 outputibias.n23 outputibias.n2 0.155672
R20934 outputibias.n23 outputibias.n22 0.155672
R20935 outputibias.n22 outputibias.n6 0.155672
R20936 outputibias.n15 outputibias.n6 0.155672
R20937 outputibias.n15 outputibias.n14 0.155672
R20938 outputibias.n61 outputibias.n33 0.155672
R20939 outputibias.n54 outputibias.n33 0.155672
R20940 outputibias.n54 outputibias.n53 0.155672
R20941 outputibias.n53 outputibias.n37 0.155672
R20942 outputibias.n46 outputibias.n37 0.155672
R20943 outputibias.n46 outputibias.n45 0.155672
R20944 outputibias.n93 outputibias.n65 0.155672
R20945 outputibias.n86 outputibias.n65 0.155672
R20946 outputibias.n86 outputibias.n85 0.155672
R20947 outputibias.n85 outputibias.n69 0.155672
R20948 outputibias.n78 outputibias.n69 0.155672
R20949 outputibias.n78 outputibias.n77 0.155672
R20950 outputibias.n125 outputibias.n97 0.155672
R20951 outputibias.n118 outputibias.n97 0.155672
R20952 outputibias.n118 outputibias.n117 0.155672
R20953 outputibias.n117 outputibias.n101 0.155672
R20954 outputibias.n110 outputibias.n101 0.155672
R20955 outputibias.n110 outputibias.n109 0.155672
R20956 output.n41 output.n15 289.615
R20957 output.n72 output.n46 289.615
R20958 output.n104 output.n78 289.615
R20959 output.n136 output.n110 289.615
R20960 output.n77 output.n45 197.26
R20961 output.n77 output.n76 196.298
R20962 output.n109 output.n108 196.298
R20963 output.n141 output.n140 196.298
R20964 output.n42 output.n41 185
R20965 output.n40 output.n39 185
R20966 output.n19 output.n18 185
R20967 output.n34 output.n33 185
R20968 output.n32 output.n31 185
R20969 output.n23 output.n22 185
R20970 output.n26 output.n25 185
R20971 output.n73 output.n72 185
R20972 output.n71 output.n70 185
R20973 output.n50 output.n49 185
R20974 output.n65 output.n64 185
R20975 output.n63 output.n62 185
R20976 output.n54 output.n53 185
R20977 output.n57 output.n56 185
R20978 output.n105 output.n104 185
R20979 output.n103 output.n102 185
R20980 output.n82 output.n81 185
R20981 output.n97 output.n96 185
R20982 output.n95 output.n94 185
R20983 output.n86 output.n85 185
R20984 output.n89 output.n88 185
R20985 output.n137 output.n136 185
R20986 output.n135 output.n134 185
R20987 output.n114 output.n113 185
R20988 output.n129 output.n128 185
R20989 output.n127 output.n126 185
R20990 output.n118 output.n117 185
R20991 output.n121 output.n120 185
R20992 output.t2 output.n24 147.661
R20993 output.t1 output.n55 147.661
R20994 output.t3 output.n87 147.661
R20995 output.t0 output.n119 147.661
R20996 output.n41 output.n40 104.615
R20997 output.n40 output.n18 104.615
R20998 output.n33 output.n18 104.615
R20999 output.n33 output.n32 104.615
R21000 output.n32 output.n22 104.615
R21001 output.n25 output.n22 104.615
R21002 output.n72 output.n71 104.615
R21003 output.n71 output.n49 104.615
R21004 output.n64 output.n49 104.615
R21005 output.n64 output.n63 104.615
R21006 output.n63 output.n53 104.615
R21007 output.n56 output.n53 104.615
R21008 output.n104 output.n103 104.615
R21009 output.n103 output.n81 104.615
R21010 output.n96 output.n81 104.615
R21011 output.n96 output.n95 104.615
R21012 output.n95 output.n85 104.615
R21013 output.n88 output.n85 104.615
R21014 output.n136 output.n135 104.615
R21015 output.n135 output.n113 104.615
R21016 output.n128 output.n113 104.615
R21017 output.n128 output.n127 104.615
R21018 output.n127 output.n117 104.615
R21019 output.n120 output.n117 104.615
R21020 output.n1 output.t9 77.056
R21021 output.n14 output.t10 76.6694
R21022 output.n1 output.n0 72.7095
R21023 output.n3 output.n2 72.7095
R21024 output.n5 output.n4 72.7095
R21025 output.n7 output.n6 72.7095
R21026 output.n9 output.n8 72.7095
R21027 output.n11 output.n10 72.7095
R21028 output.n13 output.n12 72.7095
R21029 output.n25 output.t2 52.3082
R21030 output.n56 output.t1 52.3082
R21031 output.n88 output.t3 52.3082
R21032 output.n120 output.t0 52.3082
R21033 output.n26 output.n24 15.6674
R21034 output.n57 output.n55 15.6674
R21035 output.n89 output.n87 15.6674
R21036 output.n121 output.n119 15.6674
R21037 output.n27 output.n23 12.8005
R21038 output.n58 output.n54 12.8005
R21039 output.n90 output.n86 12.8005
R21040 output.n122 output.n118 12.8005
R21041 output.n31 output.n30 12.0247
R21042 output.n62 output.n61 12.0247
R21043 output.n94 output.n93 12.0247
R21044 output.n126 output.n125 12.0247
R21045 output.n34 output.n21 11.249
R21046 output.n65 output.n52 11.249
R21047 output.n97 output.n84 11.249
R21048 output.n129 output.n116 11.249
R21049 output.n35 output.n19 10.4732
R21050 output.n66 output.n50 10.4732
R21051 output.n98 output.n82 10.4732
R21052 output.n130 output.n114 10.4732
R21053 output.n39 output.n38 9.69747
R21054 output.n70 output.n69 9.69747
R21055 output.n102 output.n101 9.69747
R21056 output.n134 output.n133 9.69747
R21057 output.n45 output.n44 9.45567
R21058 output.n76 output.n75 9.45567
R21059 output.n108 output.n107 9.45567
R21060 output.n140 output.n139 9.45567
R21061 output.n44 output.n43 9.3005
R21062 output.n17 output.n16 9.3005
R21063 output.n38 output.n37 9.3005
R21064 output.n36 output.n35 9.3005
R21065 output.n21 output.n20 9.3005
R21066 output.n30 output.n29 9.3005
R21067 output.n28 output.n27 9.3005
R21068 output.n75 output.n74 9.3005
R21069 output.n48 output.n47 9.3005
R21070 output.n69 output.n68 9.3005
R21071 output.n67 output.n66 9.3005
R21072 output.n52 output.n51 9.3005
R21073 output.n61 output.n60 9.3005
R21074 output.n59 output.n58 9.3005
R21075 output.n107 output.n106 9.3005
R21076 output.n80 output.n79 9.3005
R21077 output.n101 output.n100 9.3005
R21078 output.n99 output.n98 9.3005
R21079 output.n84 output.n83 9.3005
R21080 output.n93 output.n92 9.3005
R21081 output.n91 output.n90 9.3005
R21082 output.n139 output.n138 9.3005
R21083 output.n112 output.n111 9.3005
R21084 output.n133 output.n132 9.3005
R21085 output.n131 output.n130 9.3005
R21086 output.n116 output.n115 9.3005
R21087 output.n125 output.n124 9.3005
R21088 output.n123 output.n122 9.3005
R21089 output.n42 output.n17 8.92171
R21090 output.n73 output.n48 8.92171
R21091 output.n105 output.n80 8.92171
R21092 output.n137 output.n112 8.92171
R21093 output output.n141 8.15037
R21094 output.n43 output.n15 8.14595
R21095 output.n74 output.n46 8.14595
R21096 output.n106 output.n78 8.14595
R21097 output.n138 output.n110 8.14595
R21098 output.n45 output.n15 5.81868
R21099 output.n76 output.n46 5.81868
R21100 output.n108 output.n78 5.81868
R21101 output.n140 output.n110 5.81868
R21102 output.n43 output.n42 5.04292
R21103 output.n74 output.n73 5.04292
R21104 output.n106 output.n105 5.04292
R21105 output.n138 output.n137 5.04292
R21106 output.n28 output.n24 4.38594
R21107 output.n59 output.n55 4.38594
R21108 output.n91 output.n87 4.38594
R21109 output.n123 output.n119 4.38594
R21110 output.n39 output.n17 4.26717
R21111 output.n70 output.n48 4.26717
R21112 output.n102 output.n80 4.26717
R21113 output.n134 output.n112 4.26717
R21114 output.n0 output.t15 3.9605
R21115 output.n0 output.t19 3.9605
R21116 output.n2 output.t7 3.9605
R21117 output.n2 output.t11 3.9605
R21118 output.n4 output.t12 3.9605
R21119 output.n4 output.t17 3.9605
R21120 output.n6 output.t5 3.9605
R21121 output.n6 output.t13 3.9605
R21122 output.n8 output.t16 3.9605
R21123 output.n8 output.t14 3.9605
R21124 output.n10 output.t4 3.9605
R21125 output.n10 output.t6 3.9605
R21126 output.n12 output.t8 3.9605
R21127 output.n12 output.t18 3.9605
R21128 output.n38 output.n19 3.49141
R21129 output.n69 output.n50 3.49141
R21130 output.n101 output.n82 3.49141
R21131 output.n133 output.n114 3.49141
R21132 output.n35 output.n34 2.71565
R21133 output.n66 output.n65 2.71565
R21134 output.n98 output.n97 2.71565
R21135 output.n130 output.n129 2.71565
R21136 output.n31 output.n21 1.93989
R21137 output.n62 output.n52 1.93989
R21138 output.n94 output.n84 1.93989
R21139 output.n126 output.n116 1.93989
R21140 output.n30 output.n23 1.16414
R21141 output.n61 output.n54 1.16414
R21142 output.n93 output.n86 1.16414
R21143 output.n125 output.n118 1.16414
R21144 output.n141 output.n109 0.962709
R21145 output.n109 output.n77 0.962709
R21146 output.n27 output.n26 0.388379
R21147 output.n58 output.n57 0.388379
R21148 output.n90 output.n89 0.388379
R21149 output.n122 output.n121 0.388379
R21150 output.n14 output.n13 0.387128
R21151 output.n13 output.n11 0.387128
R21152 output.n11 output.n9 0.387128
R21153 output.n9 output.n7 0.387128
R21154 output.n7 output.n5 0.387128
R21155 output.n5 output.n3 0.387128
R21156 output.n3 output.n1 0.387128
R21157 output.n44 output.n16 0.155672
R21158 output.n37 output.n16 0.155672
R21159 output.n37 output.n36 0.155672
R21160 output.n36 output.n20 0.155672
R21161 output.n29 output.n20 0.155672
R21162 output.n29 output.n28 0.155672
R21163 output.n75 output.n47 0.155672
R21164 output.n68 output.n47 0.155672
R21165 output.n68 output.n67 0.155672
R21166 output.n67 output.n51 0.155672
R21167 output.n60 output.n51 0.155672
R21168 output.n60 output.n59 0.155672
R21169 output.n107 output.n79 0.155672
R21170 output.n100 output.n79 0.155672
R21171 output.n100 output.n99 0.155672
R21172 output.n99 output.n83 0.155672
R21173 output.n92 output.n83 0.155672
R21174 output.n92 output.n91 0.155672
R21175 output.n139 output.n111 0.155672
R21176 output.n132 output.n111 0.155672
R21177 output.n132 output.n131 0.155672
R21178 output.n131 output.n115 0.155672
R21179 output.n124 output.n115 0.155672
R21180 output.n124 output.n123 0.155672
R21181 output output.n14 0.126227
R21182 minus.n76 minus.t28 250.337
R21183 minus.n15 minus.t20 250.337
R21184 minus.n126 minus.t1 243.255
R21185 minus.n120 minus.t8 231.093
R21186 minus.n59 minus.t10 231.093
R21187 minus.n125 minus.n123 224.169
R21188 minus.n125 minus.n124 223.454
R21189 minus.n62 minus.t12 187.445
R21190 minus.n113 minus.t18 187.445
R21191 minus.n107 minus.t25 187.445
R21192 minus.n66 minus.t22 187.445
R21193 minus.n68 minus.t19 187.445
R21194 minus.n95 minus.t7 187.445
R21195 minus.n89 minus.t6 187.445
R21196 minus.n72 minus.t16 187.445
R21197 minus.n74 minus.t15 187.445
R21198 minus.n77 minus.t23 187.445
R21199 minus.n16 minus.t14 187.445
R21200 minus.n13 minus.t9 187.445
R21201 minus.n11 minus.t5 187.445
R21202 minus.n28 minus.t26 187.445
R21203 minus.n34 minus.t27 187.445
R21204 minus.n7 minus.t21 187.445
R21205 minus.n5 minus.t24 187.445
R21206 minus.n46 minus.t17 187.445
R21207 minus.n52 minus.t11 187.445
R21208 minus.n1 minus.t13 187.445
R21209 minus.n78 minus.n75 161.3
R21210 minus.n80 minus.n79 161.3
R21211 minus.n82 minus.n81 161.3
R21212 minus.n83 minus.n73 161.3
R21213 minus.n85 minus.n84 161.3
R21214 minus.n87 minus.n86 161.3
R21215 minus.n88 minus.n71 161.3
R21216 minus.n91 minus.n90 161.3
R21217 minus.n92 minus.n70 161.3
R21218 minus.n94 minus.n93 161.3
R21219 minus.n96 minus.n69 161.3
R21220 minus.n98 minus.n97 161.3
R21221 minus.n100 minus.n99 161.3
R21222 minus.n101 minus.n67 161.3
R21223 minus.n103 minus.n102 161.3
R21224 minus.n105 minus.n104 161.3
R21225 minus.n106 minus.n65 161.3
R21226 minus.n109 minus.n108 161.3
R21227 minus.n110 minus.n64 161.3
R21228 minus.n112 minus.n111 161.3
R21229 minus.n114 minus.n63 161.3
R21230 minus.n116 minus.n115 161.3
R21231 minus.n118 minus.n117 161.3
R21232 minus.n119 minus.n61 161.3
R21233 minus.n121 minus.n120 161.3
R21234 minus.n60 minus.n59 161.3
R21235 minus.n58 minus.n0 161.3
R21236 minus.n57 minus.n56 161.3
R21237 minus.n55 minus.n54 161.3
R21238 minus.n53 minus.n2 161.3
R21239 minus.n51 minus.n50 161.3
R21240 minus.n49 minus.n3 161.3
R21241 minus.n48 minus.n47 161.3
R21242 minus.n45 minus.n4 161.3
R21243 minus.n44 minus.n43 161.3
R21244 minus.n42 minus.n41 161.3
R21245 minus.n40 minus.n6 161.3
R21246 minus.n39 minus.n38 161.3
R21247 minus.n37 minus.n36 161.3
R21248 minus.n35 minus.n8 161.3
R21249 minus.n33 minus.n32 161.3
R21250 minus.n31 minus.n9 161.3
R21251 minus.n30 minus.n29 161.3
R21252 minus.n27 minus.n10 161.3
R21253 minus.n26 minus.n25 161.3
R21254 minus.n24 minus.n23 161.3
R21255 minus.n22 minus.n12 161.3
R21256 minus.n21 minus.n20 161.3
R21257 minus.n19 minus.n18 161.3
R21258 minus.n17 minus.n14 161.3
R21259 minus.n106 minus.n105 56.5617
R21260 minus.n97 minus.n96 56.5617
R21261 minus.n88 minus.n87 56.5617
R21262 minus.n27 minus.n26 56.5617
R21263 minus.n36 minus.n35 56.5617
R21264 minus.n45 minus.n44 56.5617
R21265 minus.n115 minus.n114 56.5617
R21266 minus.n79 minus.n78 56.5617
R21267 minus.n18 minus.n17 56.5617
R21268 minus.n54 minus.n53 56.5617
R21269 minus.n119 minus.n118 50.2647
R21270 minus.n58 minus.n57 50.2647
R21271 minus.n108 minus.n64 46.3896
R21272 minus.n84 minus.n83 46.3896
R21273 minus.n23 minus.n22 46.3896
R21274 minus.n47 minus.n3 46.3896
R21275 minus.n76 minus.n75 43.1929
R21276 minus.n15 minus.n14 43.1929
R21277 minus.n101 minus.n100 42.5146
R21278 minus.n94 minus.n70 42.5146
R21279 minus.n33 minus.n9 42.5146
R21280 minus.n40 minus.n39 42.5146
R21281 minus.n77 minus.n76 40.6041
R21282 minus.n16 minus.n15 40.6041
R21283 minus.n102 minus.n101 38.6395
R21284 minus.n90 minus.n70 38.6395
R21285 minus.n29 minus.n9 38.6395
R21286 minus.n41 minus.n40 38.6395
R21287 minus.n122 minus.n121 35.4191
R21288 minus.n112 minus.n64 34.7644
R21289 minus.n83 minus.n82 34.7644
R21290 minus.n22 minus.n21 34.7644
R21291 minus.n51 minus.n3 34.7644
R21292 minus.n114 minus.n113 21.8872
R21293 minus.n79 minus.n74 21.8872
R21294 minus.n18 minus.n13 21.8872
R21295 minus.n53 minus.n52 21.8872
R21296 minus.n105 minus.n66 19.9199
R21297 minus.n89 minus.n88 19.9199
R21298 minus.n28 minus.n27 19.9199
R21299 minus.n44 minus.n5 19.9199
R21300 minus.n124 minus.t0 19.8005
R21301 minus.n124 minus.t2 19.8005
R21302 minus.n123 minus.t4 19.8005
R21303 minus.n123 minus.t3 19.8005
R21304 minus.n97 minus.n68 17.9525
R21305 minus.n96 minus.n95 17.9525
R21306 minus.n35 minus.n34 17.9525
R21307 minus.n36 minus.n7 17.9525
R21308 minus.n107 minus.n106 15.9852
R21309 minus.n87 minus.n72 15.9852
R21310 minus.n26 minus.n11 15.9852
R21311 minus.n46 minus.n45 15.9852
R21312 minus.n115 minus.n62 14.0178
R21313 minus.n78 minus.n77 14.0178
R21314 minus.n17 minus.n16 14.0178
R21315 minus.n54 minus.n1 14.0178
R21316 minus.n122 minus.n60 12.1501
R21317 minus minus.n127 10.9162
R21318 minus.n118 minus.n62 10.575
R21319 minus.n57 minus.n1 10.575
R21320 minus.n120 minus.n119 9.49444
R21321 minus.n59 minus.n58 9.49444
R21322 minus.n108 minus.n107 8.60764
R21323 minus.n84 minus.n72 8.60764
R21324 minus.n23 minus.n11 8.60764
R21325 minus.n47 minus.n46 8.60764
R21326 minus.n100 minus.n68 6.6403
R21327 minus.n95 minus.n94 6.6403
R21328 minus.n34 minus.n33 6.6403
R21329 minus.n39 minus.n7 6.6403
R21330 minus.n127 minus.n126 4.80222
R21331 minus.n102 minus.n66 4.67295
R21332 minus.n90 minus.n89 4.67295
R21333 minus.n29 minus.n28 4.67295
R21334 minus.n41 minus.n5 4.67295
R21335 minus.n113 minus.n112 2.7056
R21336 minus.n82 minus.n74 2.7056
R21337 minus.n21 minus.n13 2.7056
R21338 minus.n52 minus.n51 2.7056
R21339 minus.n127 minus.n122 0.972091
R21340 minus.n126 minus.n125 0.716017
R21341 minus.n121 minus.n61 0.189894
R21342 minus.n117 minus.n61 0.189894
R21343 minus.n117 minus.n116 0.189894
R21344 minus.n116 minus.n63 0.189894
R21345 minus.n111 minus.n63 0.189894
R21346 minus.n111 minus.n110 0.189894
R21347 minus.n110 minus.n109 0.189894
R21348 minus.n109 minus.n65 0.189894
R21349 minus.n104 minus.n65 0.189894
R21350 minus.n104 minus.n103 0.189894
R21351 minus.n103 minus.n67 0.189894
R21352 minus.n99 minus.n67 0.189894
R21353 minus.n99 minus.n98 0.189894
R21354 minus.n98 minus.n69 0.189894
R21355 minus.n93 minus.n69 0.189894
R21356 minus.n93 minus.n92 0.189894
R21357 minus.n92 minus.n91 0.189894
R21358 minus.n91 minus.n71 0.189894
R21359 minus.n86 minus.n71 0.189894
R21360 minus.n86 minus.n85 0.189894
R21361 minus.n85 minus.n73 0.189894
R21362 minus.n81 minus.n73 0.189894
R21363 minus.n81 minus.n80 0.189894
R21364 minus.n80 minus.n75 0.189894
R21365 minus.n19 minus.n14 0.189894
R21366 minus.n20 minus.n19 0.189894
R21367 minus.n20 minus.n12 0.189894
R21368 minus.n24 minus.n12 0.189894
R21369 minus.n25 minus.n24 0.189894
R21370 minus.n25 minus.n10 0.189894
R21371 minus.n30 minus.n10 0.189894
R21372 minus.n31 minus.n30 0.189894
R21373 minus.n32 minus.n31 0.189894
R21374 minus.n32 minus.n8 0.189894
R21375 minus.n37 minus.n8 0.189894
R21376 minus.n38 minus.n37 0.189894
R21377 minus.n38 minus.n6 0.189894
R21378 minus.n42 minus.n6 0.189894
R21379 minus.n43 minus.n42 0.189894
R21380 minus.n43 minus.n4 0.189894
R21381 minus.n48 minus.n4 0.189894
R21382 minus.n49 minus.n48 0.189894
R21383 minus.n50 minus.n49 0.189894
R21384 minus.n50 minus.n2 0.189894
R21385 minus.n55 minus.n2 0.189894
R21386 minus.n56 minus.n55 0.189894
R21387 minus.n56 minus.n0 0.189894
R21388 minus.n60 minus.n0 0.189894
R21389 diffpairibias.n0 diffpairibias.t18 436.822
R21390 diffpairibias.n21 diffpairibias.t19 435.479
R21391 diffpairibias.n20 diffpairibias.t16 435.479
R21392 diffpairibias.n19 diffpairibias.t17 435.479
R21393 diffpairibias.n18 diffpairibias.t21 435.479
R21394 diffpairibias.n0 diffpairibias.t22 435.479
R21395 diffpairibias.n1 diffpairibias.t20 435.479
R21396 diffpairibias.n2 diffpairibias.t23 435.479
R21397 diffpairibias.n10 diffpairibias.t0 377.536
R21398 diffpairibias.n10 diffpairibias.t8 376.193
R21399 diffpairibias.n11 diffpairibias.t10 376.193
R21400 diffpairibias.n12 diffpairibias.t6 376.193
R21401 diffpairibias.n13 diffpairibias.t2 376.193
R21402 diffpairibias.n14 diffpairibias.t12 376.193
R21403 diffpairibias.n15 diffpairibias.t4 376.193
R21404 diffpairibias.n16 diffpairibias.t14 376.193
R21405 diffpairibias.n3 diffpairibias.t1 113.368
R21406 diffpairibias.n3 diffpairibias.t9 112.698
R21407 diffpairibias.n4 diffpairibias.t11 112.698
R21408 diffpairibias.n5 diffpairibias.t7 112.698
R21409 diffpairibias.n6 diffpairibias.t3 112.698
R21410 diffpairibias.n7 diffpairibias.t13 112.698
R21411 diffpairibias.n8 diffpairibias.t5 112.698
R21412 diffpairibias.n9 diffpairibias.t15 112.698
R21413 diffpairibias.n17 diffpairibias.n16 4.77242
R21414 diffpairibias.n17 diffpairibias.n9 4.30807
R21415 diffpairibias.n18 diffpairibias.n17 4.13945
R21416 diffpairibias.n16 diffpairibias.n15 1.34352
R21417 diffpairibias.n15 diffpairibias.n14 1.34352
R21418 diffpairibias.n14 diffpairibias.n13 1.34352
R21419 diffpairibias.n13 diffpairibias.n12 1.34352
R21420 diffpairibias.n12 diffpairibias.n11 1.34352
R21421 diffpairibias.n11 diffpairibias.n10 1.34352
R21422 diffpairibias.n2 diffpairibias.n1 1.34352
R21423 diffpairibias.n1 diffpairibias.n0 1.34352
R21424 diffpairibias.n19 diffpairibias.n18 1.34352
R21425 diffpairibias.n20 diffpairibias.n19 1.34352
R21426 diffpairibias.n21 diffpairibias.n20 1.34352
R21427 diffpairibias.n22 diffpairibias.n21 0.862419
R21428 diffpairibias diffpairibias.n22 0.684875
R21429 diffpairibias.n9 diffpairibias.n8 0.672012
R21430 diffpairibias.n8 diffpairibias.n7 0.672012
R21431 diffpairibias.n7 diffpairibias.n6 0.672012
R21432 diffpairibias.n6 diffpairibias.n5 0.672012
R21433 diffpairibias.n5 diffpairibias.n4 0.672012
R21434 diffpairibias.n4 diffpairibias.n3 0.672012
R21435 diffpairibias.n22 diffpairibias.n2 0.190907
C0 minus diffpairibias 5.39e-19
C1 commonsourceibias output 0.006808f
C2 vdd plus 0.072837f
C3 CSoutput minus 2.25384f
C4 plus diffpairibias 4.4e-19
C5 commonsourceibias outputibias 0.003832f
C6 vdd commonsourceibias 0.004218f
C7 CSoutput plus 0.874948f
C8 commonsourceibias diffpairibias 0.06482f
C9 CSoutput commonsourceibias 41.846302f
C10 minus plus 9.674179f
C11 minus commonsourceibias 0.515277f
C12 plus commonsourceibias 0.49873f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13881f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 67.6707f
C18 diffpairibias gnd 48.964737f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.143619p
C22 plus gnd 37.5619f
C23 minus gnd 28.67481f
C24 CSoutput gnd 0.106998p
C25 vdd gnd 0.344772p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.031832f
C74 minus.t13 gnd 0.535246f
C75 minus.n1 gnd 0.216477f
C76 minus.n2 gnd 0.031832f
C77 minus.t11 gnd 0.535246f
C78 minus.n3 gnd 0.027201f
C79 minus.n4 gnd 0.031832f
C80 minus.t17 gnd 0.535246f
C81 minus.t24 gnd 0.535246f
C82 minus.n5 gnd 0.216477f
C83 minus.n6 gnd 0.031832f
C84 minus.t21 gnd 0.535246f
C85 minus.n7 gnd 0.216477f
C86 minus.n8 gnd 0.031832f
C87 minus.t27 gnd 0.535246f
C88 minus.n9 gnd 0.025872f
C89 minus.n10 gnd 0.031832f
C90 minus.t26 gnd 0.535246f
C91 minus.t5 gnd 0.535246f
C92 minus.n11 gnd 0.216477f
C93 minus.n12 gnd 0.031832f
C94 minus.t9 gnd 0.535246f
C95 minus.n13 gnd 0.216477f
C96 minus.n14 gnd 0.135091f
C97 minus.t14 gnd 0.535246f
C98 minus.t20 gnd 0.59877f
C99 minus.n15 gnd 0.253084f
C100 minus.n16 gnd 0.247907f
C101 minus.n17 gnd 0.040787f
C102 minus.n18 gnd 0.036021f
C103 minus.n19 gnd 0.031832f
C104 minus.n20 gnd 0.031832f
C105 minus.n21 gnd 0.038039f
C106 minus.n22 gnd 0.027201f
C107 minus.n23 gnd 0.041457f
C108 minus.n24 gnd 0.031832f
C109 minus.n25 gnd 0.031832f
C110 minus.n26 gnd 0.039596f
C111 minus.n27 gnd 0.037213f
C112 minus.n28 gnd 0.216477f
C113 minus.n29 gnd 0.039874f
C114 minus.n30 gnd 0.031832f
C115 minus.n31 gnd 0.031832f
C116 minus.n32 gnd 0.031832f
C117 minus.n33 gnd 0.04095f
C118 minus.n34 gnd 0.216477f
C119 minus.n35 gnd 0.038404f
C120 minus.n36 gnd 0.038404f
C121 minus.n37 gnd 0.031832f
C122 minus.n38 gnd 0.031832f
C123 minus.n39 gnd 0.04095f
C124 minus.n40 gnd 0.025872f
C125 minus.n41 gnd 0.039874f
C126 minus.n42 gnd 0.031832f
C127 minus.n43 gnd 0.031832f
C128 minus.n44 gnd 0.037213f
C129 minus.n45 gnd 0.039596f
C130 minus.n46 gnd 0.216477f
C131 minus.n47 gnd 0.041457f
C132 minus.n48 gnd 0.031832f
C133 minus.n49 gnd 0.031832f
C134 minus.n50 gnd 0.031832f
C135 minus.n51 gnd 0.038039f
C136 minus.n52 gnd 0.216477f
C137 minus.n53 gnd 0.036021f
C138 minus.n54 gnd 0.040787f
C139 minus.n55 gnd 0.031832f
C140 minus.n56 gnd 0.031832f
C141 minus.n57 gnd 0.041526f
C142 minus.n58 gnd 0.011569f
C143 minus.t10 gnd 0.578869f
C144 minus.n59 gnd 0.250644f
C145 minus.n60 gnd 0.372897f
C146 minus.n61 gnd 0.031832f
C147 minus.t8 gnd 0.578869f
C148 minus.t12 gnd 0.535246f
C149 minus.n62 gnd 0.216477f
C150 minus.n63 gnd 0.031832f
C151 minus.t18 gnd 0.535246f
C152 minus.n64 gnd 0.027201f
C153 minus.n65 gnd 0.031832f
C154 minus.t25 gnd 0.535246f
C155 minus.t22 gnd 0.535246f
C156 minus.n66 gnd 0.216477f
C157 minus.n67 gnd 0.031832f
C158 minus.t19 gnd 0.535246f
C159 minus.n68 gnd 0.216477f
C160 minus.n69 gnd 0.031832f
C161 minus.t7 gnd 0.535246f
C162 minus.n70 gnd 0.025872f
C163 minus.n71 gnd 0.031832f
C164 minus.t6 gnd 0.535246f
C165 minus.t16 gnd 0.535246f
C166 minus.n72 gnd 0.216477f
C167 minus.n73 gnd 0.031832f
C168 minus.t15 gnd 0.535246f
C169 minus.n74 gnd 0.216477f
C170 minus.n75 gnd 0.135091f
C171 minus.t23 gnd 0.535246f
C172 minus.t28 gnd 0.59877f
C173 minus.n76 gnd 0.253084f
C174 minus.n77 gnd 0.247907f
C175 minus.n78 gnd 0.040787f
C176 minus.n79 gnd 0.036021f
C177 minus.n80 gnd 0.031832f
C178 minus.n81 gnd 0.031832f
C179 minus.n82 gnd 0.038039f
C180 minus.n83 gnd 0.027201f
C181 minus.n84 gnd 0.041457f
C182 minus.n85 gnd 0.031832f
C183 minus.n86 gnd 0.031832f
C184 minus.n87 gnd 0.039596f
C185 minus.n88 gnd 0.037213f
C186 minus.n89 gnd 0.216477f
C187 minus.n90 gnd 0.039874f
C188 minus.n91 gnd 0.031832f
C189 minus.n92 gnd 0.031832f
C190 minus.n93 gnd 0.031832f
C191 minus.n94 gnd 0.04095f
C192 minus.n95 gnd 0.216477f
C193 minus.n96 gnd 0.038404f
C194 minus.n97 gnd 0.038404f
C195 minus.n98 gnd 0.031832f
C196 minus.n99 gnd 0.031832f
C197 minus.n100 gnd 0.04095f
C198 minus.n101 gnd 0.025872f
C199 minus.n102 gnd 0.039874f
C200 minus.n103 gnd 0.031832f
C201 minus.n104 gnd 0.031832f
C202 minus.n105 gnd 0.037213f
C203 minus.n106 gnd 0.039596f
C204 minus.n107 gnd 0.216477f
C205 minus.n108 gnd 0.041457f
C206 minus.n109 gnd 0.031832f
C207 minus.n110 gnd 0.031832f
C208 minus.n111 gnd 0.031832f
C209 minus.n112 gnd 0.038039f
C210 minus.n113 gnd 0.216477f
C211 minus.n114 gnd 0.036021f
C212 minus.n115 gnd 0.040787f
C213 minus.n116 gnd 0.031832f
C214 minus.n117 gnd 0.031832f
C215 minus.n118 gnd 0.041526f
C216 minus.n119 gnd 0.011569f
C217 minus.n120 gnd 0.250644f
C218 minus.n121 gnd 1.16121f
C219 minus.n122 gnd 1.70573f
C220 minus.t4 gnd 0.009813f
C221 minus.t3 gnd 0.009813f
C222 minus.n123 gnd 0.032267f
C223 minus.t0 gnd 0.009813f
C224 minus.t2 gnd 0.009813f
C225 minus.n124 gnd 0.031825f
C226 minus.n125 gnd 0.271609f
C227 minus.t1 gnd 0.054617f
C228 minus.n126 gnd 0.148215f
C229 minus.n127 gnd 1.6183f
C230 output.t9 gnd 0.464308f
C231 output.t15 gnd 0.044422f
C232 output.t19 gnd 0.044422f
C233 output.n0 gnd 0.364624f
C234 output.n1 gnd 0.614102f
C235 output.t7 gnd 0.044422f
C236 output.t11 gnd 0.044422f
C237 output.n2 gnd 0.364624f
C238 output.n3 gnd 0.350265f
C239 output.t12 gnd 0.044422f
C240 output.t17 gnd 0.044422f
C241 output.n4 gnd 0.364624f
C242 output.n5 gnd 0.350265f
C243 output.t5 gnd 0.044422f
C244 output.t13 gnd 0.044422f
C245 output.n6 gnd 0.364624f
C246 output.n7 gnd 0.350265f
C247 output.t16 gnd 0.044422f
C248 output.t14 gnd 0.044422f
C249 output.n8 gnd 0.364624f
C250 output.n9 gnd 0.350265f
C251 output.t4 gnd 0.044422f
C252 output.t6 gnd 0.044422f
C253 output.n10 gnd 0.364624f
C254 output.n11 gnd 0.350265f
C255 output.t8 gnd 0.044422f
C256 output.t18 gnd 0.044422f
C257 output.n12 gnd 0.364624f
C258 output.n13 gnd 0.350265f
C259 output.t10 gnd 0.462979f
C260 output.n14 gnd 0.28994f
C261 output.n15 gnd 0.015803f
C262 output.n16 gnd 0.011243f
C263 output.n17 gnd 0.006041f
C264 output.n18 gnd 0.01428f
C265 output.n19 gnd 0.006397f
C266 output.n20 gnd 0.011243f
C267 output.n21 gnd 0.006041f
C268 output.n22 gnd 0.01428f
C269 output.n23 gnd 0.006397f
C270 output.n24 gnd 0.048111f
C271 output.t2 gnd 0.023274f
C272 output.n25 gnd 0.01071f
C273 output.n26 gnd 0.008435f
C274 output.n27 gnd 0.006041f
C275 output.n28 gnd 0.267512f
C276 output.n29 gnd 0.011243f
C277 output.n30 gnd 0.006041f
C278 output.n31 gnd 0.006397f
C279 output.n32 gnd 0.01428f
C280 output.n33 gnd 0.01428f
C281 output.n34 gnd 0.006397f
C282 output.n35 gnd 0.006041f
C283 output.n36 gnd 0.011243f
C284 output.n37 gnd 0.011243f
C285 output.n38 gnd 0.006041f
C286 output.n39 gnd 0.006397f
C287 output.n40 gnd 0.01428f
C288 output.n41 gnd 0.030913f
C289 output.n42 gnd 0.006397f
C290 output.n43 gnd 0.006041f
C291 output.n44 gnd 0.025987f
C292 output.n45 gnd 0.097665f
C293 output.n46 gnd 0.015803f
C294 output.n47 gnd 0.011243f
C295 output.n48 gnd 0.006041f
C296 output.n49 gnd 0.01428f
C297 output.n50 gnd 0.006397f
C298 output.n51 gnd 0.011243f
C299 output.n52 gnd 0.006041f
C300 output.n53 gnd 0.01428f
C301 output.n54 gnd 0.006397f
C302 output.n55 gnd 0.048111f
C303 output.t1 gnd 0.023274f
C304 output.n56 gnd 0.01071f
C305 output.n57 gnd 0.008435f
C306 output.n58 gnd 0.006041f
C307 output.n59 gnd 0.267512f
C308 output.n60 gnd 0.011243f
C309 output.n61 gnd 0.006041f
C310 output.n62 gnd 0.006397f
C311 output.n63 gnd 0.01428f
C312 output.n64 gnd 0.01428f
C313 output.n65 gnd 0.006397f
C314 output.n66 gnd 0.006041f
C315 output.n67 gnd 0.011243f
C316 output.n68 gnd 0.011243f
C317 output.n69 gnd 0.006041f
C318 output.n70 gnd 0.006397f
C319 output.n71 gnd 0.01428f
C320 output.n72 gnd 0.030913f
C321 output.n73 gnd 0.006397f
C322 output.n74 gnd 0.006041f
C323 output.n75 gnd 0.025987f
C324 output.n76 gnd 0.09306f
C325 output.n77 gnd 1.65264f
C326 output.n78 gnd 0.015803f
C327 output.n79 gnd 0.011243f
C328 output.n80 gnd 0.006041f
C329 output.n81 gnd 0.01428f
C330 output.n82 gnd 0.006397f
C331 output.n83 gnd 0.011243f
C332 output.n84 gnd 0.006041f
C333 output.n85 gnd 0.01428f
C334 output.n86 gnd 0.006397f
C335 output.n87 gnd 0.048111f
C336 output.t3 gnd 0.023274f
C337 output.n88 gnd 0.01071f
C338 output.n89 gnd 0.008435f
C339 output.n90 gnd 0.006041f
C340 output.n91 gnd 0.267512f
C341 output.n92 gnd 0.011243f
C342 output.n93 gnd 0.006041f
C343 output.n94 gnd 0.006397f
C344 output.n95 gnd 0.01428f
C345 output.n96 gnd 0.01428f
C346 output.n97 gnd 0.006397f
C347 output.n98 gnd 0.006041f
C348 output.n99 gnd 0.011243f
C349 output.n100 gnd 0.011243f
C350 output.n101 gnd 0.006041f
C351 output.n102 gnd 0.006397f
C352 output.n103 gnd 0.01428f
C353 output.n104 gnd 0.030913f
C354 output.n105 gnd 0.006397f
C355 output.n106 gnd 0.006041f
C356 output.n107 gnd 0.025987f
C357 output.n108 gnd 0.09306f
C358 output.n109 gnd 0.713089f
C359 output.n110 gnd 0.015803f
C360 output.n111 gnd 0.011243f
C361 output.n112 gnd 0.006041f
C362 output.n113 gnd 0.01428f
C363 output.n114 gnd 0.006397f
C364 output.n115 gnd 0.011243f
C365 output.n116 gnd 0.006041f
C366 output.n117 gnd 0.01428f
C367 output.n118 gnd 0.006397f
C368 output.n119 gnd 0.048111f
C369 output.t0 gnd 0.023274f
C370 output.n120 gnd 0.01071f
C371 output.n121 gnd 0.008435f
C372 output.n122 gnd 0.006041f
C373 output.n123 gnd 0.267512f
C374 output.n124 gnd 0.011243f
C375 output.n125 gnd 0.006041f
C376 output.n126 gnd 0.006397f
C377 output.n127 gnd 0.01428f
C378 output.n128 gnd 0.01428f
C379 output.n129 gnd 0.006397f
C380 output.n130 gnd 0.006041f
C381 output.n131 gnd 0.011243f
C382 output.n132 gnd 0.011243f
C383 output.n133 gnd 0.006041f
C384 output.n134 gnd 0.006397f
C385 output.n135 gnd 0.01428f
C386 output.n136 gnd 0.030913f
C387 output.n137 gnd 0.006397f
C388 output.n138 gnd 0.006041f
C389 output.n139 gnd 0.025987f
C390 output.n140 gnd 0.09306f
C391 output.n141 gnd 1.67353f
C392 outputibias.t10 gnd 0.11477f
C393 outputibias.t9 gnd 0.115567f
C394 outputibias.n0 gnd 0.130108f
C395 outputibias.n1 gnd 0.001372f
C396 outputibias.n2 gnd 9.76e-19
C397 outputibias.n3 gnd 5.24e-19
C398 outputibias.n4 gnd 0.001239f
C399 outputibias.n5 gnd 5.55e-19
C400 outputibias.n6 gnd 9.76e-19
C401 outputibias.n7 gnd 5.24e-19
C402 outputibias.n8 gnd 0.001239f
C403 outputibias.n9 gnd 5.55e-19
C404 outputibias.n10 gnd 0.004176f
C405 outputibias.t5 gnd 0.00202f
C406 outputibias.n11 gnd 9.3e-19
C407 outputibias.n12 gnd 7.32e-19
C408 outputibias.n13 gnd 5.24e-19
C409 outputibias.n14 gnd 0.02322f
C410 outputibias.n15 gnd 9.76e-19
C411 outputibias.n16 gnd 5.24e-19
C412 outputibias.n17 gnd 5.55e-19
C413 outputibias.n18 gnd 0.001239f
C414 outputibias.n19 gnd 0.001239f
C415 outputibias.n20 gnd 5.55e-19
C416 outputibias.n21 gnd 5.24e-19
C417 outputibias.n22 gnd 9.76e-19
C418 outputibias.n23 gnd 9.76e-19
C419 outputibias.n24 gnd 5.24e-19
C420 outputibias.n25 gnd 5.55e-19
C421 outputibias.n26 gnd 0.001239f
C422 outputibias.n27 gnd 0.002683f
C423 outputibias.n28 gnd 5.55e-19
C424 outputibias.n29 gnd 5.24e-19
C425 outputibias.n30 gnd 0.002256f
C426 outputibias.n31 gnd 0.005781f
C427 outputibias.n32 gnd 0.001372f
C428 outputibias.n33 gnd 9.76e-19
C429 outputibias.n34 gnd 5.24e-19
C430 outputibias.n35 gnd 0.001239f
C431 outputibias.n36 gnd 5.55e-19
C432 outputibias.n37 gnd 9.76e-19
C433 outputibias.n38 gnd 5.24e-19
C434 outputibias.n39 gnd 0.001239f
C435 outputibias.n40 gnd 5.55e-19
C436 outputibias.n41 gnd 0.004176f
C437 outputibias.t7 gnd 0.00202f
C438 outputibias.n42 gnd 9.3e-19
C439 outputibias.n43 gnd 7.32e-19
C440 outputibias.n44 gnd 5.24e-19
C441 outputibias.n45 gnd 0.02322f
C442 outputibias.n46 gnd 9.76e-19
C443 outputibias.n47 gnd 5.24e-19
C444 outputibias.n48 gnd 5.55e-19
C445 outputibias.n49 gnd 0.001239f
C446 outputibias.n50 gnd 0.001239f
C447 outputibias.n51 gnd 5.55e-19
C448 outputibias.n52 gnd 5.24e-19
C449 outputibias.n53 gnd 9.76e-19
C450 outputibias.n54 gnd 9.76e-19
C451 outputibias.n55 gnd 5.24e-19
C452 outputibias.n56 gnd 5.55e-19
C453 outputibias.n57 gnd 0.001239f
C454 outputibias.n58 gnd 0.002683f
C455 outputibias.n59 gnd 5.55e-19
C456 outputibias.n60 gnd 5.24e-19
C457 outputibias.n61 gnd 0.002256f
C458 outputibias.n62 gnd 0.005197f
C459 outputibias.n63 gnd 0.121892f
C460 outputibias.n64 gnd 0.001372f
C461 outputibias.n65 gnd 9.76e-19
C462 outputibias.n66 gnd 5.24e-19
C463 outputibias.n67 gnd 0.001239f
C464 outputibias.n68 gnd 5.55e-19
C465 outputibias.n69 gnd 9.76e-19
C466 outputibias.n70 gnd 5.24e-19
C467 outputibias.n71 gnd 0.001239f
C468 outputibias.n72 gnd 5.55e-19
C469 outputibias.n73 gnd 0.004176f
C470 outputibias.t1 gnd 0.00202f
C471 outputibias.n74 gnd 9.3e-19
C472 outputibias.n75 gnd 7.32e-19
C473 outputibias.n76 gnd 5.24e-19
C474 outputibias.n77 gnd 0.02322f
C475 outputibias.n78 gnd 9.76e-19
C476 outputibias.n79 gnd 5.24e-19
C477 outputibias.n80 gnd 5.55e-19
C478 outputibias.n81 gnd 0.001239f
C479 outputibias.n82 gnd 0.001239f
C480 outputibias.n83 gnd 5.55e-19
C481 outputibias.n84 gnd 5.24e-19
C482 outputibias.n85 gnd 9.76e-19
C483 outputibias.n86 gnd 9.76e-19
C484 outputibias.n87 gnd 5.24e-19
C485 outputibias.n88 gnd 5.55e-19
C486 outputibias.n89 gnd 0.001239f
C487 outputibias.n90 gnd 0.002683f
C488 outputibias.n91 gnd 5.55e-19
C489 outputibias.n92 gnd 5.24e-19
C490 outputibias.n93 gnd 0.002256f
C491 outputibias.n94 gnd 0.005197f
C492 outputibias.n95 gnd 0.064513f
C493 outputibias.n96 gnd 0.001372f
C494 outputibias.n97 gnd 9.76e-19
C495 outputibias.n98 gnd 5.24e-19
C496 outputibias.n99 gnd 0.001239f
C497 outputibias.n100 gnd 5.55e-19
C498 outputibias.n101 gnd 9.76e-19
C499 outputibias.n102 gnd 5.24e-19
C500 outputibias.n103 gnd 0.001239f
C501 outputibias.n104 gnd 5.55e-19
C502 outputibias.n105 gnd 0.004176f
C503 outputibias.t3 gnd 0.00202f
C504 outputibias.n106 gnd 9.3e-19
C505 outputibias.n107 gnd 7.32e-19
C506 outputibias.n108 gnd 5.24e-19
C507 outputibias.n109 gnd 0.02322f
C508 outputibias.n110 gnd 9.76e-19
C509 outputibias.n111 gnd 5.24e-19
C510 outputibias.n112 gnd 5.55e-19
C511 outputibias.n113 gnd 0.001239f
C512 outputibias.n114 gnd 0.001239f
C513 outputibias.n115 gnd 5.55e-19
C514 outputibias.n116 gnd 5.24e-19
C515 outputibias.n117 gnd 9.76e-19
C516 outputibias.n118 gnd 9.76e-19
C517 outputibias.n119 gnd 5.24e-19
C518 outputibias.n120 gnd 5.55e-19
C519 outputibias.n121 gnd 0.001239f
C520 outputibias.n122 gnd 0.002683f
C521 outputibias.n123 gnd 5.55e-19
C522 outputibias.n124 gnd 5.24e-19
C523 outputibias.n125 gnd 0.002256f
C524 outputibias.n126 gnd 0.005197f
C525 outputibias.n127 gnd 0.084814f
C526 outputibias.t2 gnd 0.108319f
C527 outputibias.t0 gnd 0.108319f
C528 outputibias.t6 gnd 0.108319f
C529 outputibias.t4 gnd 0.109238f
C530 outputibias.n128 gnd 0.134674f
C531 outputibias.n129 gnd 0.07244f
C532 outputibias.n130 gnd 0.079818f
C533 outputibias.n131 gnd 0.164901f
C534 outputibias.t11 gnd 0.11477f
C535 outputibias.n132 gnd 0.067481f
C536 outputibias.t8 gnd 0.11477f
C537 outputibias.n133 gnd 0.065115f
C538 outputibias.n134 gnd 0.029159f
C539 a_n3106_n452.t8 gnd 0.10001f
C540 a_n3106_n452.t19 gnd 1.03942f
C541 a_n3106_n452.n0 gnd 0.392946f
C542 a_n3106_n452.t33 gnd 1.29145f
C543 a_n3106_n452.n1 gnd 1.22854f
C544 a_n3106_n452.t47 gnd 1.03942f
C545 a_n3106_n452.n2 gnd 0.392946f
C546 a_n3106_n452.t39 gnd 0.10001f
C547 a_n3106_n452.t50 gnd 0.10001f
C548 a_n3106_n452.n3 gnd 0.816794f
C549 a_n3106_n452.n4 gnd 0.411618f
C550 a_n3106_n452.t34 gnd 0.10001f
C551 a_n3106_n452.t44 gnd 0.10001f
C552 a_n3106_n452.n5 gnd 0.816794f
C553 a_n3106_n452.n6 gnd 0.411618f
C554 a_n3106_n452.t37 gnd 0.10001f
C555 a_n3106_n452.t42 gnd 0.10001f
C556 a_n3106_n452.n7 gnd 0.816794f
C557 a_n3106_n452.n8 gnd 0.411618f
C558 a_n3106_n452.t1 gnd 0.10001f
C559 a_n3106_n452.t51 gnd 0.10001f
C560 a_n3106_n452.n9 gnd 0.816794f
C561 a_n3106_n452.n10 gnd 0.411618f
C562 a_n3106_n452.t36 gnd 0.10001f
C563 a_n3106_n452.t31 gnd 0.10001f
C564 a_n3106_n452.n11 gnd 0.816794f
C565 a_n3106_n452.n12 gnd 0.411618f
C566 a_n3106_n452.t48 gnd 1.03942f
C567 a_n3106_n452.n13 gnd 0.972974f
C568 a_n3106_n452.t54 gnd 1.29145f
C569 a_n3106_n452.n14 gnd 0.909591f
C570 a_n3106_n452.t52 gnd 1.29145f
C571 a_n3106_n452.n15 gnd 0.909591f
C572 a_n3106_n452.t40 gnd 1.29145f
C573 a_n3106_n452.n16 gnd 0.909591f
C574 a_n3106_n452.t41 gnd 1.29145f
C575 a_n3106_n452.n17 gnd 0.909591f
C576 a_n3106_n452.t55 gnd 1.29145f
C577 a_n3106_n452.n18 gnd 0.909591f
C578 a_n3106_n452.t0 gnd 1.29145f
C579 a_n3106_n452.n19 gnd 0.909591f
C580 a_n3106_n452.t53 gnd 1.29145f
C581 a_n3106_n452.n20 gnd 0.789472f
C582 a_n3106_n452.n21 gnd 0.948419f
C583 a_n3106_n452.t10 gnd 1.03941f
C584 a_n3106_n452.n22 gnd 0.645631f
C585 a_n3106_n452.t7 gnd 0.10001f
C586 a_n3106_n452.t24 gnd 0.10001f
C587 a_n3106_n452.n23 gnd 0.816793f
C588 a_n3106_n452.n24 gnd 0.41162f
C589 a_n3106_n452.t18 gnd 0.10001f
C590 a_n3106_n452.t22 gnd 0.10001f
C591 a_n3106_n452.n25 gnd 0.816793f
C592 a_n3106_n452.n26 gnd 0.41162f
C593 a_n3106_n452.t23 gnd 0.10001f
C594 a_n3106_n452.t11 gnd 0.10001f
C595 a_n3106_n452.n27 gnd 0.816793f
C596 a_n3106_n452.n28 gnd 0.41162f
C597 a_n3106_n452.t12 gnd 0.10001f
C598 a_n3106_n452.t3 gnd 0.10001f
C599 a_n3106_n452.n29 gnd 0.816793f
C600 a_n3106_n452.n30 gnd 0.41162f
C601 a_n3106_n452.t5 gnd 0.10001f
C602 a_n3106_n452.t21 gnd 0.10001f
C603 a_n3106_n452.n31 gnd 0.816793f
C604 a_n3106_n452.n32 gnd 0.41162f
C605 a_n3106_n452.t16 gnd 1.03941f
C606 a_n3106_n452.n33 gnd 0.39295f
C607 a_n3106_n452.t35 gnd 1.03941f
C608 a_n3106_n452.n34 gnd 0.39295f
C609 a_n3106_n452.t28 gnd 0.10001f
C610 a_n3106_n452.t29 gnd 0.10001f
C611 a_n3106_n452.n35 gnd 0.816793f
C612 a_n3106_n452.n36 gnd 0.41162f
C613 a_n3106_n452.t49 gnd 0.10001f
C614 a_n3106_n452.t38 gnd 0.10001f
C615 a_n3106_n452.n37 gnd 0.816793f
C616 a_n3106_n452.n38 gnd 0.41162f
C617 a_n3106_n452.t45 gnd 0.10001f
C618 a_n3106_n452.t27 gnd 0.10001f
C619 a_n3106_n452.n39 gnd 0.816793f
C620 a_n3106_n452.n40 gnd 0.41162f
C621 a_n3106_n452.t43 gnd 0.10001f
C622 a_n3106_n452.t46 gnd 0.10001f
C623 a_n3106_n452.n41 gnd 0.816793f
C624 a_n3106_n452.n42 gnd 0.41162f
C625 a_n3106_n452.t32 gnd 0.10001f
C626 a_n3106_n452.t30 gnd 0.10001f
C627 a_n3106_n452.n43 gnd 0.816793f
C628 a_n3106_n452.n44 gnd 0.41162f
C629 a_n3106_n452.t26 gnd 1.03941f
C630 a_n3106_n452.n45 gnd 0.645631f
C631 a_n3106_n452.n46 gnd 1.05146f
C632 a_n3106_n452.t6 gnd 1.03941f
C633 a_n3106_n452.n47 gnd 0.972978f
C634 a_n3106_n452.t4 gnd 0.10001f
C635 a_n3106_n452.t2 gnd 0.10001f
C636 a_n3106_n452.n48 gnd 0.816794f
C637 a_n3106_n452.n49 gnd 0.411618f
C638 a_n3106_n452.t15 gnd 0.10001f
C639 a_n3106_n452.t20 gnd 0.10001f
C640 a_n3106_n452.n50 gnd 0.816794f
C641 a_n3106_n452.n51 gnd 0.411618f
C642 a_n3106_n452.t13 gnd 0.10001f
C643 a_n3106_n452.t17 gnd 0.10001f
C644 a_n3106_n452.n52 gnd 0.816794f
C645 a_n3106_n452.n53 gnd 0.411618f
C646 a_n3106_n452.t9 gnd 0.10001f
C647 a_n3106_n452.t14 gnd 0.10001f
C648 a_n3106_n452.n54 gnd 0.816794f
C649 a_n3106_n452.n55 gnd 0.411618f
C650 a_n3106_n452.n56 gnd 0.411617f
C651 a_n3106_n452.n57 gnd 0.816796f
C652 a_n3106_n452.t25 gnd 0.10001f
C653 plus.n0 gnd 0.023652f
C654 plus.t20 gnd 0.430126f
C655 plus.t23 gnd 0.397712f
C656 plus.n1 gnd 0.160852f
C657 plus.n2 gnd 0.023652f
C658 plus.t6 gnd 0.397712f
C659 plus.n3 gnd 0.020211f
C660 plus.n4 gnd 0.023652f
C661 plus.t12 gnd 0.397712f
C662 plus.t8 gnd 0.397712f
C663 plus.n5 gnd 0.160852f
C664 plus.n6 gnd 0.023652f
C665 plus.t7 gnd 0.397712f
C666 plus.n7 gnd 0.160852f
C667 plus.n8 gnd 0.023652f
C668 plus.t19 gnd 0.397712f
C669 plus.n9 gnd 0.019224f
C670 plus.n10 gnd 0.023652f
C671 plus.t18 gnd 0.397712f
C672 plus.t27 gnd 0.397712f
C673 plus.n11 gnd 0.160852f
C674 plus.n12 gnd 0.023652f
C675 plus.t25 gnd 0.397712f
C676 plus.n13 gnd 0.160852f
C677 plus.n14 gnd 0.100378f
C678 plus.t9 gnd 0.397712f
C679 plus.t14 gnd 0.444913f
C680 plus.n15 gnd 0.188053f
C681 plus.n16 gnd 0.184206f
C682 plus.n17 gnd 0.030307f
C683 plus.n18 gnd 0.026765f
C684 plus.n19 gnd 0.023652f
C685 plus.n20 gnd 0.023652f
C686 plus.n21 gnd 0.028265f
C687 plus.n22 gnd 0.020211f
C688 plus.n23 gnd 0.030804f
C689 plus.n24 gnd 0.023652f
C690 plus.n25 gnd 0.023652f
C691 plus.n26 gnd 0.029422f
C692 plus.n27 gnd 0.027651f
C693 plus.n28 gnd 0.160852f
C694 plus.n29 gnd 0.029629f
C695 plus.n30 gnd 0.023652f
C696 plus.n31 gnd 0.023652f
C697 plus.n32 gnd 0.023652f
C698 plus.n33 gnd 0.030428f
C699 plus.n34 gnd 0.160852f
C700 plus.n35 gnd 0.028536f
C701 plus.n36 gnd 0.028536f
C702 plus.n37 gnd 0.023652f
C703 plus.n38 gnd 0.023652f
C704 plus.n39 gnd 0.030428f
C705 plus.n40 gnd 0.019224f
C706 plus.n41 gnd 0.029629f
C707 plus.n42 gnd 0.023652f
C708 plus.n43 gnd 0.023652f
C709 plus.n44 gnd 0.027651f
C710 plus.n45 gnd 0.029422f
C711 plus.n46 gnd 0.160852f
C712 plus.n47 gnd 0.030804f
C713 plus.n48 gnd 0.023652f
C714 plus.n49 gnd 0.023652f
C715 plus.n50 gnd 0.023652f
C716 plus.n51 gnd 0.028265f
C717 plus.n52 gnd 0.160852f
C718 plus.n53 gnd 0.026765f
C719 plus.n54 gnd 0.030307f
C720 plus.n55 gnd 0.023652f
C721 plus.n56 gnd 0.023652f
C722 plus.n57 gnd 0.030855f
C723 plus.n58 gnd 0.008596f
C724 plus.n59 gnd 0.18624f
C725 plus.n60 gnd 0.270994f
C726 plus.n61 gnd 0.023652f
C727 plus.t28 gnd 0.397712f
C728 plus.n62 gnd 0.160852f
C729 plus.n63 gnd 0.023652f
C730 plus.t26 gnd 0.397712f
C731 plus.n64 gnd 0.020211f
C732 plus.n65 gnd 0.023652f
C733 plus.t10 gnd 0.397712f
C734 plus.t15 gnd 0.397712f
C735 plus.n66 gnd 0.160852f
C736 plus.n67 gnd 0.023652f
C737 plus.t13 gnd 0.397712f
C738 plus.n68 gnd 0.160852f
C739 plus.n69 gnd 0.023652f
C740 plus.t17 gnd 0.397712f
C741 plus.n70 gnd 0.019224f
C742 plus.n71 gnd 0.023652f
C743 plus.t16 gnd 0.397712f
C744 plus.t21 gnd 0.397712f
C745 plus.n72 gnd 0.160852f
C746 plus.n73 gnd 0.023652f
C747 plus.t22 gnd 0.397712f
C748 plus.n74 gnd 0.160852f
C749 plus.n75 gnd 0.100378f
C750 plus.t5 gnd 0.397712f
C751 plus.t11 gnd 0.444913f
C752 plus.n76 gnd 0.188053f
C753 plus.n77 gnd 0.184206f
C754 plus.n78 gnd 0.030307f
C755 plus.n79 gnd 0.026765f
C756 plus.n80 gnd 0.023652f
C757 plus.n81 gnd 0.023652f
C758 plus.n82 gnd 0.028265f
C759 plus.n83 gnd 0.020211f
C760 plus.n84 gnd 0.030804f
C761 plus.n85 gnd 0.023652f
C762 plus.n86 gnd 0.023652f
C763 plus.n87 gnd 0.029422f
C764 plus.n88 gnd 0.027651f
C765 plus.n89 gnd 0.160852f
C766 plus.n90 gnd 0.029629f
C767 plus.n91 gnd 0.023652f
C768 plus.n92 gnd 0.023652f
C769 plus.n93 gnd 0.023652f
C770 plus.n94 gnd 0.030428f
C771 plus.n95 gnd 0.160852f
C772 plus.n96 gnd 0.028536f
C773 plus.n97 gnd 0.028536f
C774 plus.n98 gnd 0.023652f
C775 plus.n99 gnd 0.023652f
C776 plus.n100 gnd 0.030428f
C777 plus.n101 gnd 0.019224f
C778 plus.n102 gnd 0.029629f
C779 plus.n103 gnd 0.023652f
C780 plus.n104 gnd 0.023652f
C781 plus.n105 gnd 0.027651f
C782 plus.n106 gnd 0.029422f
C783 plus.n107 gnd 0.160852f
C784 plus.n108 gnd 0.030804f
C785 plus.n109 gnd 0.023652f
C786 plus.n110 gnd 0.023652f
C787 plus.n111 gnd 0.023652f
C788 plus.n112 gnd 0.028265f
C789 plus.n113 gnd 0.160852f
C790 plus.n114 gnd 0.026765f
C791 plus.n115 gnd 0.030307f
C792 plus.n116 gnd 0.023652f
C793 plus.n117 gnd 0.023652f
C794 plus.n118 gnd 0.030855f
C795 plus.n119 gnd 0.008596f
C796 plus.t24 gnd 0.430126f
C797 plus.n120 gnd 0.18624f
C798 plus.n121 gnd 0.853371f
C799 plus.n122 gnd 1.25804f
C800 plus.t1 gnd 0.040831f
C801 plus.t2 gnd 0.007291f
C802 plus.t4 gnd 0.007291f
C803 plus.n123 gnd 0.023647f
C804 plus.n124 gnd 0.183575f
C805 plus.t3 gnd 0.007291f
C806 plus.t0 gnd 0.007291f
C807 plus.n125 gnd 0.023647f
C808 plus.n126 gnd 0.137795f
C809 plus.n127 gnd 2.64316f
C810 a_n1808_13878.t11 gnd 0.185683f
C811 a_n1808_13878.t13 gnd 0.185683f
C812 a_n1808_13878.t17 gnd 0.185683f
C813 a_n1808_13878.n0 gnd 1.46451f
C814 a_n1808_13878.t8 gnd 0.185683f
C815 a_n1808_13878.t10 gnd 0.185683f
C816 a_n1808_13878.n1 gnd 1.46364f
C817 a_n1808_13878.t14 gnd 0.185683f
C818 a_n1808_13878.t9 gnd 0.185683f
C819 a_n1808_13878.n2 gnd 1.46209f
C820 a_n1808_13878.n3 gnd 2.04299f
C821 a_n1808_13878.t12 gnd 0.185683f
C822 a_n1808_13878.t19 gnd 0.185683f
C823 a_n1808_13878.n4 gnd 1.46209f
C824 a_n1808_13878.n5 gnd 3.70273f
C825 a_n1808_13878.t1 gnd 1.73864f
C826 a_n1808_13878.t4 gnd 0.185683f
C827 a_n1808_13878.t5 gnd 0.185683f
C828 a_n1808_13878.n6 gnd 1.30795f
C829 a_n1808_13878.n7 gnd 1.46144f
C830 a_n1808_13878.t0 gnd 1.73518f
C831 a_n1808_13878.n8 gnd 0.735417f
C832 a_n1808_13878.t3 gnd 1.73518f
C833 a_n1808_13878.n9 gnd 0.735417f
C834 a_n1808_13878.t6 gnd 0.185683f
C835 a_n1808_13878.t7 gnd 0.185683f
C836 a_n1808_13878.n10 gnd 1.30795f
C837 a_n1808_13878.n11 gnd 0.742539f
C838 a_n1808_13878.t2 gnd 1.73518f
C839 a_n1808_13878.n12 gnd 1.73174f
C840 a_n1808_13878.n13 gnd 2.52099f
C841 a_n1808_13878.t15 gnd 0.185683f
C842 a_n1808_13878.t16 gnd 0.185683f
C843 a_n1808_13878.n14 gnd 1.46209f
C844 a_n1808_13878.n15 gnd 1.80499f
C845 a_n1808_13878.n16 gnd 1.31424f
C846 a_n1808_13878.n17 gnd 1.46209f
C847 a_n1808_13878.t18 gnd 0.185683f
C848 a_n1986_8322.t0 gnd 38.672398f
C849 a_n1986_8322.t2 gnd 27.512402f
C850 a_n1986_8322.t3 gnd 19.268198f
C851 a_n1986_8322.t1 gnd 38.672398f
C852 a_n1986_8322.t13 gnd 0.875792f
C853 a_n1986_8322.t21 gnd 0.093533f
C854 a_n1986_8322.t16 gnd 0.093533f
C855 a_n1986_8322.n0 gnd 0.658844f
C856 a_n1986_8322.n1 gnd 0.736161f
C857 a_n1986_8322.t19 gnd 0.093533f
C858 a_n1986_8322.t18 gnd 0.093533f
C859 a_n1986_8322.n2 gnd 0.658844f
C860 a_n1986_8322.n3 gnd 0.374034f
C861 a_n1986_8322.t12 gnd 0.874048f
C862 a_n1986_8322.n4 gnd 1.39896f
C863 a_n1986_8322.t6 gnd 0.875792f
C864 a_n1986_8322.t10 gnd 0.093533f
C865 a_n1986_8322.t9 gnd 0.093533f
C866 a_n1986_8322.n5 gnd 0.658844f
C867 a_n1986_8322.n6 gnd 0.736161f
C868 a_n1986_8322.t4 gnd 0.874048f
C869 a_n1986_8322.n7 gnd 0.370446f
C870 a_n1986_8322.t7 gnd 0.874048f
C871 a_n1986_8322.n8 gnd 0.370446f
C872 a_n1986_8322.t5 gnd 0.093533f
C873 a_n1986_8322.t11 gnd 0.093533f
C874 a_n1986_8322.n9 gnd 0.658844f
C875 a_n1986_8322.n10 gnd 0.374034f
C876 a_n1986_8322.t8 gnd 0.874048f
C877 a_n1986_8322.n11 gnd 0.872317f
C878 a_n1986_8322.n12 gnd 1.59071f
C879 a_n1986_8322.n13 gnd 3.20172f
C880 a_n1986_8322.t15 gnd 0.874048f
C881 a_n1986_8322.n14 gnd 0.76652f
C882 a_n1986_8322.t14 gnd 0.093533f
C883 a_n1986_8322.t23 gnd 0.093533f
C884 a_n1986_8322.n15 gnd 0.658844f
C885 a_n1986_8322.n16 gnd 0.374034f
C886 a_n1986_8322.t20 gnd 0.093533f
C887 a_n1986_8322.t17 gnd 0.093533f
C888 a_n1986_8322.n17 gnd 0.658844f
C889 a_n1986_8322.n18 gnd 0.736159f
C890 a_n1986_8322.t22 gnd 0.875794f
C891 a_n2848_n452.n0 gnd 0.492472f
C892 a_n2848_n452.n1 gnd 0.664435f
C893 a_n2848_n452.n2 gnd 0.215942f
C894 a_n2848_n452.n3 gnd 0.282512f
C895 a_n2848_n452.n4 gnd 0.438486f
C896 a_n2848_n452.n5 gnd 2.99175f
C897 a_n2848_n452.n6 gnd 0.526038f
C898 a_n2848_n452.n7 gnd 0.204894f
C899 a_n2848_n452.n8 gnd 0.150908f
C900 a_n2848_n452.n9 gnd 0.23718f
C901 a_n2848_n452.n10 gnd 0.183194f
C902 a_n2848_n452.n11 gnd 0.204894f
C903 a_n2848_n452.n12 gnd 0.150908f
C904 a_n2848_n452.n13 gnd 0.580023f
C905 a_n2848_n452.n14 gnd 0.432289f
C906 a_n2848_n452.n15 gnd 0.215942f
C907 a_n2848_n452.n16 gnd 0.492472f
C908 a_n2848_n452.n17 gnd 0.282512f
C909 a_n2848_n452.n18 gnd 0.438486f
C910 a_n2848_n452.n19 gnd 0.215942f
C911 a_n2848_n452.n20 gnd 0.731535f
C912 a_n2848_n452.n21 gnd 0.282512f
C913 a_n2848_n452.n22 gnd 1.77783f
C914 a_n2848_n452.n23 gnd 1.17886f
C915 a_n2848_n452.n24 gnd 1.91568f
C916 a_n2848_n452.n25 gnd 0.377489f
C917 a_n2848_n452.n26 gnd 3.11576f
C918 a_n2848_n452.n27 gnd 0.377488f
C919 a_n2848_n452.n28 gnd 3.20158f
C920 a_n2848_n452.n29 gnd 0.008361f
C921 a_n2848_n452.n31 gnd 0.285666f
C922 a_n2848_n452.n32 gnd 0.008361f
C923 a_n2848_n452.n34 gnd 0.285666f
C924 a_n2848_n452.n35 gnd 0.008361f
C925 a_n2848_n452.n36 gnd 0.28526f
C926 a_n2848_n452.n37 gnd 0.008361f
C927 a_n2848_n452.n38 gnd 0.28526f
C928 a_n2848_n452.n39 gnd 0.008361f
C929 a_n2848_n452.n40 gnd 0.28526f
C930 a_n2848_n452.n41 gnd 0.008361f
C931 a_n2848_n452.n42 gnd 1.33845f
C932 a_n2848_n452.n43 gnd 0.28526f
C933 a_n2848_n452.n45 gnd 0.285666f
C934 a_n2848_n452.n46 gnd 0.008361f
C935 a_n2848_n452.n48 gnd 0.285666f
C936 a_n2848_n452.n50 gnd 0.302425f
C937 a_n2848_n452.t24 gnd 0.14978f
C938 a_n2848_n452.t20 gnd 1.40246f
C939 a_n2848_n452.t40 gnd 0.14978f
C940 a_n2848_n452.t26 gnd 0.14978f
C941 a_n2848_n452.n51 gnd 1.05505f
C942 a_n2848_n452.t23 gnd 0.696704f
C943 a_n2848_n452.n52 gnd 0.306315f
C944 a_n2848_n452.t17 gnd 0.696704f
C945 a_n2848_n452.t39 gnd 0.696704f
C946 a_n2848_n452.t56 gnd 0.696704f
C947 a_n2848_n452.n53 gnd 0.306315f
C948 a_n2848_n452.t65 gnd 0.696704f
C949 a_n2848_n452.t71 gnd 0.696704f
C950 a_n2848_n452.t31 gnd 0.696704f
C951 a_n2848_n452.t33 gnd 0.696704f
C952 a_n2848_n452.t35 gnd 0.696704f
C953 a_n2848_n452.t21 gnd 0.696704f
C954 a_n2848_n452.t75 gnd 0.711378f
C955 a_n2848_n452.t58 gnd 0.696704f
C956 a_n2848_n452.t62 gnd 0.696704f
C957 a_n2848_n452.t52 gnd 0.696704f
C958 a_n2848_n452.n54 gnd 0.306315f
C959 a_n2848_n452.t67 gnd 0.696704f
C960 a_n2848_n452.t73 gnd 0.708223f
C961 a_n2848_n452.n55 gnd 0.308933f
C962 a_n2848_n452.n56 gnd 0.302425f
C963 a_n2848_n452.n57 gnd 0.308932f
C964 a_n2848_n452.t37 gnd 0.708223f
C965 a_n2848_n452.n58 gnd 0.308933f
C966 a_n2848_n452.t29 gnd 0.696704f
C967 a_n2848_n452.n59 gnd 0.302425f
C968 a_n2848_n452.n60 gnd 0.01225f
C969 a_n2848_n452.t9 gnd 0.116496f
C970 a_n2848_n452.t3 gnd 0.116496f
C971 a_n2848_n452.n61 gnd 1.03243f
C972 a_n2848_n452.t4 gnd 0.116496f
C973 a_n2848_n452.t45 gnd 0.116496f
C974 a_n2848_n452.n62 gnd 1.0294f
C975 a_n2848_n452.n63 gnd 0.912817f
C976 a_n2848_n452.t12 gnd 0.116496f
C977 a_n2848_n452.t41 gnd 0.116496f
C978 a_n2848_n452.n64 gnd 1.0294f
C979 a_n2848_n452.t5 gnd 0.116496f
C980 a_n2848_n452.t1 gnd 0.116496f
C981 a_n2848_n452.n65 gnd 1.03243f
C982 a_n2848_n452.t42 gnd 0.116496f
C983 a_n2848_n452.t7 gnd 0.116496f
C984 a_n2848_n452.n66 gnd 1.0294f
C985 a_n2848_n452.n67 gnd 0.912817f
C986 a_n2848_n452.t2 gnd 0.116496f
C987 a_n2848_n452.t15 gnd 0.116496f
C988 a_n2848_n452.n68 gnd 1.0294f
C989 a_n2848_n452.t44 gnd 0.116496f
C990 a_n2848_n452.t10 gnd 0.116496f
C991 a_n2848_n452.n69 gnd 1.0294f
C992 a_n2848_n452.n70 gnd 3.15028f
C993 a_n2848_n452.t6 gnd 0.116496f
C994 a_n2848_n452.t0 gnd 0.116496f
C995 a_n2848_n452.n71 gnd 1.0294f
C996 a_n2848_n452.n72 gnd 0.449443f
C997 a_n2848_n452.t47 gnd 0.116496f
C998 a_n2848_n452.t11 gnd 0.116496f
C999 a_n2848_n452.n73 gnd 1.0294f
C1000 a_n2848_n452.t46 gnd 0.116496f
C1001 a_n2848_n452.t43 gnd 0.116496f
C1002 a_n2848_n452.n74 gnd 1.03243f
C1003 a_n2848_n452.t16 gnd 0.116496f
C1004 a_n2848_n452.t13 gnd 0.116496f
C1005 a_n2848_n452.n75 gnd 1.0294f
C1006 a_n2848_n452.n76 gnd 0.912815f
C1007 a_n2848_n452.t14 gnd 0.116496f
C1008 a_n2848_n452.t8 gnd 0.116496f
C1009 a_n2848_n452.n77 gnd 1.0294f
C1010 a_n2848_n452.n78 gnd 0.2971f
C1011 a_n2848_n452.n79 gnd 0.01225f
C1012 a_n2848_n452.n80 gnd 0.296767f
C1013 a_n2848_n452.n81 gnd 0.531228f
C1014 a_n2848_n452.t38 gnd 1.40246f
C1015 a_n2848_n452.t30 gnd 0.14978f
C1016 a_n2848_n452.t22 gnd 0.14978f
C1017 a_n2848_n452.n82 gnd 1.05505f
C1018 a_n2848_n452.t36 gnd 0.14978f
C1019 a_n2848_n452.t34 gnd 0.14978f
C1020 a_n2848_n452.n83 gnd 1.05505f
C1021 a_n2848_n452.t32 gnd 1.39967f
C1022 a_n2848_n452.n84 gnd 1.14458f
C1023 a_n2848_n452.n85 gnd 0.786935f
C1024 a_n2848_n452.t57 gnd 0.696704f
C1025 a_n2848_n452.t66 gnd 0.696704f
C1026 a_n2848_n452.t48 gnd 0.696704f
C1027 a_n2848_n452.n86 gnd 0.306315f
C1028 a_n2848_n452.t68 gnd 0.696704f
C1029 a_n2848_n452.t53 gnd 0.696704f
C1030 a_n2848_n452.t54 gnd 0.696704f
C1031 a_n2848_n452.n87 gnd 0.306315f
C1032 a_n2848_n452.t72 gnd 0.696704f
C1033 a_n2848_n452.t61 gnd 0.696704f
C1034 a_n2848_n452.t60 gnd 0.696704f
C1035 a_n2848_n452.n88 gnd 0.306315f
C1036 a_n2848_n452.t64 gnd 0.696704f
C1037 a_n2848_n452.t55 gnd 0.696704f
C1038 a_n2848_n452.t49 gnd 0.696704f
C1039 a_n2848_n452.n89 gnd 0.306315f
C1040 a_n2848_n452.t69 gnd 0.708378f
C1041 a_n2848_n452.n90 gnd 0.302425f
C1042 a_n2848_n452.n91 gnd 0.296933f
C1043 a_n2848_n452.t74 gnd 0.708378f
C1044 a_n2848_n452.n92 gnd 0.302425f
C1045 a_n2848_n452.n93 gnd 0.296933f
C1046 a_n2848_n452.t63 gnd 0.708378f
C1047 a_n2848_n452.n94 gnd 0.302425f
C1048 a_n2848_n452.n95 gnd 0.296933f
C1049 a_n2848_n452.t59 gnd 0.708378f
C1050 a_n2848_n452.n96 gnd 0.302425f
C1051 a_n2848_n452.n97 gnd 0.296933f
C1052 a_n2848_n452.n98 gnd 1.0063f
C1053 a_n2848_n452.t70 gnd 0.711378f
C1054 a_n2848_n452.n99 gnd 0.308932f
C1055 a_n2848_n452.t50 gnd 0.696704f
C1056 a_n2848_n452.n100 gnd 0.302425f
C1057 a_n2848_n452.n101 gnd 0.308933f
C1058 a_n2848_n452.t51 gnd 0.708223f
C1059 a_n2848_n452.t19 gnd 0.711378f
C1060 a_n2848_n452.n102 gnd 0.308932f
C1061 a_n2848_n452.t25 gnd 0.696704f
C1062 a_n2848_n452.n103 gnd 0.302425f
C1063 a_n2848_n452.n104 gnd 0.308933f
C1064 a_n2848_n452.t27 gnd 0.708223f
C1065 a_n2848_n452.n105 gnd 1.13204f
C1066 a_n2848_n452.t28 gnd 1.39967f
C1067 a_n2848_n452.n106 gnd 1.05505f
C1068 a_n2848_n452.t18 gnd 0.14978f
C1069 vdd.t9 gnd 0.032933f
C1070 vdd.t102 gnd 0.032933f
C1071 vdd.n0 gnd 0.259746f
C1072 vdd.t94 gnd 0.032933f
C1073 vdd.t199 gnd 0.032933f
C1074 vdd.n1 gnd 0.259317f
C1075 vdd.n2 gnd 0.23914f
C1076 vdd.t106 gnd 0.032933f
C1077 vdd.t92 gnd 0.032933f
C1078 vdd.n3 gnd 0.259317f
C1079 vdd.n4 gnd 0.120942f
C1080 vdd.t195 gnd 0.032933f
C1081 vdd.t193 gnd 0.032933f
C1082 vdd.n5 gnd 0.259317f
C1083 vdd.n6 gnd 0.113482f
C1084 vdd.t96 gnd 0.032933f
C1085 vdd.t108 gnd 0.032933f
C1086 vdd.n7 gnd 0.259746f
C1087 vdd.t1 gnd 0.032933f
C1088 vdd.t197 gnd 0.032933f
C1089 vdd.n8 gnd 0.259317f
C1090 vdd.n9 gnd 0.23914f
C1091 vdd.t4 gnd 0.032933f
C1092 vdd.t12 gnd 0.032933f
C1093 vdd.n10 gnd 0.259317f
C1094 vdd.n11 gnd 0.120942f
C1095 vdd.t99 gnd 0.032933f
C1096 vdd.t6 gnd 0.032933f
C1097 vdd.n12 gnd 0.259317f
C1098 vdd.n13 gnd 0.113482f
C1099 vdd.n14 gnd 0.080229f
C1100 vdd.t177 gnd 0.018296f
C1101 vdd.t187 gnd 0.018296f
C1102 vdd.n15 gnd 0.168407f
C1103 vdd.t188 gnd 0.018296f
C1104 vdd.t182 gnd 0.018296f
C1105 vdd.n16 gnd 0.167914f
C1106 vdd.n17 gnd 0.292223f
C1107 vdd.t179 gnd 0.018296f
C1108 vdd.t189 gnd 0.018296f
C1109 vdd.n18 gnd 0.167914f
C1110 vdd.n19 gnd 0.120896f
C1111 vdd.t176 gnd 0.018296f
C1112 vdd.t181 gnd 0.018296f
C1113 vdd.n20 gnd 0.168407f
C1114 vdd.t190 gnd 0.018296f
C1115 vdd.t186 gnd 0.018296f
C1116 vdd.n21 gnd 0.167914f
C1117 vdd.n22 gnd 0.292223f
C1118 vdd.t184 gnd 0.018296f
C1119 vdd.t180 gnd 0.018296f
C1120 vdd.n23 gnd 0.167914f
C1121 vdd.n24 gnd 0.120896f
C1122 vdd.t178 gnd 0.018296f
C1123 vdd.t191 gnd 0.018296f
C1124 vdd.n25 gnd 0.167914f
C1125 vdd.t183 gnd 0.018296f
C1126 vdd.t185 gnd 0.018296f
C1127 vdd.n26 gnd 0.167914f
C1128 vdd.n27 gnd 18.208302f
C1129 vdd.n28 gnd 6.72294f
C1130 vdd.n29 gnd 0.00499f
C1131 vdd.n30 gnd 0.004631f
C1132 vdd.n31 gnd 0.002561f
C1133 vdd.n32 gnd 0.005881f
C1134 vdd.n33 gnd 0.002488f
C1135 vdd.n34 gnd 0.002635f
C1136 vdd.n35 gnd 0.004631f
C1137 vdd.n36 gnd 0.002488f
C1138 vdd.n37 gnd 0.005881f
C1139 vdd.n38 gnd 0.002635f
C1140 vdd.n39 gnd 0.004631f
C1141 vdd.n40 gnd 0.002488f
C1142 vdd.n41 gnd 0.004411f
C1143 vdd.n42 gnd 0.004424f
C1144 vdd.t115 gnd 0.012636f
C1145 vdd.n43 gnd 0.028114f
C1146 vdd.n44 gnd 0.146311f
C1147 vdd.n45 gnd 0.002488f
C1148 vdd.n46 gnd 0.002635f
C1149 vdd.n47 gnd 0.005881f
C1150 vdd.n48 gnd 0.005881f
C1151 vdd.n49 gnd 0.002635f
C1152 vdd.n50 gnd 0.002488f
C1153 vdd.n51 gnd 0.004631f
C1154 vdd.n52 gnd 0.004631f
C1155 vdd.n53 gnd 0.002488f
C1156 vdd.n54 gnd 0.002635f
C1157 vdd.n55 gnd 0.005881f
C1158 vdd.n56 gnd 0.005881f
C1159 vdd.n57 gnd 0.002635f
C1160 vdd.n58 gnd 0.002488f
C1161 vdd.n59 gnd 0.004631f
C1162 vdd.n60 gnd 0.004631f
C1163 vdd.n61 gnd 0.002488f
C1164 vdd.n62 gnd 0.002635f
C1165 vdd.n63 gnd 0.005881f
C1166 vdd.n64 gnd 0.005881f
C1167 vdd.n65 gnd 0.013905f
C1168 vdd.n66 gnd 0.002561f
C1169 vdd.n67 gnd 0.002488f
C1170 vdd.n68 gnd 0.011968f
C1171 vdd.n69 gnd 0.008356f
C1172 vdd.t167 gnd 0.029274f
C1173 vdd.t141 gnd 0.029274f
C1174 vdd.n70 gnd 0.201188f
C1175 vdd.n71 gnd 0.158204f
C1176 vdd.t174 gnd 0.029274f
C1177 vdd.t130 gnd 0.029274f
C1178 vdd.n72 gnd 0.201188f
C1179 vdd.n73 gnd 0.127669f
C1180 vdd.t160 gnd 0.029274f
C1181 vdd.t135 gnd 0.029274f
C1182 vdd.n74 gnd 0.201188f
C1183 vdd.n75 gnd 0.127669f
C1184 vdd.n76 gnd 0.00499f
C1185 vdd.n77 gnd 0.004631f
C1186 vdd.n78 gnd 0.002561f
C1187 vdd.n79 gnd 0.005881f
C1188 vdd.n80 gnd 0.002488f
C1189 vdd.n81 gnd 0.002635f
C1190 vdd.n82 gnd 0.004631f
C1191 vdd.n83 gnd 0.002488f
C1192 vdd.n84 gnd 0.005881f
C1193 vdd.n85 gnd 0.002635f
C1194 vdd.n86 gnd 0.004631f
C1195 vdd.n87 gnd 0.002488f
C1196 vdd.n88 gnd 0.004411f
C1197 vdd.n89 gnd 0.004424f
C1198 vdd.t173 gnd 0.012636f
C1199 vdd.n90 gnd 0.028114f
C1200 vdd.n91 gnd 0.146311f
C1201 vdd.n92 gnd 0.002488f
C1202 vdd.n93 gnd 0.002635f
C1203 vdd.n94 gnd 0.005881f
C1204 vdd.n95 gnd 0.005881f
C1205 vdd.n96 gnd 0.002635f
C1206 vdd.n97 gnd 0.002488f
C1207 vdd.n98 gnd 0.004631f
C1208 vdd.n99 gnd 0.004631f
C1209 vdd.n100 gnd 0.002488f
C1210 vdd.n101 gnd 0.002635f
C1211 vdd.n102 gnd 0.005881f
C1212 vdd.n103 gnd 0.005881f
C1213 vdd.n104 gnd 0.002635f
C1214 vdd.n105 gnd 0.002488f
C1215 vdd.n106 gnd 0.004631f
C1216 vdd.n107 gnd 0.004631f
C1217 vdd.n108 gnd 0.002488f
C1218 vdd.n109 gnd 0.002635f
C1219 vdd.n110 gnd 0.005881f
C1220 vdd.n111 gnd 0.005881f
C1221 vdd.n112 gnd 0.013905f
C1222 vdd.n113 gnd 0.002561f
C1223 vdd.n114 gnd 0.002488f
C1224 vdd.n115 gnd 0.011968f
C1225 vdd.n116 gnd 0.008094f
C1226 vdd.n117 gnd 0.094987f
C1227 vdd.n118 gnd 0.00499f
C1228 vdd.n119 gnd 0.004631f
C1229 vdd.n120 gnd 0.002561f
C1230 vdd.n121 gnd 0.005881f
C1231 vdd.n122 gnd 0.002488f
C1232 vdd.n123 gnd 0.002635f
C1233 vdd.n124 gnd 0.004631f
C1234 vdd.n125 gnd 0.002488f
C1235 vdd.n126 gnd 0.005881f
C1236 vdd.n127 gnd 0.002635f
C1237 vdd.n128 gnd 0.004631f
C1238 vdd.n129 gnd 0.002488f
C1239 vdd.n130 gnd 0.004411f
C1240 vdd.n131 gnd 0.004424f
C1241 vdd.t142 gnd 0.012636f
C1242 vdd.n132 gnd 0.028114f
C1243 vdd.n133 gnd 0.146311f
C1244 vdd.n134 gnd 0.002488f
C1245 vdd.n135 gnd 0.002635f
C1246 vdd.n136 gnd 0.005881f
C1247 vdd.n137 gnd 0.005881f
C1248 vdd.n138 gnd 0.002635f
C1249 vdd.n139 gnd 0.002488f
C1250 vdd.n140 gnd 0.004631f
C1251 vdd.n141 gnd 0.004631f
C1252 vdd.n142 gnd 0.002488f
C1253 vdd.n143 gnd 0.002635f
C1254 vdd.n144 gnd 0.005881f
C1255 vdd.n145 gnd 0.005881f
C1256 vdd.n146 gnd 0.002635f
C1257 vdd.n147 gnd 0.002488f
C1258 vdd.n148 gnd 0.004631f
C1259 vdd.n149 gnd 0.004631f
C1260 vdd.n150 gnd 0.002488f
C1261 vdd.n151 gnd 0.002635f
C1262 vdd.n152 gnd 0.005881f
C1263 vdd.n153 gnd 0.005881f
C1264 vdd.n154 gnd 0.013905f
C1265 vdd.n155 gnd 0.002561f
C1266 vdd.n156 gnd 0.002488f
C1267 vdd.n157 gnd 0.011968f
C1268 vdd.n158 gnd 0.008356f
C1269 vdd.t144 gnd 0.029274f
C1270 vdd.t155 gnd 0.029274f
C1271 vdd.n159 gnd 0.201188f
C1272 vdd.n160 gnd 0.158204f
C1273 vdd.t119 gnd 0.029274f
C1274 vdd.t138 gnd 0.029274f
C1275 vdd.n161 gnd 0.201188f
C1276 vdd.n162 gnd 0.127669f
C1277 vdd.t154 gnd 0.029274f
C1278 vdd.t175 gnd 0.029274f
C1279 vdd.n163 gnd 0.201188f
C1280 vdd.n164 gnd 0.127669f
C1281 vdd.n165 gnd 0.00499f
C1282 vdd.n166 gnd 0.004631f
C1283 vdd.n167 gnd 0.002561f
C1284 vdd.n168 gnd 0.005881f
C1285 vdd.n169 gnd 0.002488f
C1286 vdd.n170 gnd 0.002635f
C1287 vdd.n171 gnd 0.004631f
C1288 vdd.n172 gnd 0.002488f
C1289 vdd.n173 gnd 0.005881f
C1290 vdd.n174 gnd 0.002635f
C1291 vdd.n175 gnd 0.004631f
C1292 vdd.n176 gnd 0.002488f
C1293 vdd.n177 gnd 0.004411f
C1294 vdd.n178 gnd 0.004424f
C1295 vdd.t132 gnd 0.012636f
C1296 vdd.n179 gnd 0.028114f
C1297 vdd.n180 gnd 0.146311f
C1298 vdd.n181 gnd 0.002488f
C1299 vdd.n182 gnd 0.002635f
C1300 vdd.n183 gnd 0.005881f
C1301 vdd.n184 gnd 0.005881f
C1302 vdd.n185 gnd 0.002635f
C1303 vdd.n186 gnd 0.002488f
C1304 vdd.n187 gnd 0.004631f
C1305 vdd.n188 gnd 0.004631f
C1306 vdd.n189 gnd 0.002488f
C1307 vdd.n190 gnd 0.002635f
C1308 vdd.n191 gnd 0.005881f
C1309 vdd.n192 gnd 0.005881f
C1310 vdd.n193 gnd 0.002635f
C1311 vdd.n194 gnd 0.002488f
C1312 vdd.n195 gnd 0.004631f
C1313 vdd.n196 gnd 0.004631f
C1314 vdd.n197 gnd 0.002488f
C1315 vdd.n198 gnd 0.002635f
C1316 vdd.n199 gnd 0.005881f
C1317 vdd.n200 gnd 0.005881f
C1318 vdd.n201 gnd 0.013905f
C1319 vdd.n202 gnd 0.002561f
C1320 vdd.n203 gnd 0.002488f
C1321 vdd.n204 gnd 0.011968f
C1322 vdd.n205 gnd 0.008094f
C1323 vdd.n206 gnd 0.056507f
C1324 vdd.n207 gnd 0.203611f
C1325 vdd.n208 gnd 0.00499f
C1326 vdd.n209 gnd 0.004631f
C1327 vdd.n210 gnd 0.002561f
C1328 vdd.n211 gnd 0.005881f
C1329 vdd.n212 gnd 0.002488f
C1330 vdd.n213 gnd 0.002635f
C1331 vdd.n214 gnd 0.004631f
C1332 vdd.n215 gnd 0.002488f
C1333 vdd.n216 gnd 0.005881f
C1334 vdd.n217 gnd 0.002635f
C1335 vdd.n218 gnd 0.004631f
C1336 vdd.n219 gnd 0.002488f
C1337 vdd.n220 gnd 0.004411f
C1338 vdd.n221 gnd 0.004424f
C1339 vdd.t147 gnd 0.012636f
C1340 vdd.n222 gnd 0.028114f
C1341 vdd.n223 gnd 0.146311f
C1342 vdd.n224 gnd 0.002488f
C1343 vdd.n225 gnd 0.002635f
C1344 vdd.n226 gnd 0.005881f
C1345 vdd.n227 gnd 0.005881f
C1346 vdd.n228 gnd 0.002635f
C1347 vdd.n229 gnd 0.002488f
C1348 vdd.n230 gnd 0.004631f
C1349 vdd.n231 gnd 0.004631f
C1350 vdd.n232 gnd 0.002488f
C1351 vdd.n233 gnd 0.002635f
C1352 vdd.n234 gnd 0.005881f
C1353 vdd.n235 gnd 0.005881f
C1354 vdd.n236 gnd 0.002635f
C1355 vdd.n237 gnd 0.002488f
C1356 vdd.n238 gnd 0.004631f
C1357 vdd.n239 gnd 0.004631f
C1358 vdd.n240 gnd 0.002488f
C1359 vdd.n241 gnd 0.002635f
C1360 vdd.n242 gnd 0.005881f
C1361 vdd.n243 gnd 0.005881f
C1362 vdd.n244 gnd 0.013905f
C1363 vdd.n245 gnd 0.002561f
C1364 vdd.n246 gnd 0.002488f
C1365 vdd.n247 gnd 0.011968f
C1366 vdd.n248 gnd 0.008356f
C1367 vdd.t148 gnd 0.029274f
C1368 vdd.t164 gnd 0.029274f
C1369 vdd.n249 gnd 0.201188f
C1370 vdd.n250 gnd 0.158204f
C1371 vdd.t125 gnd 0.029274f
C1372 vdd.t146 gnd 0.029274f
C1373 vdd.n251 gnd 0.201188f
C1374 vdd.n252 gnd 0.127669f
C1375 vdd.t159 gnd 0.029274f
C1376 vdd.t123 gnd 0.029274f
C1377 vdd.n253 gnd 0.201188f
C1378 vdd.n254 gnd 0.127669f
C1379 vdd.n255 gnd 0.00499f
C1380 vdd.n256 gnd 0.004631f
C1381 vdd.n257 gnd 0.002561f
C1382 vdd.n258 gnd 0.005881f
C1383 vdd.n259 gnd 0.002488f
C1384 vdd.n260 gnd 0.002635f
C1385 vdd.n261 gnd 0.004631f
C1386 vdd.n262 gnd 0.002488f
C1387 vdd.n263 gnd 0.005881f
C1388 vdd.n264 gnd 0.002635f
C1389 vdd.n265 gnd 0.004631f
C1390 vdd.n266 gnd 0.002488f
C1391 vdd.n267 gnd 0.004411f
C1392 vdd.n268 gnd 0.004424f
C1393 vdd.t136 gnd 0.012636f
C1394 vdd.n269 gnd 0.028114f
C1395 vdd.n270 gnd 0.146311f
C1396 vdd.n271 gnd 0.002488f
C1397 vdd.n272 gnd 0.002635f
C1398 vdd.n273 gnd 0.005881f
C1399 vdd.n274 gnd 0.005881f
C1400 vdd.n275 gnd 0.002635f
C1401 vdd.n276 gnd 0.002488f
C1402 vdd.n277 gnd 0.004631f
C1403 vdd.n278 gnd 0.004631f
C1404 vdd.n279 gnd 0.002488f
C1405 vdd.n280 gnd 0.002635f
C1406 vdd.n281 gnd 0.005881f
C1407 vdd.n282 gnd 0.005881f
C1408 vdd.n283 gnd 0.002635f
C1409 vdd.n284 gnd 0.002488f
C1410 vdd.n285 gnd 0.004631f
C1411 vdd.n286 gnd 0.004631f
C1412 vdd.n287 gnd 0.002488f
C1413 vdd.n288 gnd 0.002635f
C1414 vdd.n289 gnd 0.005881f
C1415 vdd.n290 gnd 0.005881f
C1416 vdd.n291 gnd 0.013905f
C1417 vdd.n292 gnd 0.002561f
C1418 vdd.n293 gnd 0.002488f
C1419 vdd.n294 gnd 0.011968f
C1420 vdd.n295 gnd 0.008094f
C1421 vdd.n296 gnd 0.056507f
C1422 vdd.n297 gnd 0.220385f
C1423 vdd.n298 gnd 0.006988f
C1424 vdd.n299 gnd 0.009093f
C1425 vdd.n300 gnd 0.007318f
C1426 vdd.n301 gnd 0.007318f
C1427 vdd.n302 gnd 0.009093f
C1428 vdd.n303 gnd 0.009093f
C1429 vdd.n304 gnd 0.664388f
C1430 vdd.n305 gnd 0.009093f
C1431 vdd.n306 gnd 0.009093f
C1432 vdd.n307 gnd 0.009093f
C1433 vdd.n308 gnd 0.720141f
C1434 vdd.n309 gnd 0.009093f
C1435 vdd.n310 gnd 0.009093f
C1436 vdd.n311 gnd 0.009093f
C1437 vdd.n312 gnd 0.009093f
C1438 vdd.n313 gnd 0.007318f
C1439 vdd.n314 gnd 0.009093f
C1440 vdd.t122 gnd 0.464607f
C1441 vdd.n315 gnd 0.009093f
C1442 vdd.n316 gnd 0.009093f
C1443 vdd.n317 gnd 0.009093f
C1444 vdd.n318 gnd 0.929214f
C1445 vdd.n319 gnd 0.009093f
C1446 vdd.n320 gnd 0.009093f
C1447 vdd.n321 gnd 0.009093f
C1448 vdd.n322 gnd 0.009093f
C1449 vdd.n323 gnd 0.009093f
C1450 vdd.n324 gnd 0.007318f
C1451 vdd.n325 gnd 0.009093f
C1452 vdd.n326 gnd 0.009093f
C1453 vdd.n327 gnd 0.009093f
C1454 vdd.n328 gnd 0.022159f
C1455 vdd.n329 gnd 2.22082f
C1456 vdd.n330 gnd 0.022667f
C1457 vdd.n331 gnd 0.009093f
C1458 vdd.n332 gnd 0.009093f
C1459 vdd.n334 gnd 0.009093f
C1460 vdd.n335 gnd 0.009093f
C1461 vdd.n336 gnd 0.007318f
C1462 vdd.n337 gnd 0.007318f
C1463 vdd.n338 gnd 0.009093f
C1464 vdd.n339 gnd 0.009093f
C1465 vdd.n340 gnd 0.009093f
C1466 vdd.n341 gnd 0.009093f
C1467 vdd.n342 gnd 0.009093f
C1468 vdd.n343 gnd 0.009093f
C1469 vdd.n344 gnd 0.007318f
C1470 vdd.n346 gnd 0.009093f
C1471 vdd.n347 gnd 0.009093f
C1472 vdd.n348 gnd 0.009093f
C1473 vdd.n349 gnd 0.009093f
C1474 vdd.n350 gnd 0.009093f
C1475 vdd.n351 gnd 0.007318f
C1476 vdd.n353 gnd 0.009093f
C1477 vdd.n354 gnd 0.009093f
C1478 vdd.n355 gnd 0.009093f
C1479 vdd.n356 gnd 0.009093f
C1480 vdd.n357 gnd 0.009093f
C1481 vdd.n358 gnd 0.007318f
C1482 vdd.n360 gnd 0.009093f
C1483 vdd.n361 gnd 0.009093f
C1484 vdd.n362 gnd 0.009093f
C1485 vdd.n363 gnd 0.009093f
C1486 vdd.n364 gnd 0.006111f
C1487 vdd.t45 gnd 0.111862f
C1488 vdd.t44 gnd 0.11955f
C1489 vdd.t43 gnd 0.14609f
C1490 vdd.n365 gnd 0.187267f
C1491 vdd.n366 gnd 0.15807f
C1492 vdd.n368 gnd 0.009093f
C1493 vdd.n369 gnd 0.009093f
C1494 vdd.n370 gnd 0.007318f
C1495 vdd.n371 gnd 0.009093f
C1496 vdd.n373 gnd 0.009093f
C1497 vdd.n374 gnd 0.009093f
C1498 vdd.n375 gnd 0.009093f
C1499 vdd.n376 gnd 0.009093f
C1500 vdd.n377 gnd 0.007318f
C1501 vdd.n379 gnd 0.009093f
C1502 vdd.n380 gnd 0.009093f
C1503 vdd.n381 gnd 0.009093f
C1504 vdd.n382 gnd 0.009093f
C1505 vdd.n383 gnd 0.009093f
C1506 vdd.n384 gnd 0.007318f
C1507 vdd.n386 gnd 0.009093f
C1508 vdd.n387 gnd 0.009093f
C1509 vdd.n388 gnd 0.009093f
C1510 vdd.n389 gnd 0.009093f
C1511 vdd.n390 gnd 0.009093f
C1512 vdd.n391 gnd 0.007318f
C1513 vdd.n393 gnd 0.009093f
C1514 vdd.n394 gnd 0.009093f
C1515 vdd.n395 gnd 0.009093f
C1516 vdd.n396 gnd 0.009093f
C1517 vdd.n397 gnd 0.009093f
C1518 vdd.n398 gnd 0.007318f
C1519 vdd.n400 gnd 0.009093f
C1520 vdd.n401 gnd 0.009093f
C1521 vdd.n402 gnd 0.009093f
C1522 vdd.n403 gnd 0.009093f
C1523 vdd.n404 gnd 0.007245f
C1524 vdd.t39 gnd 0.111862f
C1525 vdd.t38 gnd 0.11955f
C1526 vdd.t36 gnd 0.14609f
C1527 vdd.n405 gnd 0.187267f
C1528 vdd.n406 gnd 0.15807f
C1529 vdd.n408 gnd 0.009093f
C1530 vdd.n409 gnd 0.009093f
C1531 vdd.n410 gnd 0.007318f
C1532 vdd.n411 gnd 0.009093f
C1533 vdd.n413 gnd 0.009093f
C1534 vdd.n414 gnd 0.009093f
C1535 vdd.n415 gnd 0.009093f
C1536 vdd.n416 gnd 0.009093f
C1537 vdd.n417 gnd 0.007318f
C1538 vdd.n419 gnd 0.009093f
C1539 vdd.n420 gnd 0.009093f
C1540 vdd.n421 gnd 0.009093f
C1541 vdd.n422 gnd 0.009093f
C1542 vdd.n423 gnd 0.009093f
C1543 vdd.n424 gnd 0.007318f
C1544 vdd.n426 gnd 0.009093f
C1545 vdd.n427 gnd 0.009093f
C1546 vdd.n428 gnd 0.009093f
C1547 vdd.n429 gnd 0.009093f
C1548 vdd.n430 gnd 0.009093f
C1549 vdd.n431 gnd 0.007318f
C1550 vdd.n433 gnd 0.009093f
C1551 vdd.n434 gnd 0.009093f
C1552 vdd.n435 gnd 0.009093f
C1553 vdd.n436 gnd 0.009093f
C1554 vdd.n437 gnd 0.009093f
C1555 vdd.n438 gnd 0.007318f
C1556 vdd.n440 gnd 0.009093f
C1557 vdd.n441 gnd 0.009093f
C1558 vdd.n442 gnd 0.009093f
C1559 vdd.n443 gnd 0.009093f
C1560 vdd.n444 gnd 0.009093f
C1561 vdd.n445 gnd 0.009093f
C1562 vdd.n446 gnd 0.007318f
C1563 vdd.n447 gnd 0.009093f
C1564 vdd.n448 gnd 0.009093f
C1565 vdd.n449 gnd 0.007318f
C1566 vdd.n450 gnd 0.009093f
C1567 vdd.n451 gnd 0.007318f
C1568 vdd.n452 gnd 0.009093f
C1569 vdd.n453 gnd 0.007318f
C1570 vdd.n454 gnd 0.009093f
C1571 vdd.n455 gnd 0.009093f
C1572 vdd.n456 gnd 0.506422f
C1573 vdd.t118 gnd 0.464607f
C1574 vdd.n457 gnd 0.009093f
C1575 vdd.n458 gnd 0.007318f
C1576 vdd.n459 gnd 0.009093f
C1577 vdd.n460 gnd 0.007318f
C1578 vdd.n461 gnd 0.009093f
C1579 vdd.t143 gnd 0.464607f
C1580 vdd.n462 gnd 0.009093f
C1581 vdd.n463 gnd 0.007318f
C1582 vdd.n464 gnd 0.009093f
C1583 vdd.n465 gnd 0.007318f
C1584 vdd.n466 gnd 0.009093f
C1585 vdd.t114 gnd 0.464607f
C1586 vdd.n467 gnd 0.580759f
C1587 vdd.n468 gnd 0.009093f
C1588 vdd.n469 gnd 0.007318f
C1589 vdd.n470 gnd 0.009093f
C1590 vdd.n471 gnd 0.007318f
C1591 vdd.n472 gnd 0.009093f
C1592 vdd.n473 gnd 0.929214f
C1593 vdd.n474 gnd 0.009093f
C1594 vdd.n475 gnd 0.007318f
C1595 vdd.n476 gnd 0.022159f
C1596 vdd.n477 gnd 0.006074f
C1597 vdd.n478 gnd 0.022159f
C1598 vdd.t15 gnd 0.464607f
C1599 vdd.n479 gnd 0.022159f
C1600 vdd.n480 gnd 0.006074f
C1601 vdd.n481 gnd 0.00782f
C1602 vdd.n482 gnd 0.007318f
C1603 vdd.n483 gnd 0.009093f
C1604 vdd.n484 gnd 6.40228f
C1605 vdd.n515 gnd 0.022667f
C1606 vdd.n516 gnd 1.27767f
C1607 vdd.n517 gnd 0.009093f
C1608 vdd.n518 gnd 0.007318f
C1609 vdd.n519 gnd 0.005819f
C1610 vdd.n520 gnd 0.014858f
C1611 vdd.n521 gnd 0.007318f
C1612 vdd.n522 gnd 0.009093f
C1613 vdd.n523 gnd 0.009093f
C1614 vdd.n524 gnd 0.009093f
C1615 vdd.n525 gnd 0.009093f
C1616 vdd.n526 gnd 0.009093f
C1617 vdd.n527 gnd 0.009093f
C1618 vdd.n528 gnd 0.009093f
C1619 vdd.n529 gnd 0.009093f
C1620 vdd.n530 gnd 0.009093f
C1621 vdd.n531 gnd 0.009093f
C1622 vdd.n532 gnd 0.009093f
C1623 vdd.n533 gnd 0.009093f
C1624 vdd.n534 gnd 0.009093f
C1625 vdd.n535 gnd 0.009093f
C1626 vdd.n536 gnd 0.006111f
C1627 vdd.n537 gnd 0.009093f
C1628 vdd.n538 gnd 0.009093f
C1629 vdd.n539 gnd 0.009093f
C1630 vdd.n540 gnd 0.009093f
C1631 vdd.n541 gnd 0.009093f
C1632 vdd.n542 gnd 0.009093f
C1633 vdd.n543 gnd 0.009093f
C1634 vdd.n544 gnd 0.009093f
C1635 vdd.n545 gnd 0.009093f
C1636 vdd.n546 gnd 0.009093f
C1637 vdd.n547 gnd 0.009093f
C1638 vdd.n548 gnd 0.009093f
C1639 vdd.n549 gnd 0.009093f
C1640 vdd.n550 gnd 0.009093f
C1641 vdd.n551 gnd 0.009093f
C1642 vdd.n552 gnd 0.009093f
C1643 vdd.n553 gnd 0.009093f
C1644 vdd.n554 gnd 0.009093f
C1645 vdd.n555 gnd 0.009093f
C1646 vdd.n556 gnd 0.007245f
C1647 vdd.t16 gnd 0.111862f
C1648 vdd.t17 gnd 0.11955f
C1649 vdd.t14 gnd 0.14609f
C1650 vdd.n557 gnd 0.187267f
C1651 vdd.n558 gnd 0.157338f
C1652 vdd.n559 gnd 0.009093f
C1653 vdd.n560 gnd 0.009093f
C1654 vdd.n561 gnd 0.009093f
C1655 vdd.n562 gnd 0.009093f
C1656 vdd.n563 gnd 0.009093f
C1657 vdd.n564 gnd 0.009093f
C1658 vdd.n565 gnd 0.009093f
C1659 vdd.n566 gnd 0.009093f
C1660 vdd.n567 gnd 0.009093f
C1661 vdd.n568 gnd 0.009093f
C1662 vdd.n569 gnd 0.009093f
C1663 vdd.n570 gnd 0.009093f
C1664 vdd.n571 gnd 0.009093f
C1665 vdd.n572 gnd 0.005819f
C1666 vdd.n575 gnd 0.006183f
C1667 vdd.n576 gnd 0.006183f
C1668 vdd.n577 gnd 0.006183f
C1669 vdd.n578 gnd 0.006183f
C1670 vdd.n579 gnd 0.006183f
C1671 vdd.n580 gnd 0.006183f
C1672 vdd.n582 gnd 0.006183f
C1673 vdd.n583 gnd 0.006183f
C1674 vdd.n585 gnd 0.006183f
C1675 vdd.n586 gnd 0.004501f
C1676 vdd.n588 gnd 0.006183f
C1677 vdd.t60 gnd 0.249851f
C1678 vdd.t59 gnd 0.255754f
C1679 vdd.t58 gnd 0.163112f
C1680 vdd.n589 gnd 0.088153f
C1681 vdd.n590 gnd 0.050003f
C1682 vdd.n591 gnd 0.008836f
C1683 vdd.n592 gnd 0.014451f
C1684 vdd.n594 gnd 0.006183f
C1685 vdd.n595 gnd 0.631866f
C1686 vdd.n596 gnd 0.013698f
C1687 vdd.n597 gnd 0.013698f
C1688 vdd.n598 gnd 0.006183f
C1689 vdd.n599 gnd 0.014671f
C1690 vdd.n600 gnd 0.006183f
C1691 vdd.n601 gnd 0.006183f
C1692 vdd.n602 gnd 0.006183f
C1693 vdd.n603 gnd 0.006183f
C1694 vdd.n604 gnd 0.006183f
C1695 vdd.n606 gnd 0.006183f
C1696 vdd.n607 gnd 0.006183f
C1697 vdd.n609 gnd 0.006183f
C1698 vdd.n610 gnd 0.006183f
C1699 vdd.n612 gnd 0.006183f
C1700 vdd.n613 gnd 0.006183f
C1701 vdd.n615 gnd 0.006183f
C1702 vdd.n616 gnd 0.006183f
C1703 vdd.n618 gnd 0.006183f
C1704 vdd.n619 gnd 0.006183f
C1705 vdd.n621 gnd 0.006183f
C1706 vdd.t53 gnd 0.249851f
C1707 vdd.t52 gnd 0.255754f
C1708 vdd.t50 gnd 0.163112f
C1709 vdd.n622 gnd 0.088153f
C1710 vdd.n623 gnd 0.050003f
C1711 vdd.n624 gnd 0.006183f
C1712 vdd.n626 gnd 0.006183f
C1713 vdd.n627 gnd 0.006183f
C1714 vdd.t51 gnd 0.315933f
C1715 vdd.n628 gnd 0.006183f
C1716 vdd.n629 gnd 0.006183f
C1717 vdd.n630 gnd 0.006183f
C1718 vdd.n631 gnd 0.006183f
C1719 vdd.n632 gnd 0.006183f
C1720 vdd.n633 gnd 0.631866f
C1721 vdd.n634 gnd 0.006183f
C1722 vdd.n635 gnd 0.006183f
C1723 vdd.n636 gnd 0.552882f
C1724 vdd.n637 gnd 0.006183f
C1725 vdd.n638 gnd 0.006183f
C1726 vdd.n639 gnd 0.005456f
C1727 vdd.n640 gnd 0.006183f
C1728 vdd.n641 gnd 0.557528f
C1729 vdd.n642 gnd 0.006183f
C1730 vdd.n643 gnd 0.006183f
C1731 vdd.n644 gnd 0.006183f
C1732 vdd.n645 gnd 0.006183f
C1733 vdd.n646 gnd 0.006183f
C1734 vdd.n647 gnd 0.631866f
C1735 vdd.n648 gnd 0.006183f
C1736 vdd.n649 gnd 0.006183f
C1737 vdd.t30 gnd 0.28341f
C1738 vdd.t100 gnd 0.074337f
C1739 vdd.n650 gnd 0.006183f
C1740 vdd.n651 gnd 0.006183f
C1741 vdd.n652 gnd 0.006183f
C1742 vdd.t103 gnd 0.315933f
C1743 vdd.n653 gnd 0.006183f
C1744 vdd.n654 gnd 0.006183f
C1745 vdd.n655 gnd 0.006183f
C1746 vdd.n656 gnd 0.006183f
C1747 vdd.n657 gnd 0.006183f
C1748 vdd.t90 gnd 0.315933f
C1749 vdd.n658 gnd 0.006183f
C1750 vdd.n659 gnd 0.006183f
C1751 vdd.n660 gnd 0.525006f
C1752 vdd.n661 gnd 0.006183f
C1753 vdd.n662 gnd 0.006183f
C1754 vdd.n663 gnd 0.006183f
C1755 vdd.n664 gnd 0.385624f
C1756 vdd.n665 gnd 0.006183f
C1757 vdd.n666 gnd 0.006183f
C1758 vdd.t107 gnd 0.315933f
C1759 vdd.n667 gnd 0.006183f
C1760 vdd.n668 gnd 0.006183f
C1761 vdd.n669 gnd 0.006183f
C1762 vdd.n670 gnd 0.525006f
C1763 vdd.n671 gnd 0.006183f
C1764 vdd.n672 gnd 0.006183f
C1765 vdd.t111 gnd 0.269472f
C1766 vdd.t95 gnd 0.246242f
C1767 vdd.n673 gnd 0.006183f
C1768 vdd.n674 gnd 0.006183f
C1769 vdd.n675 gnd 0.006183f
C1770 vdd.t196 gnd 0.315933f
C1771 vdd.n676 gnd 0.006183f
C1772 vdd.n677 gnd 0.006183f
C1773 vdd.t10 gnd 0.315933f
C1774 vdd.n678 gnd 0.006183f
C1775 vdd.n679 gnd 0.006183f
C1776 vdd.n680 gnd 0.006183f
C1777 vdd.t13 gnd 0.232304f
C1778 vdd.n681 gnd 0.006183f
C1779 vdd.n682 gnd 0.006183f
C1780 vdd.n683 gnd 0.538944f
C1781 vdd.n684 gnd 0.006183f
C1782 vdd.n685 gnd 0.006183f
C1783 vdd.n686 gnd 0.006183f
C1784 vdd.n687 gnd 0.631866f
C1785 vdd.n688 gnd 0.006183f
C1786 vdd.n689 gnd 0.006183f
C1787 vdd.t0 gnd 0.28341f
C1788 vdd.n690 gnd 0.399562f
C1789 vdd.n691 gnd 0.006183f
C1790 vdd.n692 gnd 0.006183f
C1791 vdd.n693 gnd 0.006183f
C1792 vdd.t11 gnd 0.315933f
C1793 vdd.n694 gnd 0.006183f
C1794 vdd.n695 gnd 0.006183f
C1795 vdd.n696 gnd 0.006183f
C1796 vdd.n697 gnd 0.006183f
C1797 vdd.n698 gnd 0.006183f
C1798 vdd.t3 gnd 0.631866f
C1799 vdd.n699 gnd 0.006183f
C1800 vdd.n700 gnd 0.006183f
C1801 vdd.t55 gnd 0.315933f
C1802 vdd.n701 gnd 0.006183f
C1803 vdd.n702 gnd 0.014671f
C1804 vdd.n703 gnd 0.014671f
C1805 vdd.t5 gnd 0.594697f
C1806 vdd.n704 gnd 0.013698f
C1807 vdd.n705 gnd 0.013698f
C1808 vdd.n706 gnd 0.014671f
C1809 vdd.n707 gnd 0.006183f
C1810 vdd.n708 gnd 0.006183f
C1811 vdd.t194 gnd 0.594697f
C1812 vdd.n726 gnd 0.014671f
C1813 vdd.n744 gnd 0.013698f
C1814 vdd.n745 gnd 0.006183f
C1815 vdd.n746 gnd 0.013698f
C1816 vdd.t80 gnd 0.249851f
C1817 vdd.t79 gnd 0.255754f
C1818 vdd.t78 gnd 0.163112f
C1819 vdd.n747 gnd 0.088153f
C1820 vdd.n748 gnd 0.050003f
C1821 vdd.n749 gnd 0.014451f
C1822 vdd.n750 gnd 0.006183f
C1823 vdd.t91 gnd 0.631866f
C1824 vdd.n751 gnd 0.013698f
C1825 vdd.n752 gnd 0.006183f
C1826 vdd.n753 gnd 0.014671f
C1827 vdd.n754 gnd 0.006183f
C1828 vdd.t49 gnd 0.249851f
C1829 vdd.t48 gnd 0.255754f
C1830 vdd.t46 gnd 0.163112f
C1831 vdd.n755 gnd 0.088153f
C1832 vdd.n756 gnd 0.050003f
C1833 vdd.n757 gnd 0.008836f
C1834 vdd.n758 gnd 0.006183f
C1835 vdd.n759 gnd 0.006183f
C1836 vdd.t47 gnd 0.315933f
C1837 vdd.n760 gnd 0.006183f
C1838 vdd.n761 gnd 0.006183f
C1839 vdd.n762 gnd 0.006183f
C1840 vdd.n763 gnd 0.006183f
C1841 vdd.n764 gnd 0.006183f
C1842 vdd.n765 gnd 0.006183f
C1843 vdd.n766 gnd 0.631866f
C1844 vdd.n767 gnd 0.006183f
C1845 vdd.n768 gnd 0.006183f
C1846 vdd.t105 gnd 0.315933f
C1847 vdd.n769 gnd 0.006183f
C1848 vdd.n770 gnd 0.006183f
C1849 vdd.n771 gnd 0.006183f
C1850 vdd.n772 gnd 0.006183f
C1851 vdd.n773 gnd 0.399562f
C1852 vdd.n774 gnd 0.006183f
C1853 vdd.n775 gnd 0.006183f
C1854 vdd.n776 gnd 0.006183f
C1855 vdd.n777 gnd 0.006183f
C1856 vdd.n778 gnd 0.006183f
C1857 vdd.n779 gnd 0.538944f
C1858 vdd.n780 gnd 0.006183f
C1859 vdd.n781 gnd 0.006183f
C1860 vdd.t198 gnd 0.28341f
C1861 vdd.t110 gnd 0.232304f
C1862 vdd.n782 gnd 0.006183f
C1863 vdd.n783 gnd 0.006183f
C1864 vdd.n784 gnd 0.006183f
C1865 vdd.t2 gnd 0.315933f
C1866 vdd.n785 gnd 0.006183f
C1867 vdd.n786 gnd 0.006183f
C1868 vdd.t93 gnd 0.315933f
C1869 vdd.n787 gnd 0.006183f
C1870 vdd.n788 gnd 0.006183f
C1871 vdd.n789 gnd 0.006183f
C1872 vdd.t101 gnd 0.246242f
C1873 vdd.n790 gnd 0.006183f
C1874 vdd.n791 gnd 0.006183f
C1875 vdd.n792 gnd 0.525006f
C1876 vdd.n793 gnd 0.006183f
C1877 vdd.n794 gnd 0.006183f
C1878 vdd.n795 gnd 0.006183f
C1879 vdd.t8 gnd 0.315933f
C1880 vdd.n796 gnd 0.006183f
C1881 vdd.n797 gnd 0.006183f
C1882 vdd.t7 gnd 0.269472f
C1883 vdd.n798 gnd 0.385624f
C1884 vdd.n799 gnd 0.006183f
C1885 vdd.n800 gnd 0.006183f
C1886 vdd.n801 gnd 0.006183f
C1887 vdd.n802 gnd 0.525006f
C1888 vdd.n803 gnd 0.006183f
C1889 vdd.n804 gnd 0.006183f
C1890 vdd.t109 gnd 0.315933f
C1891 vdd.n805 gnd 0.006183f
C1892 vdd.n806 gnd 0.006183f
C1893 vdd.n807 gnd 0.006183f
C1894 vdd.n808 gnd 0.631866f
C1895 vdd.n809 gnd 0.006183f
C1896 vdd.n810 gnd 0.006183f
C1897 vdd.t104 gnd 0.315933f
C1898 vdd.n811 gnd 0.006183f
C1899 vdd.n812 gnd 0.006183f
C1900 vdd.n813 gnd 0.006183f
C1901 vdd.t97 gnd 0.074337f
C1902 vdd.n814 gnd 0.006183f
C1903 vdd.n815 gnd 0.006183f
C1904 vdd.n816 gnd 0.006183f
C1905 vdd.t67 gnd 0.255754f
C1906 vdd.t65 gnd 0.163112f
C1907 vdd.t68 gnd 0.255754f
C1908 vdd.n817 gnd 0.143744f
C1909 vdd.n818 gnd 0.006183f
C1910 vdd.n819 gnd 0.006183f
C1911 vdd.n820 gnd 0.631866f
C1912 vdd.n821 gnd 0.006183f
C1913 vdd.n822 gnd 0.006183f
C1914 vdd.t66 gnd 0.28341f
C1915 vdd.n823 gnd 0.557528f
C1916 vdd.n824 gnd 0.006183f
C1917 vdd.n825 gnd 0.006183f
C1918 vdd.n826 gnd 0.006183f
C1919 vdd.n827 gnd 0.552882f
C1920 vdd.n828 gnd 0.006183f
C1921 vdd.n829 gnd 0.006183f
C1922 vdd.n830 gnd 0.006183f
C1923 vdd.n831 gnd 0.006183f
C1924 vdd.n832 gnd 0.006183f
C1925 vdd.n833 gnd 0.631866f
C1926 vdd.n834 gnd 0.006183f
C1927 vdd.n835 gnd 0.006183f
C1928 vdd.t62 gnd 0.315933f
C1929 vdd.n836 gnd 0.006183f
C1930 vdd.n837 gnd 0.014671f
C1931 vdd.n838 gnd 0.014671f
C1932 vdd.n839 gnd 6.40228f
C1933 vdd.n840 gnd 0.013698f
C1934 vdd.n841 gnd 0.013698f
C1935 vdd.n842 gnd 0.014671f
C1936 vdd.n843 gnd 0.006183f
C1937 vdd.n844 gnd 0.006183f
C1938 vdd.n845 gnd 0.006183f
C1939 vdd.n846 gnd 0.006183f
C1940 vdd.n847 gnd 0.006183f
C1941 vdd.n848 gnd 0.006183f
C1942 vdd.n849 gnd 0.006183f
C1943 vdd.n850 gnd 0.006183f
C1944 vdd.n852 gnd 0.006183f
C1945 vdd.n853 gnd 0.006183f
C1946 vdd.n854 gnd 0.005819f
C1947 vdd.n857 gnd 0.022667f
C1948 vdd.n858 gnd 0.007318f
C1949 vdd.n859 gnd 0.009093f
C1950 vdd.n861 gnd 0.009093f
C1951 vdd.n862 gnd 0.006074f
C1952 vdd.t22 gnd 0.464607f
C1953 vdd.n863 gnd 6.7368f
C1954 vdd.n864 gnd 0.009093f
C1955 vdd.n865 gnd 0.022667f
C1956 vdd.n866 gnd 0.007318f
C1957 vdd.n867 gnd 0.009093f
C1958 vdd.n868 gnd 0.007318f
C1959 vdd.n869 gnd 0.009093f
C1960 vdd.n870 gnd 0.929214f
C1961 vdd.n871 gnd 0.009093f
C1962 vdd.n872 gnd 0.007318f
C1963 vdd.n873 gnd 0.007318f
C1964 vdd.n874 gnd 0.009093f
C1965 vdd.n875 gnd 0.007318f
C1966 vdd.n876 gnd 0.009093f
C1967 vdd.t112 gnd 0.464607f
C1968 vdd.n877 gnd 0.009093f
C1969 vdd.n878 gnd 0.007318f
C1970 vdd.n879 gnd 0.009093f
C1971 vdd.n880 gnd 0.007318f
C1972 vdd.n881 gnd 0.009093f
C1973 vdd.t165 gnd 0.464607f
C1974 vdd.n882 gnd 0.009093f
C1975 vdd.n883 gnd 0.007318f
C1976 vdd.n884 gnd 0.009093f
C1977 vdd.n885 gnd 0.007318f
C1978 vdd.n886 gnd 0.009093f
C1979 vdd.n887 gnd 0.729433f
C1980 vdd.n888 gnd 0.771248f
C1981 vdd.t120 gnd 0.464607f
C1982 vdd.n889 gnd 0.009093f
C1983 vdd.n890 gnd 0.007318f
C1984 vdd.n891 gnd 0.00499f
C1985 vdd.n892 gnd 0.004631f
C1986 vdd.n893 gnd 0.002561f
C1987 vdd.n894 gnd 0.005881f
C1988 vdd.n895 gnd 0.002488f
C1989 vdd.n896 gnd 0.002635f
C1990 vdd.n897 gnd 0.004631f
C1991 vdd.n898 gnd 0.002488f
C1992 vdd.n899 gnd 0.005881f
C1993 vdd.n900 gnd 0.002635f
C1994 vdd.n901 gnd 0.004631f
C1995 vdd.n902 gnd 0.002488f
C1996 vdd.n903 gnd 0.004411f
C1997 vdd.n904 gnd 0.004424f
C1998 vdd.t113 gnd 0.012636f
C1999 vdd.n905 gnd 0.028114f
C2000 vdd.n906 gnd 0.146311f
C2001 vdd.n907 gnd 0.002488f
C2002 vdd.n908 gnd 0.002635f
C2003 vdd.n909 gnd 0.005881f
C2004 vdd.n910 gnd 0.005881f
C2005 vdd.n911 gnd 0.002635f
C2006 vdd.n912 gnd 0.002488f
C2007 vdd.n913 gnd 0.004631f
C2008 vdd.n914 gnd 0.004631f
C2009 vdd.n915 gnd 0.002488f
C2010 vdd.n916 gnd 0.002635f
C2011 vdd.n917 gnd 0.005881f
C2012 vdd.n918 gnd 0.005881f
C2013 vdd.n919 gnd 0.002635f
C2014 vdd.n920 gnd 0.002488f
C2015 vdd.n921 gnd 0.004631f
C2016 vdd.n922 gnd 0.004631f
C2017 vdd.n923 gnd 0.002488f
C2018 vdd.n924 gnd 0.002635f
C2019 vdd.n925 gnd 0.005881f
C2020 vdd.n926 gnd 0.005881f
C2021 vdd.n927 gnd 0.013905f
C2022 vdd.n928 gnd 0.002561f
C2023 vdd.n929 gnd 0.002488f
C2024 vdd.n930 gnd 0.011968f
C2025 vdd.n931 gnd 0.008356f
C2026 vdd.t139 gnd 0.029274f
C2027 vdd.t168 gnd 0.029274f
C2028 vdd.n932 gnd 0.201188f
C2029 vdd.n933 gnd 0.158204f
C2030 vdd.t128 gnd 0.029274f
C2031 vdd.t156 gnd 0.029274f
C2032 vdd.n934 gnd 0.201188f
C2033 vdd.n935 gnd 0.127669f
C2034 vdd.t134 gnd 0.029274f
C2035 vdd.t162 gnd 0.029274f
C2036 vdd.n936 gnd 0.201188f
C2037 vdd.n937 gnd 0.127669f
C2038 vdd.n938 gnd 0.00499f
C2039 vdd.n939 gnd 0.004631f
C2040 vdd.n940 gnd 0.002561f
C2041 vdd.n941 gnd 0.005881f
C2042 vdd.n942 gnd 0.002488f
C2043 vdd.n943 gnd 0.002635f
C2044 vdd.n944 gnd 0.004631f
C2045 vdd.n945 gnd 0.002488f
C2046 vdd.n946 gnd 0.005881f
C2047 vdd.n947 gnd 0.002635f
C2048 vdd.n948 gnd 0.004631f
C2049 vdd.n949 gnd 0.002488f
C2050 vdd.n950 gnd 0.004411f
C2051 vdd.n951 gnd 0.004424f
C2052 vdd.t172 gnd 0.012636f
C2053 vdd.n952 gnd 0.028114f
C2054 vdd.n953 gnd 0.146311f
C2055 vdd.n954 gnd 0.002488f
C2056 vdd.n955 gnd 0.002635f
C2057 vdd.n956 gnd 0.005881f
C2058 vdd.n957 gnd 0.005881f
C2059 vdd.n958 gnd 0.002635f
C2060 vdd.n959 gnd 0.002488f
C2061 vdd.n960 gnd 0.004631f
C2062 vdd.n961 gnd 0.004631f
C2063 vdd.n962 gnd 0.002488f
C2064 vdd.n963 gnd 0.002635f
C2065 vdd.n964 gnd 0.005881f
C2066 vdd.n965 gnd 0.005881f
C2067 vdd.n966 gnd 0.002635f
C2068 vdd.n967 gnd 0.002488f
C2069 vdd.n968 gnd 0.004631f
C2070 vdd.n969 gnd 0.004631f
C2071 vdd.n970 gnd 0.002488f
C2072 vdd.n971 gnd 0.002635f
C2073 vdd.n972 gnd 0.005881f
C2074 vdd.n973 gnd 0.005881f
C2075 vdd.n974 gnd 0.013905f
C2076 vdd.n975 gnd 0.002561f
C2077 vdd.n976 gnd 0.002488f
C2078 vdd.n977 gnd 0.011968f
C2079 vdd.n978 gnd 0.008094f
C2080 vdd.n979 gnd 0.094987f
C2081 vdd.n980 gnd 0.00499f
C2082 vdd.n981 gnd 0.004631f
C2083 vdd.n982 gnd 0.002561f
C2084 vdd.n983 gnd 0.005881f
C2085 vdd.n984 gnd 0.002488f
C2086 vdd.n985 gnd 0.002635f
C2087 vdd.n986 gnd 0.004631f
C2088 vdd.n987 gnd 0.002488f
C2089 vdd.n988 gnd 0.005881f
C2090 vdd.n989 gnd 0.002635f
C2091 vdd.n990 gnd 0.004631f
C2092 vdd.n991 gnd 0.002488f
C2093 vdd.n992 gnd 0.004411f
C2094 vdd.n993 gnd 0.004424f
C2095 vdd.t163 gnd 0.012636f
C2096 vdd.n994 gnd 0.028114f
C2097 vdd.n995 gnd 0.146311f
C2098 vdd.n996 gnd 0.002488f
C2099 vdd.n997 gnd 0.002635f
C2100 vdd.n998 gnd 0.005881f
C2101 vdd.n999 gnd 0.005881f
C2102 vdd.n1000 gnd 0.002635f
C2103 vdd.n1001 gnd 0.002488f
C2104 vdd.n1002 gnd 0.004631f
C2105 vdd.n1003 gnd 0.004631f
C2106 vdd.n1004 gnd 0.002488f
C2107 vdd.n1005 gnd 0.002635f
C2108 vdd.n1006 gnd 0.005881f
C2109 vdd.n1007 gnd 0.005881f
C2110 vdd.n1008 gnd 0.002635f
C2111 vdd.n1009 gnd 0.002488f
C2112 vdd.n1010 gnd 0.004631f
C2113 vdd.n1011 gnd 0.004631f
C2114 vdd.n1012 gnd 0.002488f
C2115 vdd.n1013 gnd 0.002635f
C2116 vdd.n1014 gnd 0.005881f
C2117 vdd.n1015 gnd 0.005881f
C2118 vdd.n1016 gnd 0.013905f
C2119 vdd.n1017 gnd 0.002561f
C2120 vdd.n1018 gnd 0.002488f
C2121 vdd.n1019 gnd 0.011968f
C2122 vdd.n1020 gnd 0.008356f
C2123 vdd.t121 gnd 0.029274f
C2124 vdd.t166 gnd 0.029274f
C2125 vdd.n1021 gnd 0.201188f
C2126 vdd.n1022 gnd 0.158204f
C2127 vdd.t161 gnd 0.029274f
C2128 vdd.t152 gnd 0.029274f
C2129 vdd.n1023 gnd 0.201188f
C2130 vdd.n1024 gnd 0.127669f
C2131 vdd.t137 gnd 0.029274f
C2132 vdd.t117 gnd 0.029274f
C2133 vdd.n1025 gnd 0.201188f
C2134 vdd.n1026 gnd 0.127669f
C2135 vdd.n1027 gnd 0.00499f
C2136 vdd.n1028 gnd 0.004631f
C2137 vdd.n1029 gnd 0.002561f
C2138 vdd.n1030 gnd 0.005881f
C2139 vdd.n1031 gnd 0.002488f
C2140 vdd.n1032 gnd 0.002635f
C2141 vdd.n1033 gnd 0.004631f
C2142 vdd.n1034 gnd 0.002488f
C2143 vdd.n1035 gnd 0.005881f
C2144 vdd.n1036 gnd 0.002635f
C2145 vdd.n1037 gnd 0.004631f
C2146 vdd.n1038 gnd 0.002488f
C2147 vdd.n1039 gnd 0.004411f
C2148 vdd.n1040 gnd 0.004424f
C2149 vdd.t150 gnd 0.012636f
C2150 vdd.n1041 gnd 0.028114f
C2151 vdd.n1042 gnd 0.146311f
C2152 vdd.n1043 gnd 0.002488f
C2153 vdd.n1044 gnd 0.002635f
C2154 vdd.n1045 gnd 0.005881f
C2155 vdd.n1046 gnd 0.005881f
C2156 vdd.n1047 gnd 0.002635f
C2157 vdd.n1048 gnd 0.002488f
C2158 vdd.n1049 gnd 0.004631f
C2159 vdd.n1050 gnd 0.004631f
C2160 vdd.n1051 gnd 0.002488f
C2161 vdd.n1052 gnd 0.002635f
C2162 vdd.n1053 gnd 0.005881f
C2163 vdd.n1054 gnd 0.005881f
C2164 vdd.n1055 gnd 0.002635f
C2165 vdd.n1056 gnd 0.002488f
C2166 vdd.n1057 gnd 0.004631f
C2167 vdd.n1058 gnd 0.004631f
C2168 vdd.n1059 gnd 0.002488f
C2169 vdd.n1060 gnd 0.002635f
C2170 vdd.n1061 gnd 0.005881f
C2171 vdd.n1062 gnd 0.005881f
C2172 vdd.n1063 gnd 0.013905f
C2173 vdd.n1064 gnd 0.002561f
C2174 vdd.n1065 gnd 0.002488f
C2175 vdd.n1066 gnd 0.011968f
C2176 vdd.n1067 gnd 0.008094f
C2177 vdd.n1068 gnd 0.056507f
C2178 vdd.n1069 gnd 0.203611f
C2179 vdd.n1070 gnd 0.00499f
C2180 vdd.n1071 gnd 0.004631f
C2181 vdd.n1072 gnd 0.002561f
C2182 vdd.n1073 gnd 0.005881f
C2183 vdd.n1074 gnd 0.002488f
C2184 vdd.n1075 gnd 0.002635f
C2185 vdd.n1076 gnd 0.004631f
C2186 vdd.n1077 gnd 0.002488f
C2187 vdd.n1078 gnd 0.005881f
C2188 vdd.n1079 gnd 0.002635f
C2189 vdd.n1080 gnd 0.004631f
C2190 vdd.n1081 gnd 0.002488f
C2191 vdd.n1082 gnd 0.004411f
C2192 vdd.n1083 gnd 0.004424f
C2193 vdd.t171 gnd 0.012636f
C2194 vdd.n1084 gnd 0.028114f
C2195 vdd.n1085 gnd 0.146311f
C2196 vdd.n1086 gnd 0.002488f
C2197 vdd.n1087 gnd 0.002635f
C2198 vdd.n1088 gnd 0.005881f
C2199 vdd.n1089 gnd 0.005881f
C2200 vdd.n1090 gnd 0.002635f
C2201 vdd.n1091 gnd 0.002488f
C2202 vdd.n1092 gnd 0.004631f
C2203 vdd.n1093 gnd 0.004631f
C2204 vdd.n1094 gnd 0.002488f
C2205 vdd.n1095 gnd 0.002635f
C2206 vdd.n1096 gnd 0.005881f
C2207 vdd.n1097 gnd 0.005881f
C2208 vdd.n1098 gnd 0.002635f
C2209 vdd.n1099 gnd 0.002488f
C2210 vdd.n1100 gnd 0.004631f
C2211 vdd.n1101 gnd 0.004631f
C2212 vdd.n1102 gnd 0.002488f
C2213 vdd.n1103 gnd 0.002635f
C2214 vdd.n1104 gnd 0.005881f
C2215 vdd.n1105 gnd 0.005881f
C2216 vdd.n1106 gnd 0.013905f
C2217 vdd.n1107 gnd 0.002561f
C2218 vdd.n1108 gnd 0.002488f
C2219 vdd.n1109 gnd 0.011968f
C2220 vdd.n1110 gnd 0.008356f
C2221 vdd.t126 gnd 0.029274f
C2222 vdd.t170 gnd 0.029274f
C2223 vdd.n1111 gnd 0.201188f
C2224 vdd.n1112 gnd 0.158204f
C2225 vdd.t169 gnd 0.029274f
C2226 vdd.t158 gnd 0.029274f
C2227 vdd.n1113 gnd 0.201188f
C2228 vdd.n1114 gnd 0.127669f
C2229 vdd.t145 gnd 0.029274f
C2230 vdd.t124 gnd 0.029274f
C2231 vdd.n1115 gnd 0.201188f
C2232 vdd.n1116 gnd 0.127669f
C2233 vdd.n1117 gnd 0.00499f
C2234 vdd.n1118 gnd 0.004631f
C2235 vdd.n1119 gnd 0.002561f
C2236 vdd.n1120 gnd 0.005881f
C2237 vdd.n1121 gnd 0.002488f
C2238 vdd.n1122 gnd 0.002635f
C2239 vdd.n1123 gnd 0.004631f
C2240 vdd.n1124 gnd 0.002488f
C2241 vdd.n1125 gnd 0.005881f
C2242 vdd.n1126 gnd 0.002635f
C2243 vdd.n1127 gnd 0.004631f
C2244 vdd.n1128 gnd 0.002488f
C2245 vdd.n1129 gnd 0.004411f
C2246 vdd.n1130 gnd 0.004424f
C2247 vdd.t157 gnd 0.012636f
C2248 vdd.n1131 gnd 0.028114f
C2249 vdd.n1132 gnd 0.146311f
C2250 vdd.n1133 gnd 0.002488f
C2251 vdd.n1134 gnd 0.002635f
C2252 vdd.n1135 gnd 0.005881f
C2253 vdd.n1136 gnd 0.005881f
C2254 vdd.n1137 gnd 0.002635f
C2255 vdd.n1138 gnd 0.002488f
C2256 vdd.n1139 gnd 0.004631f
C2257 vdd.n1140 gnd 0.004631f
C2258 vdd.n1141 gnd 0.002488f
C2259 vdd.n1142 gnd 0.002635f
C2260 vdd.n1143 gnd 0.005881f
C2261 vdd.n1144 gnd 0.005881f
C2262 vdd.n1145 gnd 0.002635f
C2263 vdd.n1146 gnd 0.002488f
C2264 vdd.n1147 gnd 0.004631f
C2265 vdd.n1148 gnd 0.004631f
C2266 vdd.n1149 gnd 0.002488f
C2267 vdd.n1150 gnd 0.002635f
C2268 vdd.n1151 gnd 0.005881f
C2269 vdd.n1152 gnd 0.005881f
C2270 vdd.n1153 gnd 0.013905f
C2271 vdd.n1154 gnd 0.002561f
C2272 vdd.n1155 gnd 0.002488f
C2273 vdd.n1156 gnd 0.011968f
C2274 vdd.n1157 gnd 0.008094f
C2275 vdd.n1158 gnd 0.056507f
C2276 vdd.n1159 gnd 0.220385f
C2277 vdd.n1160 gnd 1.85217f
C2278 vdd.n1161 gnd 0.536312f
C2279 vdd.n1162 gnd 0.007318f
C2280 vdd.n1163 gnd 0.009093f
C2281 vdd.n1164 gnd 0.571467f
C2282 vdd.n1165 gnd 0.009093f
C2283 vdd.n1166 gnd 0.007318f
C2284 vdd.n1167 gnd 0.009093f
C2285 vdd.n1168 gnd 0.007318f
C2286 vdd.n1169 gnd 0.009093f
C2287 vdd.t116 gnd 0.464607f
C2288 vdd.t127 gnd 0.464607f
C2289 vdd.n1170 gnd 0.009093f
C2290 vdd.n1171 gnd 0.007318f
C2291 vdd.n1172 gnd 0.009093f
C2292 vdd.n1173 gnd 0.007318f
C2293 vdd.n1174 gnd 0.009093f
C2294 vdd.t133 gnd 0.464607f
C2295 vdd.n1175 gnd 0.009093f
C2296 vdd.n1176 gnd 0.007318f
C2297 vdd.n1177 gnd 0.009093f
C2298 vdd.n1178 gnd 0.007318f
C2299 vdd.n1179 gnd 0.009093f
C2300 vdd.t149 gnd 0.464607f
C2301 vdd.n1180 gnd 0.67368f
C2302 vdd.n1181 gnd 0.009093f
C2303 vdd.n1182 gnd 0.007318f
C2304 vdd.n1183 gnd 0.009093f
C2305 vdd.n1184 gnd 0.007318f
C2306 vdd.n1185 gnd 0.009093f
C2307 vdd.n1186 gnd 0.929214f
C2308 vdd.n1187 gnd 0.009093f
C2309 vdd.n1188 gnd 0.007318f
C2310 vdd.n1189 gnd 0.022159f
C2311 vdd.n1190 gnd 0.006074f
C2312 vdd.n1191 gnd 0.022159f
C2313 vdd.t26 gnd 0.464607f
C2314 vdd.n1192 gnd 0.022159f
C2315 vdd.n1193 gnd 0.006074f
C2316 vdd.n1194 gnd 0.009093f
C2317 vdd.n1195 gnd 0.007318f
C2318 vdd.n1196 gnd 0.009093f
C2319 vdd.n1227 gnd 0.022667f
C2320 vdd.n1228 gnd 1.37059f
C2321 vdd.n1229 gnd 0.009093f
C2322 vdd.n1230 gnd 0.007318f
C2323 vdd.n1231 gnd 0.009093f
C2324 vdd.n1232 gnd 0.009093f
C2325 vdd.n1233 gnd 0.009093f
C2326 vdd.n1234 gnd 0.009093f
C2327 vdd.n1235 gnd 0.009093f
C2328 vdd.n1236 gnd 0.007318f
C2329 vdd.n1237 gnd 0.009093f
C2330 vdd.n1238 gnd 0.009093f
C2331 vdd.n1239 gnd 0.009093f
C2332 vdd.n1240 gnd 0.009093f
C2333 vdd.n1241 gnd 0.009093f
C2334 vdd.n1242 gnd 0.007318f
C2335 vdd.n1243 gnd 0.009093f
C2336 vdd.n1244 gnd 0.009093f
C2337 vdd.n1245 gnd 0.009093f
C2338 vdd.n1246 gnd 0.009093f
C2339 vdd.n1247 gnd 0.009093f
C2340 vdd.n1248 gnd 0.007318f
C2341 vdd.n1249 gnd 0.009093f
C2342 vdd.n1250 gnd 0.009093f
C2343 vdd.n1251 gnd 0.009093f
C2344 vdd.n1252 gnd 0.009093f
C2345 vdd.n1253 gnd 0.009093f
C2346 vdd.t76 gnd 0.111862f
C2347 vdd.t77 gnd 0.11955f
C2348 vdd.t75 gnd 0.14609f
C2349 vdd.n1254 gnd 0.187267f
C2350 vdd.n1255 gnd 0.15807f
C2351 vdd.n1256 gnd 0.015661f
C2352 vdd.n1257 gnd 0.009093f
C2353 vdd.n1258 gnd 0.009093f
C2354 vdd.n1259 gnd 0.009093f
C2355 vdd.n1260 gnd 0.009093f
C2356 vdd.n1261 gnd 0.009093f
C2357 vdd.n1262 gnd 0.007318f
C2358 vdd.n1263 gnd 0.009093f
C2359 vdd.n1264 gnd 0.009093f
C2360 vdd.n1265 gnd 0.009093f
C2361 vdd.n1266 gnd 0.009093f
C2362 vdd.n1267 gnd 0.009093f
C2363 vdd.n1268 gnd 0.007318f
C2364 vdd.n1269 gnd 0.009093f
C2365 vdd.n1270 gnd 0.009093f
C2366 vdd.n1271 gnd 0.009093f
C2367 vdd.n1272 gnd 0.009093f
C2368 vdd.n1273 gnd 0.009093f
C2369 vdd.n1274 gnd 0.007318f
C2370 vdd.n1275 gnd 0.009093f
C2371 vdd.n1276 gnd 0.009093f
C2372 vdd.n1277 gnd 0.009093f
C2373 vdd.n1278 gnd 0.009093f
C2374 vdd.n1279 gnd 0.009093f
C2375 vdd.n1280 gnd 0.007318f
C2376 vdd.n1281 gnd 0.009093f
C2377 vdd.n1282 gnd 0.009093f
C2378 vdd.n1283 gnd 0.009093f
C2379 vdd.n1284 gnd 0.009093f
C2380 vdd.n1285 gnd 0.009093f
C2381 vdd.n1286 gnd 0.007318f
C2382 vdd.n1287 gnd 0.009093f
C2383 vdd.n1288 gnd 0.009093f
C2384 vdd.n1289 gnd 0.009093f
C2385 vdd.n1290 gnd 0.009093f
C2386 vdd.n1291 gnd 0.007318f
C2387 vdd.n1292 gnd 0.009093f
C2388 vdd.n1293 gnd 0.009093f
C2389 vdd.n1294 gnd 0.009093f
C2390 vdd.n1295 gnd 0.009093f
C2391 vdd.n1296 gnd 0.009093f
C2392 vdd.n1297 gnd 0.007318f
C2393 vdd.n1298 gnd 0.009093f
C2394 vdd.n1299 gnd 0.009093f
C2395 vdd.n1300 gnd 0.009093f
C2396 vdd.n1301 gnd 0.009093f
C2397 vdd.n1302 gnd 0.009093f
C2398 vdd.n1303 gnd 0.007318f
C2399 vdd.n1304 gnd 0.009093f
C2400 vdd.n1305 gnd 0.009093f
C2401 vdd.n1306 gnd 0.009093f
C2402 vdd.n1307 gnd 0.009093f
C2403 vdd.n1308 gnd 0.009093f
C2404 vdd.n1309 gnd 0.007318f
C2405 vdd.n1310 gnd 0.009093f
C2406 vdd.n1311 gnd 0.009093f
C2407 vdd.n1312 gnd 0.009093f
C2408 vdd.n1313 gnd 0.009093f
C2409 vdd.n1314 gnd 0.009093f
C2410 vdd.n1315 gnd 0.007318f
C2411 vdd.n1316 gnd 0.009093f
C2412 vdd.n1317 gnd 0.009093f
C2413 vdd.n1318 gnd 0.009093f
C2414 vdd.n1319 gnd 0.009093f
C2415 vdd.t27 gnd 0.111862f
C2416 vdd.t28 gnd 0.11955f
C2417 vdd.t25 gnd 0.14609f
C2418 vdd.n1320 gnd 0.187267f
C2419 vdd.n1321 gnd 0.15807f
C2420 vdd.n1322 gnd 0.012002f
C2421 vdd.n1323 gnd 0.003476f
C2422 vdd.n1324 gnd 0.022667f
C2423 vdd.n1325 gnd 0.009093f
C2424 vdd.n1326 gnd 0.003842f
C2425 vdd.n1327 gnd 0.007318f
C2426 vdd.n1328 gnd 0.007318f
C2427 vdd.n1329 gnd 0.009093f
C2428 vdd.n1330 gnd 0.009093f
C2429 vdd.n1331 gnd 0.009093f
C2430 vdd.n1332 gnd 0.007318f
C2431 vdd.n1333 gnd 0.007318f
C2432 vdd.n1334 gnd 0.007318f
C2433 vdd.n1335 gnd 0.009093f
C2434 vdd.n1336 gnd 0.009093f
C2435 vdd.n1337 gnd 0.009093f
C2436 vdd.n1338 gnd 0.007318f
C2437 vdd.n1339 gnd 0.007318f
C2438 vdd.n1340 gnd 0.007318f
C2439 vdd.n1341 gnd 0.009093f
C2440 vdd.n1342 gnd 0.009093f
C2441 vdd.n1343 gnd 0.009093f
C2442 vdd.n1344 gnd 0.007318f
C2443 vdd.n1345 gnd 0.007318f
C2444 vdd.n1346 gnd 0.007318f
C2445 vdd.n1347 gnd 0.009093f
C2446 vdd.n1348 gnd 0.009093f
C2447 vdd.n1349 gnd 0.009093f
C2448 vdd.n1350 gnd 0.007318f
C2449 vdd.n1351 gnd 0.007318f
C2450 vdd.n1352 gnd 0.007318f
C2451 vdd.n1353 gnd 0.009093f
C2452 vdd.n1354 gnd 0.009093f
C2453 vdd.n1355 gnd 0.009093f
C2454 vdd.n1356 gnd 0.007245f
C2455 vdd.n1357 gnd 0.009093f
C2456 vdd.t73 gnd 0.111862f
C2457 vdd.t74 gnd 0.11955f
C2458 vdd.t72 gnd 0.14609f
C2459 vdd.n1358 gnd 0.187267f
C2460 vdd.n1359 gnd 0.15807f
C2461 vdd.n1360 gnd 0.015661f
C2462 vdd.n1361 gnd 0.004977f
C2463 vdd.n1362 gnd 0.009093f
C2464 vdd.n1363 gnd 0.009093f
C2465 vdd.n1364 gnd 0.009093f
C2466 vdd.n1365 gnd 0.007318f
C2467 vdd.n1366 gnd 0.007318f
C2468 vdd.n1367 gnd 0.007318f
C2469 vdd.n1368 gnd 0.009093f
C2470 vdd.n1369 gnd 0.009093f
C2471 vdd.n1370 gnd 0.009093f
C2472 vdd.n1371 gnd 0.007318f
C2473 vdd.n1372 gnd 0.007318f
C2474 vdd.n1373 gnd 0.007318f
C2475 vdd.n1374 gnd 0.009093f
C2476 vdd.n1375 gnd 0.009093f
C2477 vdd.n1376 gnd 0.009093f
C2478 vdd.n1377 gnd 0.007318f
C2479 vdd.n1378 gnd 0.007318f
C2480 vdd.n1379 gnd 0.007318f
C2481 vdd.n1380 gnd 0.009093f
C2482 vdd.n1381 gnd 0.009093f
C2483 vdd.n1382 gnd 0.009093f
C2484 vdd.n1383 gnd 0.007318f
C2485 vdd.n1384 gnd 0.007318f
C2486 vdd.n1385 gnd 0.007318f
C2487 vdd.n1386 gnd 0.009093f
C2488 vdd.n1387 gnd 0.009093f
C2489 vdd.n1388 gnd 0.009093f
C2490 vdd.n1389 gnd 0.007318f
C2491 vdd.n1390 gnd 0.007318f
C2492 vdd.n1391 gnd 0.006111f
C2493 vdd.n1392 gnd 0.009093f
C2494 vdd.n1393 gnd 0.009093f
C2495 vdd.n1394 gnd 0.009093f
C2496 vdd.n1395 gnd 0.006111f
C2497 vdd.n1396 gnd 0.007318f
C2498 vdd.n1397 gnd 0.007318f
C2499 vdd.n1398 gnd 0.009093f
C2500 vdd.n1399 gnd 0.009093f
C2501 vdd.n1400 gnd 0.009093f
C2502 vdd.n1401 gnd 0.007318f
C2503 vdd.n1402 gnd 0.007318f
C2504 vdd.n1403 gnd 0.007318f
C2505 vdd.n1404 gnd 0.009093f
C2506 vdd.n1405 gnd 0.009093f
C2507 vdd.n1406 gnd 0.009093f
C2508 vdd.n1407 gnd 0.007318f
C2509 vdd.n1408 gnd 0.007318f
C2510 vdd.n1409 gnd 0.007318f
C2511 vdd.n1410 gnd 0.009093f
C2512 vdd.n1411 gnd 0.009093f
C2513 vdd.n1412 gnd 0.009093f
C2514 vdd.n1413 gnd 0.007318f
C2515 vdd.n1414 gnd 0.007318f
C2516 vdd.n1415 gnd 0.007318f
C2517 vdd.n1416 gnd 0.009093f
C2518 vdd.n1417 gnd 0.009093f
C2519 vdd.n1418 gnd 0.009093f
C2520 vdd.n1419 gnd 0.007318f
C2521 vdd.n1420 gnd 0.009093f
C2522 vdd.n1421 gnd 2.22082f
C2523 vdd.n1423 gnd 0.022667f
C2524 vdd.n1424 gnd 0.006074f
C2525 vdd.n1425 gnd 0.022667f
C2526 vdd.n1426 gnd 0.022159f
C2527 vdd.n1427 gnd 0.009093f
C2528 vdd.n1428 gnd 0.007318f
C2529 vdd.n1429 gnd 0.009093f
C2530 vdd.n1430 gnd 0.487837f
C2531 vdd.n1431 gnd 0.009093f
C2532 vdd.n1432 gnd 0.007318f
C2533 vdd.n1433 gnd 0.009093f
C2534 vdd.n1434 gnd 0.009093f
C2535 vdd.n1435 gnd 0.009093f
C2536 vdd.n1436 gnd 0.007318f
C2537 vdd.n1437 gnd 0.009093f
C2538 vdd.n1438 gnd 0.831647f
C2539 vdd.n1439 gnd 0.929214f
C2540 vdd.n1440 gnd 0.009093f
C2541 vdd.n1441 gnd 0.007318f
C2542 vdd.n1442 gnd 0.009093f
C2543 vdd.n1443 gnd 0.009093f
C2544 vdd.n1444 gnd 0.009093f
C2545 vdd.n1445 gnd 0.007318f
C2546 vdd.n1446 gnd 0.009093f
C2547 vdd.n1447 gnd 0.562174f
C2548 vdd.n1448 gnd 0.009093f
C2549 vdd.n1449 gnd 0.007318f
C2550 vdd.n1450 gnd 0.009093f
C2551 vdd.n1451 gnd 0.009093f
C2552 vdd.n1452 gnd 0.009093f
C2553 vdd.n1453 gnd 0.007318f
C2554 vdd.n1454 gnd 0.009093f
C2555 vdd.n1455 gnd 0.515714f
C2556 vdd.n1456 gnd 0.720141f
C2557 vdd.n1457 gnd 0.009093f
C2558 vdd.n1458 gnd 0.007318f
C2559 vdd.n1459 gnd 0.009093f
C2560 vdd.n1460 gnd 0.009093f
C2561 vdd.n1461 gnd 0.006988f
C2562 vdd.n1462 gnd 0.009093f
C2563 vdd.n1463 gnd 0.007318f
C2564 vdd.n1464 gnd 0.009093f
C2565 vdd.n1465 gnd 0.771248f
C2566 vdd.n1466 gnd 0.009093f
C2567 vdd.n1467 gnd 0.007318f
C2568 vdd.n1468 gnd 0.009093f
C2569 vdd.n1469 gnd 0.009093f
C2570 vdd.n1470 gnd 0.009093f
C2571 vdd.n1471 gnd 0.007318f
C2572 vdd.n1472 gnd 0.009093f
C2573 vdd.t151 gnd 0.464607f
C2574 vdd.n1473 gnd 0.664388f
C2575 vdd.n1474 gnd 0.009093f
C2576 vdd.n1475 gnd 0.007318f
C2577 vdd.n1476 gnd 0.006988f
C2578 vdd.n1477 gnd 0.009093f
C2579 vdd.n1478 gnd 0.009093f
C2580 vdd.n1479 gnd 0.007318f
C2581 vdd.n1480 gnd 0.009093f
C2582 vdd.n1481 gnd 0.506422f
C2583 vdd.n1482 gnd 0.009093f
C2584 vdd.n1483 gnd 0.007318f
C2585 vdd.n1484 gnd 0.009093f
C2586 vdd.n1485 gnd 0.009093f
C2587 vdd.n1486 gnd 0.009093f
C2588 vdd.n1487 gnd 0.007318f
C2589 vdd.n1488 gnd 0.009093f
C2590 vdd.n1489 gnd 0.655096f
C2591 vdd.n1490 gnd 0.580759f
C2592 vdd.n1491 gnd 0.009093f
C2593 vdd.n1492 gnd 0.007318f
C2594 vdd.n1493 gnd 0.009093f
C2595 vdd.n1494 gnd 0.009093f
C2596 vdd.n1495 gnd 0.009093f
C2597 vdd.n1496 gnd 0.007318f
C2598 vdd.n1497 gnd 0.009093f
C2599 vdd.n1498 gnd 0.738725f
C2600 vdd.n1499 gnd 0.009093f
C2601 vdd.n1500 gnd 0.007318f
C2602 vdd.n1501 gnd 0.009093f
C2603 vdd.n1502 gnd 0.009093f
C2604 vdd.n1503 gnd 0.022159f
C2605 vdd.n1504 gnd 0.009093f
C2606 vdd.n1505 gnd 0.009093f
C2607 vdd.n1506 gnd 0.007318f
C2608 vdd.n1507 gnd 0.009093f
C2609 vdd.n1508 gnd 0.580759f
C2610 vdd.n1509 gnd 0.929214f
C2611 vdd.n1510 gnd 0.009093f
C2612 vdd.n1511 gnd 0.007318f
C2613 vdd.n1512 gnd 0.009093f
C2614 vdd.n1513 gnd 0.009093f
C2615 vdd.n1514 gnd 0.00782f
C2616 vdd.n1515 gnd 0.007318f
C2617 vdd.n1517 gnd 0.009093f
C2618 vdd.n1519 gnd 0.007318f
C2619 vdd.n1520 gnd 0.009093f
C2620 vdd.n1521 gnd 0.007318f
C2621 vdd.n1523 gnd 0.009093f
C2622 vdd.n1524 gnd 0.007318f
C2623 vdd.n1525 gnd 0.009093f
C2624 vdd.n1526 gnd 0.009093f
C2625 vdd.n1527 gnd 0.009093f
C2626 vdd.n1528 gnd 0.009093f
C2627 vdd.n1529 gnd 0.009093f
C2628 vdd.n1530 gnd 0.007318f
C2629 vdd.n1532 gnd 0.009093f
C2630 vdd.n1533 gnd 0.009093f
C2631 vdd.n1534 gnd 0.009093f
C2632 vdd.n1535 gnd 0.009093f
C2633 vdd.n1536 gnd 0.009093f
C2634 vdd.n1537 gnd 0.007318f
C2635 vdd.n1539 gnd 0.009093f
C2636 vdd.n1540 gnd 0.009093f
C2637 vdd.n1541 gnd 0.009093f
C2638 vdd.n1542 gnd 0.009093f
C2639 vdd.n1543 gnd 0.006111f
C2640 vdd.t42 gnd 0.111862f
C2641 vdd.t41 gnd 0.11955f
C2642 vdd.t40 gnd 0.14609f
C2643 vdd.n1544 gnd 0.187267f
C2644 vdd.n1545 gnd 0.157338f
C2645 vdd.n1547 gnd 0.009093f
C2646 vdd.n1548 gnd 0.009093f
C2647 vdd.n1549 gnd 0.007318f
C2648 vdd.n1550 gnd 0.009093f
C2649 vdd.n1552 gnd 0.009093f
C2650 vdd.n1553 gnd 0.009093f
C2651 vdd.n1554 gnd 0.009093f
C2652 vdd.n1555 gnd 0.009093f
C2653 vdd.n1556 gnd 0.007318f
C2654 vdd.n1558 gnd 0.009093f
C2655 vdd.n1559 gnd 0.009093f
C2656 vdd.n1560 gnd 0.009093f
C2657 vdd.n1561 gnd 0.009093f
C2658 vdd.n1562 gnd 0.009093f
C2659 vdd.n1563 gnd 0.007318f
C2660 vdd.n1565 gnd 0.009093f
C2661 vdd.n1566 gnd 0.009093f
C2662 vdd.n1567 gnd 0.009093f
C2663 vdd.n1568 gnd 0.009093f
C2664 vdd.n1569 gnd 0.009093f
C2665 vdd.n1570 gnd 0.007318f
C2666 vdd.n1572 gnd 0.009093f
C2667 vdd.n1573 gnd 0.009093f
C2668 vdd.n1574 gnd 0.009093f
C2669 vdd.n1575 gnd 0.009093f
C2670 vdd.n1576 gnd 0.009093f
C2671 vdd.n1577 gnd 0.007318f
C2672 vdd.n1579 gnd 0.009093f
C2673 vdd.n1580 gnd 0.009093f
C2674 vdd.n1581 gnd 0.009093f
C2675 vdd.n1582 gnd 0.009093f
C2676 vdd.n1583 gnd 0.007245f
C2677 vdd.t35 gnd 0.111862f
C2678 vdd.t34 gnd 0.11955f
C2679 vdd.t33 gnd 0.14609f
C2680 vdd.n1584 gnd 0.187267f
C2681 vdd.n1585 gnd 0.157338f
C2682 vdd.n1587 gnd 0.009093f
C2683 vdd.n1588 gnd 0.009093f
C2684 vdd.n1589 gnd 0.007318f
C2685 vdd.n1590 gnd 0.009093f
C2686 vdd.n1592 gnd 0.009093f
C2687 vdd.n1593 gnd 0.009093f
C2688 vdd.n1594 gnd 0.009093f
C2689 vdd.n1595 gnd 0.009093f
C2690 vdd.n1596 gnd 0.007318f
C2691 vdd.n1598 gnd 0.009093f
C2692 vdd.n1599 gnd 0.009093f
C2693 vdd.n1600 gnd 0.009093f
C2694 vdd.n1601 gnd 0.009093f
C2695 vdd.n1602 gnd 0.009093f
C2696 vdd.n1603 gnd 0.007318f
C2697 vdd.n1605 gnd 0.009093f
C2698 vdd.n1606 gnd 0.009093f
C2699 vdd.n1607 gnd 0.009093f
C2700 vdd.n1608 gnd 0.009093f
C2701 vdd.n1609 gnd 0.009093f
C2702 vdd.n1610 gnd 0.009093f
C2703 vdd.n1611 gnd 0.007318f
C2704 vdd.n1613 gnd 0.009093f
C2705 vdd.n1615 gnd 0.009093f
C2706 vdd.n1616 gnd 0.007318f
C2707 vdd.n1617 gnd 0.007318f
C2708 vdd.n1618 gnd 0.009093f
C2709 vdd.n1620 gnd 0.009093f
C2710 vdd.n1621 gnd 0.007318f
C2711 vdd.n1622 gnd 0.007318f
C2712 vdd.n1623 gnd 0.009093f
C2713 vdd.n1625 gnd 0.009093f
C2714 vdd.n1626 gnd 0.009093f
C2715 vdd.n1627 gnd 0.007318f
C2716 vdd.n1628 gnd 0.007318f
C2717 vdd.n1629 gnd 0.007318f
C2718 vdd.n1630 gnd 0.009093f
C2719 vdd.n1632 gnd 0.009093f
C2720 vdd.n1633 gnd 0.009093f
C2721 vdd.n1634 gnd 0.007318f
C2722 vdd.n1635 gnd 0.007318f
C2723 vdd.n1636 gnd 0.007318f
C2724 vdd.n1637 gnd 0.009093f
C2725 vdd.n1639 gnd 0.009093f
C2726 vdd.n1640 gnd 0.009093f
C2727 vdd.n1641 gnd 0.007318f
C2728 vdd.n1642 gnd 0.007318f
C2729 vdd.n1643 gnd 0.007318f
C2730 vdd.n1644 gnd 0.009093f
C2731 vdd.n1646 gnd 0.009093f
C2732 vdd.n1647 gnd 0.009093f
C2733 vdd.n1648 gnd 0.007318f
C2734 vdd.n1649 gnd 0.009093f
C2735 vdd.n1650 gnd 0.009093f
C2736 vdd.n1651 gnd 0.009093f
C2737 vdd.n1652 gnd 0.01493f
C2738 vdd.n1653 gnd 0.004977f
C2739 vdd.n1654 gnd 0.007318f
C2740 vdd.n1655 gnd 0.009093f
C2741 vdd.n1657 gnd 0.009093f
C2742 vdd.n1658 gnd 0.009093f
C2743 vdd.n1659 gnd 0.007318f
C2744 vdd.n1660 gnd 0.007318f
C2745 vdd.n1661 gnd 0.007318f
C2746 vdd.n1662 gnd 0.009093f
C2747 vdd.n1664 gnd 0.009093f
C2748 vdd.n1665 gnd 0.009093f
C2749 vdd.n1666 gnd 0.007318f
C2750 vdd.n1667 gnd 0.007318f
C2751 vdd.n1668 gnd 0.007318f
C2752 vdd.n1669 gnd 0.009093f
C2753 vdd.n1671 gnd 0.009093f
C2754 vdd.n1672 gnd 0.009093f
C2755 vdd.n1673 gnd 0.007318f
C2756 vdd.n1674 gnd 0.007318f
C2757 vdd.n1675 gnd 0.007318f
C2758 vdd.n1676 gnd 0.009093f
C2759 vdd.n1678 gnd 0.009093f
C2760 vdd.n1679 gnd 0.009093f
C2761 vdd.n1680 gnd 0.007318f
C2762 vdd.n1681 gnd 0.007318f
C2763 vdd.n1682 gnd 0.007318f
C2764 vdd.n1683 gnd 0.009093f
C2765 vdd.n1685 gnd 0.009093f
C2766 vdd.n1686 gnd 0.009093f
C2767 vdd.n1687 gnd 0.007318f
C2768 vdd.n1688 gnd 0.009093f
C2769 vdd.n1689 gnd 0.009093f
C2770 vdd.n1690 gnd 0.009093f
C2771 vdd.n1691 gnd 0.01493f
C2772 vdd.n1692 gnd 0.006111f
C2773 vdd.n1693 gnd 0.007318f
C2774 vdd.n1694 gnd 0.009093f
C2775 vdd.n1696 gnd 0.009093f
C2776 vdd.n1697 gnd 0.009093f
C2777 vdd.n1698 gnd 0.007318f
C2778 vdd.n1699 gnd 0.007318f
C2779 vdd.n1700 gnd 0.007318f
C2780 vdd.n1701 gnd 0.009093f
C2781 vdd.n1703 gnd 0.009093f
C2782 vdd.n1704 gnd 0.009093f
C2783 vdd.n1705 gnd 0.007318f
C2784 vdd.n1706 gnd 0.007318f
C2785 vdd.n1707 gnd 0.007318f
C2786 vdd.n1708 gnd 0.009093f
C2787 vdd.n1710 gnd 0.009093f
C2788 vdd.n1711 gnd 0.009093f
C2789 vdd.n1713 gnd 0.009093f
C2790 vdd.n1714 gnd 0.007318f
C2791 vdd.n1715 gnd 0.005819f
C2792 vdd.n1716 gnd 0.006183f
C2793 vdd.n1717 gnd 0.006183f
C2794 vdd.n1718 gnd 0.006183f
C2795 vdd.n1719 gnd 0.006183f
C2796 vdd.n1720 gnd 0.006183f
C2797 vdd.n1721 gnd 0.006183f
C2798 vdd.n1722 gnd 0.006183f
C2799 vdd.n1723 gnd 0.006183f
C2800 vdd.n1725 gnd 0.006183f
C2801 vdd.n1726 gnd 0.006183f
C2802 vdd.n1727 gnd 0.006183f
C2803 vdd.n1728 gnd 0.006183f
C2804 vdd.n1729 gnd 0.006183f
C2805 vdd.n1731 gnd 0.006183f
C2806 vdd.n1733 gnd 0.006183f
C2807 vdd.n1734 gnd 0.006183f
C2808 vdd.n1735 gnd 0.006183f
C2809 vdd.n1736 gnd 0.006183f
C2810 vdd.n1737 gnd 0.006183f
C2811 vdd.n1739 gnd 0.006183f
C2812 vdd.n1741 gnd 0.006183f
C2813 vdd.n1742 gnd 0.006183f
C2814 vdd.n1743 gnd 0.006183f
C2815 vdd.n1744 gnd 0.006183f
C2816 vdd.n1745 gnd 0.006183f
C2817 vdd.n1747 gnd 0.006183f
C2818 vdd.n1749 gnd 0.006183f
C2819 vdd.n1750 gnd 0.006183f
C2820 vdd.n1751 gnd 0.006183f
C2821 vdd.n1752 gnd 0.006183f
C2822 vdd.n1753 gnd 0.006183f
C2823 vdd.n1755 gnd 0.006183f
C2824 vdd.n1756 gnd 0.006183f
C2825 vdd.n1757 gnd 0.006183f
C2826 vdd.n1758 gnd 0.006183f
C2827 vdd.n1759 gnd 0.006183f
C2828 vdd.n1760 gnd 0.006183f
C2829 vdd.n1761 gnd 0.006183f
C2830 vdd.n1762 gnd 0.006183f
C2831 vdd.n1763 gnd 0.004501f
C2832 vdd.n1764 gnd 0.006183f
C2833 vdd.t88 gnd 0.249851f
C2834 vdd.t89 gnd 0.255754f
C2835 vdd.t87 gnd 0.163112f
C2836 vdd.n1765 gnd 0.088153f
C2837 vdd.n1766 gnd 0.050003f
C2838 vdd.n1767 gnd 0.008836f
C2839 vdd.n1768 gnd 0.006183f
C2840 vdd.n1769 gnd 0.006183f
C2841 vdd.n1770 gnd 0.376332f
C2842 vdd.n1771 gnd 0.006183f
C2843 vdd.n1772 gnd 0.006183f
C2844 vdd.n1773 gnd 0.006183f
C2845 vdd.n1774 gnd 0.006183f
C2846 vdd.n1775 gnd 0.006183f
C2847 vdd.n1776 gnd 0.006183f
C2848 vdd.n1777 gnd 0.006183f
C2849 vdd.n1778 gnd 0.006183f
C2850 vdd.n1779 gnd 0.006183f
C2851 vdd.n1780 gnd 0.006183f
C2852 vdd.n1781 gnd 0.006183f
C2853 vdd.n1782 gnd 0.006183f
C2854 vdd.n1783 gnd 0.006183f
C2855 vdd.n1784 gnd 0.006183f
C2856 vdd.n1785 gnd 0.006183f
C2857 vdd.n1786 gnd 0.006183f
C2858 vdd.n1787 gnd 0.006183f
C2859 vdd.n1788 gnd 0.006183f
C2860 vdd.n1789 gnd 0.006183f
C2861 vdd.n1790 gnd 0.006183f
C2862 vdd.t63 gnd 0.249851f
C2863 vdd.t64 gnd 0.255754f
C2864 vdd.t61 gnd 0.163112f
C2865 vdd.n1791 gnd 0.088153f
C2866 vdd.n1792 gnd 0.050003f
C2867 vdd.n1793 gnd 0.006183f
C2868 vdd.n1794 gnd 0.006183f
C2869 vdd.n1795 gnd 0.006183f
C2870 vdd.n1796 gnd 0.006183f
C2871 vdd.n1797 gnd 0.006183f
C2872 vdd.n1798 gnd 0.006183f
C2873 vdd.n1800 gnd 0.006183f
C2874 vdd.n1801 gnd 0.006183f
C2875 vdd.n1802 gnd 0.006183f
C2876 vdd.n1803 gnd 0.006183f
C2877 vdd.n1805 gnd 0.006183f
C2878 vdd.n1807 gnd 0.006183f
C2879 vdd.n1808 gnd 0.006183f
C2880 vdd.n1809 gnd 0.006183f
C2881 vdd.n1810 gnd 0.006183f
C2882 vdd.n1811 gnd 0.006183f
C2883 vdd.n1813 gnd 0.006183f
C2884 vdd.n1815 gnd 0.006183f
C2885 vdd.n1816 gnd 0.006183f
C2886 vdd.n1817 gnd 0.006183f
C2887 vdd.n1818 gnd 0.006183f
C2888 vdd.n1819 gnd 0.006183f
C2889 vdd.n1821 gnd 0.006183f
C2890 vdd.n1823 gnd 0.006183f
C2891 vdd.n1824 gnd 0.006183f
C2892 vdd.n1825 gnd 0.004501f
C2893 vdd.n1826 gnd 0.008836f
C2894 vdd.n1827 gnd 0.004774f
C2895 vdd.n1828 gnd 0.006183f
C2896 vdd.n1830 gnd 0.006183f
C2897 vdd.n1831 gnd 0.014671f
C2898 vdd.n1832 gnd 0.014671f
C2899 vdd.n1833 gnd 0.013698f
C2900 vdd.n1834 gnd 0.006183f
C2901 vdd.n1835 gnd 0.006183f
C2902 vdd.n1836 gnd 0.006183f
C2903 vdd.n1837 gnd 0.006183f
C2904 vdd.n1838 gnd 0.006183f
C2905 vdd.n1839 gnd 0.006183f
C2906 vdd.n1840 gnd 0.006183f
C2907 vdd.n1841 gnd 0.006183f
C2908 vdd.n1842 gnd 0.006183f
C2909 vdd.n1843 gnd 0.006183f
C2910 vdd.n1844 gnd 0.006183f
C2911 vdd.n1845 gnd 0.006183f
C2912 vdd.n1846 gnd 0.006183f
C2913 vdd.n1847 gnd 0.006183f
C2914 vdd.n1848 gnd 0.006183f
C2915 vdd.n1849 gnd 0.006183f
C2916 vdd.n1850 gnd 0.006183f
C2917 vdd.n1851 gnd 0.006183f
C2918 vdd.n1852 gnd 0.006183f
C2919 vdd.n1853 gnd 0.006183f
C2920 vdd.n1854 gnd 0.006183f
C2921 vdd.n1855 gnd 0.006183f
C2922 vdd.n1856 gnd 0.006183f
C2923 vdd.n1857 gnd 0.006183f
C2924 vdd.n1858 gnd 0.006183f
C2925 vdd.n1859 gnd 0.006183f
C2926 vdd.n1860 gnd 0.006183f
C2927 vdd.n1861 gnd 0.006183f
C2928 vdd.n1862 gnd 0.006183f
C2929 vdd.n1863 gnd 0.006183f
C2930 vdd.n1864 gnd 0.006183f
C2931 vdd.n1865 gnd 0.006183f
C2932 vdd.n1866 gnd 0.006183f
C2933 vdd.n1867 gnd 0.006183f
C2934 vdd.n1868 gnd 0.006183f
C2935 vdd.n1869 gnd 0.006183f
C2936 vdd.n1870 gnd 0.006183f
C2937 vdd.n1871 gnd 0.199781f
C2938 vdd.n1872 gnd 0.006183f
C2939 vdd.n1873 gnd 0.006183f
C2940 vdd.n1874 gnd 0.006183f
C2941 vdd.n1875 gnd 0.006183f
C2942 vdd.n1876 gnd 0.006183f
C2943 vdd.n1877 gnd 0.006183f
C2944 vdd.n1878 gnd 0.006183f
C2945 vdd.n1879 gnd 0.006183f
C2946 vdd.n1880 gnd 0.006183f
C2947 vdd.n1881 gnd 0.006183f
C2948 vdd.n1882 gnd 0.006183f
C2949 vdd.n1883 gnd 0.006183f
C2950 vdd.n1884 gnd 0.006183f
C2951 vdd.n1885 gnd 0.006183f
C2952 vdd.n1886 gnd 0.006183f
C2953 vdd.n1887 gnd 0.006183f
C2954 vdd.n1888 gnd 0.006183f
C2955 vdd.n1889 gnd 0.006183f
C2956 vdd.n1890 gnd 0.006183f
C2957 vdd.n1891 gnd 0.006183f
C2958 vdd.n1892 gnd 0.013698f
C2959 vdd.n1894 gnd 0.014671f
C2960 vdd.n1895 gnd 0.014671f
C2961 vdd.n1896 gnd 0.006183f
C2962 vdd.n1897 gnd 0.004774f
C2963 vdd.n1898 gnd 0.006183f
C2964 vdd.n1900 gnd 0.006183f
C2965 vdd.n1902 gnd 0.006183f
C2966 vdd.n1903 gnd 0.006183f
C2967 vdd.n1904 gnd 0.006183f
C2968 vdd.n1905 gnd 0.006183f
C2969 vdd.n1906 gnd 0.006183f
C2970 vdd.n1908 gnd 0.006183f
C2971 vdd.n1910 gnd 0.006183f
C2972 vdd.n1911 gnd 0.006183f
C2973 vdd.n1912 gnd 0.006183f
C2974 vdd.n1913 gnd 0.006183f
C2975 vdd.n1914 gnd 0.006183f
C2976 vdd.n1916 gnd 0.006183f
C2977 vdd.n1918 gnd 0.006183f
C2978 vdd.n1919 gnd 0.006183f
C2979 vdd.n1920 gnd 0.006183f
C2980 vdd.n1921 gnd 0.006183f
C2981 vdd.n1922 gnd 0.006183f
C2982 vdd.n1924 gnd 0.006183f
C2983 vdd.n1926 gnd 0.006183f
C2984 vdd.n1927 gnd 0.006183f
C2985 vdd.n1928 gnd 0.018442f
C2986 vdd.n1929 gnd 0.546711f
C2987 vdd.n1931 gnd 0.007318f
C2988 vdd.n1932 gnd 0.007318f
C2989 vdd.n1933 gnd 0.009093f
C2990 vdd.n1935 gnd 0.009093f
C2991 vdd.n1936 gnd 0.009093f
C2992 vdd.n1937 gnd 0.007318f
C2993 vdd.n1938 gnd 0.006074f
C2994 vdd.n1939 gnd 0.022667f
C2995 vdd.n1940 gnd 0.022159f
C2996 vdd.n1941 gnd 0.006074f
C2997 vdd.n1942 gnd 0.022159f
C2998 vdd.n1943 gnd 1.27767f
C2999 vdd.n1944 gnd 0.022159f
C3000 vdd.n1945 gnd 0.022667f
C3001 vdd.n1946 gnd 0.003476f
C3002 vdd.t24 gnd 0.111862f
C3003 vdd.t23 gnd 0.11955f
C3004 vdd.t21 gnd 0.14609f
C3005 vdd.n1947 gnd 0.187267f
C3006 vdd.n1948 gnd 0.157338f
C3007 vdd.n1949 gnd 0.01127f
C3008 vdd.n1950 gnd 0.003842f
C3009 vdd.n1951 gnd 0.00782f
C3010 vdd.n1952 gnd 0.546711f
C3011 vdd.n1953 gnd 0.018442f
C3012 vdd.n1954 gnd 0.006183f
C3013 vdd.n1955 gnd 0.006183f
C3014 vdd.n1956 gnd 0.006183f
C3015 vdd.n1958 gnd 0.006183f
C3016 vdd.n1960 gnd 0.006183f
C3017 vdd.n1961 gnd 0.006183f
C3018 vdd.n1962 gnd 0.006183f
C3019 vdd.n1963 gnd 0.006183f
C3020 vdd.n1964 gnd 0.006183f
C3021 vdd.n1966 gnd 0.006183f
C3022 vdd.n1968 gnd 0.006183f
C3023 vdd.n1969 gnd 0.006183f
C3024 vdd.n1970 gnd 0.006183f
C3025 vdd.n1971 gnd 0.006183f
C3026 vdd.n1972 gnd 0.006183f
C3027 vdd.n1974 gnd 0.006183f
C3028 vdd.n1976 gnd 0.006183f
C3029 vdd.n1977 gnd 0.006183f
C3030 vdd.n1978 gnd 0.006183f
C3031 vdd.n1979 gnd 0.006183f
C3032 vdd.n1980 gnd 0.006183f
C3033 vdd.n1982 gnd 0.006183f
C3034 vdd.n1984 gnd 0.006183f
C3035 vdd.n1985 gnd 0.006183f
C3036 vdd.n1986 gnd 0.014671f
C3037 vdd.n1987 gnd 0.013698f
C3038 vdd.n1988 gnd 0.013698f
C3039 vdd.n1989 gnd 0.91063f
C3040 vdd.n1990 gnd 0.013698f
C3041 vdd.n1991 gnd 0.013698f
C3042 vdd.n1992 gnd 0.006183f
C3043 vdd.n1993 gnd 0.006183f
C3044 vdd.n1994 gnd 0.006183f
C3045 vdd.n1995 gnd 0.394916f
C3046 vdd.n1996 gnd 0.006183f
C3047 vdd.n1997 gnd 0.006183f
C3048 vdd.n1998 gnd 0.006183f
C3049 vdd.n1999 gnd 0.006183f
C3050 vdd.n2000 gnd 0.006183f
C3051 vdd.n2001 gnd 0.631866f
C3052 vdd.n2002 gnd 0.006183f
C3053 vdd.n2003 gnd 0.006183f
C3054 vdd.n2004 gnd 0.006183f
C3055 vdd.n2005 gnd 0.006183f
C3056 vdd.n2006 gnd 0.006183f
C3057 vdd.n2007 gnd 0.631866f
C3058 vdd.n2008 gnd 0.006183f
C3059 vdd.n2009 gnd 0.006183f
C3060 vdd.n2010 gnd 0.005456f
C3061 vdd.n2011 gnd 0.017911f
C3062 vdd.n2012 gnd 0.003819f
C3063 vdd.n2013 gnd 0.006183f
C3064 vdd.n2014 gnd 0.348455f
C3065 vdd.n2015 gnd 0.006183f
C3066 vdd.n2016 gnd 0.006183f
C3067 vdd.n2017 gnd 0.006183f
C3068 vdd.n2018 gnd 0.006183f
C3069 vdd.n2019 gnd 0.006183f
C3070 vdd.n2020 gnd 0.422792f
C3071 vdd.n2021 gnd 0.006183f
C3072 vdd.n2022 gnd 0.006183f
C3073 vdd.n2023 gnd 0.006183f
C3074 vdd.n2024 gnd 0.006183f
C3075 vdd.n2025 gnd 0.006183f
C3076 vdd.n2026 gnd 0.562174f
C3077 vdd.n2027 gnd 0.006183f
C3078 vdd.n2028 gnd 0.006183f
C3079 vdd.n2029 gnd 0.006183f
C3080 vdd.n2030 gnd 0.006183f
C3081 vdd.n2031 gnd 0.006183f
C3082 vdd.n2032 gnd 0.501776f
C3083 vdd.n2033 gnd 0.006183f
C3084 vdd.n2034 gnd 0.006183f
C3085 vdd.n2035 gnd 0.006183f
C3086 vdd.n2036 gnd 0.006183f
C3087 vdd.n2037 gnd 0.006183f
C3088 vdd.n2038 gnd 0.362393f
C3089 vdd.n2039 gnd 0.006183f
C3090 vdd.n2040 gnd 0.006183f
C3091 vdd.n2041 gnd 0.006183f
C3092 vdd.n2042 gnd 0.006183f
C3093 vdd.n2043 gnd 0.006183f
C3094 vdd.n2044 gnd 0.199781f
C3095 vdd.n2045 gnd 0.006183f
C3096 vdd.n2046 gnd 0.006183f
C3097 vdd.n2047 gnd 0.006183f
C3098 vdd.n2048 gnd 0.006183f
C3099 vdd.n2049 gnd 0.006183f
C3100 vdd.n2050 gnd 0.348455f
C3101 vdd.n2051 gnd 0.006183f
C3102 vdd.n2052 gnd 0.006183f
C3103 vdd.n2053 gnd 0.006183f
C3104 vdd.n2054 gnd 0.006183f
C3105 vdd.n2055 gnd 0.006183f
C3106 vdd.n2056 gnd 0.631866f
C3107 vdd.n2057 gnd 0.006183f
C3108 vdd.n2058 gnd 0.006183f
C3109 vdd.n2059 gnd 0.006183f
C3110 vdd.n2060 gnd 0.006183f
C3111 vdd.n2061 gnd 0.006183f
C3112 vdd.n2062 gnd 0.006183f
C3113 vdd.n2063 gnd 0.006183f
C3114 vdd.n2064 gnd 0.492483f
C3115 vdd.n2065 gnd 0.006183f
C3116 vdd.n2066 gnd 0.006183f
C3117 vdd.n2067 gnd 0.006183f
C3118 vdd.n2068 gnd 0.006183f
C3119 vdd.n2069 gnd 0.006183f
C3120 vdd.n2070 gnd 0.006183f
C3121 vdd.n2071 gnd 0.394916f
C3122 vdd.n2072 gnd 0.006183f
C3123 vdd.n2073 gnd 0.006183f
C3124 vdd.n2074 gnd 0.006183f
C3125 vdd.n2075 gnd 0.014451f
C3126 vdd.n2076 gnd 0.013918f
C3127 vdd.n2077 gnd 0.006183f
C3128 vdd.n2078 gnd 0.006183f
C3129 vdd.n2079 gnd 0.004774f
C3130 vdd.n2080 gnd 0.006183f
C3131 vdd.n2081 gnd 0.006183f
C3132 vdd.n2082 gnd 0.004501f
C3133 vdd.n2083 gnd 0.006183f
C3134 vdd.n2084 gnd 0.006183f
C3135 vdd.n2085 gnd 0.006183f
C3136 vdd.n2086 gnd 0.006183f
C3137 vdd.n2087 gnd 0.006183f
C3138 vdd.n2088 gnd 0.006183f
C3139 vdd.n2089 gnd 0.006183f
C3140 vdd.n2090 gnd 0.006183f
C3141 vdd.n2091 gnd 0.006183f
C3142 vdd.n2092 gnd 0.006183f
C3143 vdd.n2093 gnd 0.006183f
C3144 vdd.n2094 gnd 0.006183f
C3145 vdd.n2095 gnd 0.006183f
C3146 vdd.n2096 gnd 0.006183f
C3147 vdd.n2097 gnd 0.006183f
C3148 vdd.n2098 gnd 0.006183f
C3149 vdd.n2099 gnd 0.006183f
C3150 vdd.n2100 gnd 0.006183f
C3151 vdd.n2101 gnd 0.006183f
C3152 vdd.n2102 gnd 0.006183f
C3153 vdd.n2103 gnd 0.006183f
C3154 vdd.n2104 gnd 0.006183f
C3155 vdd.n2105 gnd 0.006183f
C3156 vdd.n2106 gnd 0.006183f
C3157 vdd.n2107 gnd 0.006183f
C3158 vdd.n2108 gnd 0.006183f
C3159 vdd.n2109 gnd 0.006183f
C3160 vdd.n2110 gnd 0.006183f
C3161 vdd.n2111 gnd 0.006183f
C3162 vdd.n2112 gnd 0.006183f
C3163 vdd.n2113 gnd 0.006183f
C3164 vdd.n2114 gnd 0.006183f
C3165 vdd.n2115 gnd 0.006183f
C3166 vdd.n2116 gnd 0.006183f
C3167 vdd.n2117 gnd 0.006183f
C3168 vdd.n2118 gnd 0.006183f
C3169 vdd.n2119 gnd 0.006183f
C3170 vdd.n2120 gnd 0.006183f
C3171 vdd.n2121 gnd 0.006183f
C3172 vdd.n2122 gnd 0.006183f
C3173 vdd.n2123 gnd 0.006183f
C3174 vdd.n2124 gnd 0.006183f
C3175 vdd.n2125 gnd 0.006183f
C3176 vdd.n2126 gnd 0.006183f
C3177 vdd.n2127 gnd 0.006183f
C3178 vdd.n2128 gnd 0.006183f
C3179 vdd.n2129 gnd 0.006183f
C3180 vdd.n2130 gnd 0.006183f
C3181 vdd.n2131 gnd 0.006183f
C3182 vdd.n2132 gnd 0.006183f
C3183 vdd.n2133 gnd 0.006183f
C3184 vdd.n2134 gnd 0.006183f
C3185 vdd.n2135 gnd 0.006183f
C3186 vdd.n2136 gnd 0.006183f
C3187 vdd.n2137 gnd 0.006183f
C3188 vdd.n2138 gnd 0.006183f
C3189 vdd.n2139 gnd 0.006183f
C3190 vdd.n2140 gnd 0.006183f
C3191 vdd.n2141 gnd 0.006183f
C3192 vdd.n2142 gnd 0.006183f
C3193 vdd.n2143 gnd 0.014671f
C3194 vdd.n2144 gnd 0.013698f
C3195 vdd.n2145 gnd 0.013698f
C3196 vdd.n2146 gnd 0.771248f
C3197 vdd.n2147 gnd 0.013698f
C3198 vdd.n2148 gnd 0.014671f
C3199 vdd.n2149 gnd 0.013918f
C3200 vdd.n2150 gnd 0.006183f
C3201 vdd.n2151 gnd 0.006183f
C3202 vdd.n2152 gnd 0.006183f
C3203 vdd.n2153 gnd 0.004774f
C3204 vdd.n2154 gnd 0.008836f
C3205 vdd.n2155 gnd 0.004501f
C3206 vdd.n2156 gnd 0.006183f
C3207 vdd.n2157 gnd 0.006183f
C3208 vdd.n2158 gnd 0.006183f
C3209 vdd.n2159 gnd 0.006183f
C3210 vdd.n2160 gnd 0.006183f
C3211 vdd.n2161 gnd 0.006183f
C3212 vdd.n2162 gnd 0.006183f
C3213 vdd.n2163 gnd 0.006183f
C3214 vdd.n2164 gnd 0.006183f
C3215 vdd.n2165 gnd 0.006183f
C3216 vdd.n2166 gnd 0.006183f
C3217 vdd.n2167 gnd 0.006183f
C3218 vdd.n2168 gnd 0.006183f
C3219 vdd.n2169 gnd 0.006183f
C3220 vdd.n2170 gnd 0.006183f
C3221 vdd.n2171 gnd 0.006183f
C3222 vdd.n2172 gnd 0.006183f
C3223 vdd.n2173 gnd 0.006183f
C3224 vdd.n2174 gnd 0.006183f
C3225 vdd.n2175 gnd 0.006183f
C3226 vdd.n2176 gnd 0.006183f
C3227 vdd.n2177 gnd 0.006183f
C3228 vdd.n2178 gnd 0.006183f
C3229 vdd.n2179 gnd 0.006183f
C3230 vdd.n2180 gnd 0.006183f
C3231 vdd.n2181 gnd 0.006183f
C3232 vdd.n2182 gnd 0.006183f
C3233 vdd.n2183 gnd 0.006183f
C3234 vdd.n2184 gnd 0.006183f
C3235 vdd.n2185 gnd 0.006183f
C3236 vdd.n2186 gnd 0.006183f
C3237 vdd.n2187 gnd 0.006183f
C3238 vdd.n2188 gnd 0.006183f
C3239 vdd.n2189 gnd 0.006183f
C3240 vdd.n2190 gnd 0.006183f
C3241 vdd.n2191 gnd 0.006183f
C3242 vdd.n2192 gnd 0.006183f
C3243 vdd.n2193 gnd 0.006183f
C3244 vdd.n2194 gnd 0.006183f
C3245 vdd.n2195 gnd 0.006183f
C3246 vdd.n2196 gnd 0.006183f
C3247 vdd.n2197 gnd 0.006183f
C3248 vdd.n2198 gnd 0.006183f
C3249 vdd.n2199 gnd 0.006183f
C3250 vdd.n2200 gnd 0.006183f
C3251 vdd.n2201 gnd 0.006183f
C3252 vdd.n2202 gnd 0.006183f
C3253 vdd.n2203 gnd 0.006183f
C3254 vdd.n2204 gnd 0.006183f
C3255 vdd.n2205 gnd 0.006183f
C3256 vdd.n2206 gnd 0.006183f
C3257 vdd.n2207 gnd 0.006183f
C3258 vdd.n2208 gnd 0.006183f
C3259 vdd.n2209 gnd 0.006183f
C3260 vdd.n2210 gnd 0.006183f
C3261 vdd.n2211 gnd 0.006183f
C3262 vdd.n2212 gnd 0.006183f
C3263 vdd.n2213 gnd 0.006183f
C3264 vdd.n2214 gnd 0.006183f
C3265 vdd.n2215 gnd 0.006183f
C3266 vdd.n2216 gnd 0.014671f
C3267 vdd.n2217 gnd 0.014671f
C3268 vdd.n2218 gnd 0.771248f
C3269 vdd.t192 gnd 2.74118f
C3270 vdd.t98 gnd 2.74118f
C3271 vdd.n2251 gnd 0.014671f
C3272 vdd.n2252 gnd 0.006183f
C3273 vdd.t56 gnd 0.249851f
C3274 vdd.t57 gnd 0.255754f
C3275 vdd.t54 gnd 0.163112f
C3276 vdd.n2253 gnd 0.088153f
C3277 vdd.n2254 gnd 0.050003f
C3278 vdd.n2255 gnd 0.006183f
C3279 vdd.t70 gnd 0.249851f
C3280 vdd.t71 gnd 0.255754f
C3281 vdd.t69 gnd 0.163112f
C3282 vdd.n2256 gnd 0.088153f
C3283 vdd.n2257 gnd 0.050003f
C3284 vdd.n2258 gnd 0.008836f
C3285 vdd.n2259 gnd 0.006183f
C3286 vdd.n2260 gnd 0.006183f
C3287 vdd.n2261 gnd 0.006183f
C3288 vdd.n2262 gnd 0.006183f
C3289 vdd.n2263 gnd 0.006183f
C3290 vdd.n2264 gnd 0.006183f
C3291 vdd.n2265 gnd 0.006183f
C3292 vdd.n2266 gnd 0.006183f
C3293 vdd.n2267 gnd 0.006183f
C3294 vdd.n2268 gnd 0.006183f
C3295 vdd.n2269 gnd 0.006183f
C3296 vdd.n2270 gnd 0.006183f
C3297 vdd.n2271 gnd 0.006183f
C3298 vdd.n2272 gnd 0.006183f
C3299 vdd.n2273 gnd 0.006183f
C3300 vdd.n2274 gnd 0.006183f
C3301 vdd.n2275 gnd 0.006183f
C3302 vdd.n2276 gnd 0.006183f
C3303 vdd.n2277 gnd 0.006183f
C3304 vdd.n2278 gnd 0.006183f
C3305 vdd.n2279 gnd 0.006183f
C3306 vdd.n2280 gnd 0.006183f
C3307 vdd.n2281 gnd 0.006183f
C3308 vdd.n2282 gnd 0.006183f
C3309 vdd.n2283 gnd 0.006183f
C3310 vdd.n2284 gnd 0.006183f
C3311 vdd.n2285 gnd 0.006183f
C3312 vdd.n2286 gnd 0.006183f
C3313 vdd.n2287 gnd 0.006183f
C3314 vdd.n2288 gnd 0.006183f
C3315 vdd.n2289 gnd 0.006183f
C3316 vdd.n2290 gnd 0.006183f
C3317 vdd.n2291 gnd 0.006183f
C3318 vdd.n2292 gnd 0.006183f
C3319 vdd.n2293 gnd 0.006183f
C3320 vdd.n2294 gnd 0.006183f
C3321 vdd.n2295 gnd 0.006183f
C3322 vdd.n2296 gnd 0.006183f
C3323 vdd.n2297 gnd 0.006183f
C3324 vdd.n2298 gnd 0.006183f
C3325 vdd.n2299 gnd 0.006183f
C3326 vdd.n2300 gnd 0.006183f
C3327 vdd.n2301 gnd 0.006183f
C3328 vdd.n2302 gnd 0.006183f
C3329 vdd.n2303 gnd 0.006183f
C3330 vdd.n2304 gnd 0.006183f
C3331 vdd.n2305 gnd 0.006183f
C3332 vdd.n2306 gnd 0.006183f
C3333 vdd.n2307 gnd 0.006183f
C3334 vdd.n2308 gnd 0.006183f
C3335 vdd.n2309 gnd 0.006183f
C3336 vdd.n2310 gnd 0.006183f
C3337 vdd.n2311 gnd 0.006183f
C3338 vdd.n2312 gnd 0.006183f
C3339 vdd.n2313 gnd 0.006183f
C3340 vdd.n2314 gnd 0.006183f
C3341 vdd.n2315 gnd 0.004501f
C3342 vdd.n2316 gnd 0.006183f
C3343 vdd.n2317 gnd 0.006183f
C3344 vdd.n2318 gnd 0.004774f
C3345 vdd.n2319 gnd 0.006183f
C3346 vdd.n2320 gnd 0.006183f
C3347 vdd.n2321 gnd 0.014671f
C3348 vdd.n2322 gnd 0.013698f
C3349 vdd.n2323 gnd 0.006183f
C3350 vdd.n2324 gnd 0.006183f
C3351 vdd.n2325 gnd 0.006183f
C3352 vdd.n2326 gnd 0.006183f
C3353 vdd.n2327 gnd 0.006183f
C3354 vdd.n2328 gnd 0.006183f
C3355 vdd.n2329 gnd 0.006183f
C3356 vdd.n2330 gnd 0.006183f
C3357 vdd.n2331 gnd 0.006183f
C3358 vdd.n2332 gnd 0.006183f
C3359 vdd.n2333 gnd 0.006183f
C3360 vdd.n2334 gnd 0.006183f
C3361 vdd.n2335 gnd 0.006183f
C3362 vdd.n2336 gnd 0.006183f
C3363 vdd.n2337 gnd 0.006183f
C3364 vdd.n2338 gnd 0.006183f
C3365 vdd.n2339 gnd 0.006183f
C3366 vdd.n2340 gnd 0.006183f
C3367 vdd.n2341 gnd 0.006183f
C3368 vdd.n2342 gnd 0.006183f
C3369 vdd.n2343 gnd 0.006183f
C3370 vdd.n2344 gnd 0.006183f
C3371 vdd.n2345 gnd 0.006183f
C3372 vdd.n2346 gnd 0.006183f
C3373 vdd.n2347 gnd 0.006183f
C3374 vdd.n2348 gnd 0.006183f
C3375 vdd.n2349 gnd 0.006183f
C3376 vdd.n2350 gnd 0.006183f
C3377 vdd.n2351 gnd 0.006183f
C3378 vdd.n2352 gnd 0.006183f
C3379 vdd.n2353 gnd 0.006183f
C3380 vdd.n2354 gnd 0.006183f
C3381 vdd.n2355 gnd 0.006183f
C3382 vdd.n2356 gnd 0.006183f
C3383 vdd.n2357 gnd 0.006183f
C3384 vdd.n2358 gnd 0.006183f
C3385 vdd.n2359 gnd 0.006183f
C3386 vdd.n2360 gnd 0.006183f
C3387 vdd.n2361 gnd 0.006183f
C3388 vdd.n2362 gnd 0.006183f
C3389 vdd.n2363 gnd 0.006183f
C3390 vdd.n2364 gnd 0.006183f
C3391 vdd.n2365 gnd 0.006183f
C3392 vdd.n2366 gnd 0.006183f
C3393 vdd.n2367 gnd 0.006183f
C3394 vdd.n2368 gnd 0.006183f
C3395 vdd.n2369 gnd 0.006183f
C3396 vdd.n2370 gnd 0.006183f
C3397 vdd.n2371 gnd 0.006183f
C3398 vdd.n2372 gnd 0.006183f
C3399 vdd.n2373 gnd 0.006183f
C3400 vdd.n2374 gnd 0.199781f
C3401 vdd.n2375 gnd 0.006183f
C3402 vdd.n2376 gnd 0.006183f
C3403 vdd.n2377 gnd 0.006183f
C3404 vdd.n2378 gnd 0.006183f
C3405 vdd.n2379 gnd 0.006183f
C3406 vdd.n2380 gnd 0.006183f
C3407 vdd.n2381 gnd 0.006183f
C3408 vdd.n2382 gnd 0.006183f
C3409 vdd.n2383 gnd 0.006183f
C3410 vdd.n2384 gnd 0.006183f
C3411 vdd.n2385 gnd 0.006183f
C3412 vdd.n2386 gnd 0.006183f
C3413 vdd.n2387 gnd 0.006183f
C3414 vdd.n2388 gnd 0.006183f
C3415 vdd.n2389 gnd 0.006183f
C3416 vdd.n2390 gnd 0.006183f
C3417 vdd.n2391 gnd 0.006183f
C3418 vdd.n2392 gnd 0.006183f
C3419 vdd.n2393 gnd 0.006183f
C3420 vdd.n2394 gnd 0.006183f
C3421 vdd.n2395 gnd 0.376332f
C3422 vdd.n2396 gnd 0.006183f
C3423 vdd.n2397 gnd 0.006183f
C3424 vdd.n2398 gnd 0.006183f
C3425 vdd.n2399 gnd 0.006183f
C3426 vdd.n2400 gnd 0.006183f
C3427 vdd.n2401 gnd 0.013698f
C3428 vdd.n2402 gnd 0.014671f
C3429 vdd.n2403 gnd 0.014671f
C3430 vdd.n2404 gnd 0.006183f
C3431 vdd.n2405 gnd 0.006183f
C3432 vdd.n2406 gnd 0.006183f
C3433 vdd.n2407 gnd 0.004774f
C3434 vdd.n2408 gnd 0.008836f
C3435 vdd.n2409 gnd 0.004501f
C3436 vdd.n2410 gnd 0.006183f
C3437 vdd.n2411 gnd 0.006183f
C3438 vdd.n2412 gnd 0.006183f
C3439 vdd.n2413 gnd 0.006183f
C3440 vdd.n2414 gnd 0.006183f
C3441 vdd.n2415 gnd 0.006183f
C3442 vdd.n2416 gnd 0.006183f
C3443 vdd.n2417 gnd 0.006183f
C3444 vdd.n2418 gnd 0.006183f
C3445 vdd.n2419 gnd 0.006183f
C3446 vdd.n2420 gnd 0.006183f
C3447 vdd.n2421 gnd 0.006183f
C3448 vdd.n2422 gnd 0.006183f
C3449 vdd.n2423 gnd 0.006183f
C3450 vdd.n2424 gnd 0.006183f
C3451 vdd.n2425 gnd 0.006183f
C3452 vdd.n2426 gnd 0.006183f
C3453 vdd.n2427 gnd 0.006183f
C3454 vdd.n2428 gnd 0.006183f
C3455 vdd.n2429 gnd 0.006183f
C3456 vdd.n2430 gnd 0.006183f
C3457 vdd.n2431 gnd 0.006183f
C3458 vdd.n2432 gnd 0.006183f
C3459 vdd.n2433 gnd 0.006183f
C3460 vdd.n2434 gnd 0.006183f
C3461 vdd.n2435 gnd 0.006183f
C3462 vdd.n2436 gnd 0.006183f
C3463 vdd.n2437 gnd 0.006183f
C3464 vdd.n2438 gnd 0.006183f
C3465 vdd.n2439 gnd 0.006183f
C3466 vdd.n2440 gnd 0.006183f
C3467 vdd.n2441 gnd 0.006183f
C3468 vdd.n2442 gnd 0.006183f
C3469 vdd.n2443 gnd 0.006183f
C3470 vdd.n2444 gnd 0.006183f
C3471 vdd.n2445 gnd 0.006183f
C3472 vdd.n2446 gnd 0.006183f
C3473 vdd.n2447 gnd 0.006183f
C3474 vdd.n2448 gnd 0.006183f
C3475 vdd.n2449 gnd 0.006183f
C3476 vdd.n2450 gnd 0.006183f
C3477 vdd.n2451 gnd 0.006183f
C3478 vdd.n2452 gnd 0.006183f
C3479 vdd.n2453 gnd 0.006183f
C3480 vdd.n2454 gnd 0.006183f
C3481 vdd.n2455 gnd 0.006183f
C3482 vdd.n2456 gnd 0.006183f
C3483 vdd.n2457 gnd 0.006183f
C3484 vdd.n2458 gnd 0.006183f
C3485 vdd.n2459 gnd 0.006183f
C3486 vdd.n2460 gnd 0.006183f
C3487 vdd.n2461 gnd 0.006183f
C3488 vdd.n2462 gnd 0.006183f
C3489 vdd.n2463 gnd 0.006183f
C3490 vdd.n2464 gnd 0.006183f
C3491 vdd.n2465 gnd 0.006183f
C3492 vdd.n2466 gnd 0.006183f
C3493 vdd.n2467 gnd 0.006183f
C3494 vdd.n2468 gnd 0.006183f
C3495 vdd.n2469 gnd 0.006183f
C3496 vdd.n2471 gnd 0.771248f
C3497 vdd.n2473 gnd 0.006183f
C3498 vdd.n2474 gnd 0.006183f
C3499 vdd.n2475 gnd 0.014671f
C3500 vdd.n2476 gnd 0.013698f
C3501 vdd.n2477 gnd 0.013698f
C3502 vdd.n2478 gnd 0.771248f
C3503 vdd.n2479 gnd 0.013698f
C3504 vdd.n2480 gnd 0.013698f
C3505 vdd.n2481 gnd 0.006183f
C3506 vdd.n2482 gnd 0.006183f
C3507 vdd.n2483 gnd 0.006183f
C3508 vdd.n2484 gnd 0.394916f
C3509 vdd.n2485 gnd 0.006183f
C3510 vdd.n2486 gnd 0.006183f
C3511 vdd.n2487 gnd 0.006183f
C3512 vdd.n2488 gnd 0.006183f
C3513 vdd.n2489 gnd 0.006183f
C3514 vdd.n2490 gnd 0.492483f
C3515 vdd.n2491 gnd 0.006183f
C3516 vdd.n2492 gnd 0.006183f
C3517 vdd.n2493 gnd 0.006183f
C3518 vdd.n2494 gnd 0.006183f
C3519 vdd.n2495 gnd 0.006183f
C3520 vdd.n2496 gnd 0.631866f
C3521 vdd.n2497 gnd 0.006183f
C3522 vdd.n2498 gnd 0.006183f
C3523 vdd.n2499 gnd 0.006183f
C3524 vdd.n2500 gnd 0.006183f
C3525 vdd.n2501 gnd 0.006183f
C3526 vdd.n2502 gnd 0.348455f
C3527 vdd.n2503 gnd 0.006183f
C3528 vdd.n2504 gnd 0.006183f
C3529 vdd.n2505 gnd 0.006183f
C3530 vdd.n2506 gnd 0.006183f
C3531 vdd.n2507 gnd 0.006183f
C3532 vdd.n2508 gnd 0.199781f
C3533 vdd.n2509 gnd 0.006183f
C3534 vdd.n2510 gnd 0.006183f
C3535 vdd.n2511 gnd 0.006183f
C3536 vdd.n2512 gnd 0.006183f
C3537 vdd.n2513 gnd 0.006183f
C3538 vdd.n2514 gnd 0.362393f
C3539 vdd.n2515 gnd 0.006183f
C3540 vdd.n2516 gnd 0.006183f
C3541 vdd.n2517 gnd 0.006183f
C3542 vdd.n2518 gnd 0.006183f
C3543 vdd.n2519 gnd 0.006183f
C3544 vdd.n2520 gnd 0.501776f
C3545 vdd.n2521 gnd 0.006183f
C3546 vdd.n2522 gnd 0.006183f
C3547 vdd.n2523 gnd 0.006183f
C3548 vdd.n2524 gnd 0.006183f
C3549 vdd.n2525 gnd 0.006183f
C3550 vdd.n2526 gnd 0.562174f
C3551 vdd.n2527 gnd 0.006183f
C3552 vdd.n2528 gnd 0.006183f
C3553 vdd.n2529 gnd 0.006183f
C3554 vdd.n2530 gnd 0.006183f
C3555 vdd.n2531 gnd 0.006183f
C3556 vdd.n2532 gnd 0.422792f
C3557 vdd.n2533 gnd 0.006183f
C3558 vdd.n2534 gnd 0.006183f
C3559 vdd.n2535 gnd 0.006183f
C3560 vdd.t31 gnd 0.255754f
C3561 vdd.t29 gnd 0.163112f
C3562 vdd.t32 gnd 0.255754f
C3563 vdd.n2536 gnd 0.143744f
C3564 vdd.n2537 gnd 0.017911f
C3565 vdd.n2538 gnd 0.003819f
C3566 vdd.n2539 gnd 0.006183f
C3567 vdd.n2540 gnd 0.348455f
C3568 vdd.n2541 gnd 0.006183f
C3569 vdd.n2542 gnd 0.006183f
C3570 vdd.n2543 gnd 0.006183f
C3571 vdd.n2544 gnd 0.006183f
C3572 vdd.n2545 gnd 0.006183f
C3573 vdd.n2546 gnd 0.631866f
C3574 vdd.n2547 gnd 0.006183f
C3575 vdd.n2548 gnd 0.006183f
C3576 vdd.n2549 gnd 0.006183f
C3577 vdd.n2550 gnd 0.006183f
C3578 vdd.n2551 gnd 0.006183f
C3579 vdd.n2552 gnd 0.006183f
C3580 vdd.n2554 gnd 0.006183f
C3581 vdd.n2555 gnd 0.006183f
C3582 vdd.n2557 gnd 0.006183f
C3583 vdd.n2558 gnd 0.006183f
C3584 vdd.n2561 gnd 0.006183f
C3585 vdd.n2562 gnd 0.006183f
C3586 vdd.n2563 gnd 0.006183f
C3587 vdd.n2564 gnd 0.006183f
C3588 vdd.n2566 gnd 0.006183f
C3589 vdd.n2567 gnd 0.006183f
C3590 vdd.n2568 gnd 0.006183f
C3591 vdd.n2569 gnd 0.006183f
C3592 vdd.n2570 gnd 0.006183f
C3593 vdd.n2571 gnd 0.006183f
C3594 vdd.n2573 gnd 0.006183f
C3595 vdd.n2574 gnd 0.006183f
C3596 vdd.n2575 gnd 0.006183f
C3597 vdd.n2576 gnd 0.006183f
C3598 vdd.n2577 gnd 0.006183f
C3599 vdd.n2578 gnd 0.006183f
C3600 vdd.n2580 gnd 0.006183f
C3601 vdd.n2581 gnd 0.006183f
C3602 vdd.n2582 gnd 0.006183f
C3603 vdd.n2583 gnd 0.006183f
C3604 vdd.n2584 gnd 0.006183f
C3605 vdd.n2585 gnd 0.006183f
C3606 vdd.n2587 gnd 0.006183f
C3607 vdd.n2588 gnd 0.014671f
C3608 vdd.n2589 gnd 0.014671f
C3609 vdd.n2590 gnd 0.013698f
C3610 vdd.n2591 gnd 0.006183f
C3611 vdd.n2592 gnd 0.006183f
C3612 vdd.n2593 gnd 0.006183f
C3613 vdd.n2594 gnd 0.006183f
C3614 vdd.n2595 gnd 0.006183f
C3615 vdd.n2596 gnd 0.006183f
C3616 vdd.n2597 gnd 0.631866f
C3617 vdd.n2598 gnd 0.006183f
C3618 vdd.n2599 gnd 0.006183f
C3619 vdd.n2600 gnd 0.006183f
C3620 vdd.n2601 gnd 0.006183f
C3621 vdd.n2602 gnd 0.006183f
C3622 vdd.n2603 gnd 0.394916f
C3623 vdd.n2604 gnd 0.006183f
C3624 vdd.n2605 gnd 0.006183f
C3625 vdd.n2606 gnd 0.006183f
C3626 vdd.n2607 gnd 0.014451f
C3627 vdd.n2608 gnd 0.013918f
C3628 vdd.n2609 gnd 0.014671f
C3629 vdd.n2611 gnd 0.006183f
C3630 vdd.n2612 gnd 0.006183f
C3631 vdd.n2613 gnd 0.004774f
C3632 vdd.n2614 gnd 0.008836f
C3633 vdd.n2615 gnd 0.004501f
C3634 vdd.n2616 gnd 0.006183f
C3635 vdd.n2617 gnd 0.006183f
C3636 vdd.n2619 gnd 0.006183f
C3637 vdd.n2620 gnd 0.006183f
C3638 vdd.n2621 gnd 0.006183f
C3639 vdd.n2622 gnd 0.006183f
C3640 vdd.n2623 gnd 0.006183f
C3641 vdd.n2624 gnd 0.006183f
C3642 vdd.n2626 gnd 0.006183f
C3643 vdd.n2627 gnd 0.006183f
C3644 vdd.n2628 gnd 0.006183f
C3645 vdd.n2629 gnd 0.006183f
C3646 vdd.n2630 gnd 0.006183f
C3647 vdd.n2631 gnd 0.006183f
C3648 vdd.n2633 gnd 0.006183f
C3649 vdd.n2634 gnd 0.006183f
C3650 vdd.n2635 gnd 0.006183f
C3651 vdd.n2636 gnd 0.006183f
C3652 vdd.n2637 gnd 0.006183f
C3653 vdd.n2638 gnd 0.006183f
C3654 vdd.n2640 gnd 0.006183f
C3655 vdd.n2641 gnd 0.006183f
C3656 vdd.n2642 gnd 0.006183f
C3657 vdd.n2644 gnd 0.006183f
C3658 vdd.n2645 gnd 0.006183f
C3659 vdd.n2646 gnd 0.006183f
C3660 vdd.n2647 gnd 0.006183f
C3661 vdd.n2648 gnd 0.006183f
C3662 vdd.n2649 gnd 0.006183f
C3663 vdd.n2651 gnd 0.006183f
C3664 vdd.n2652 gnd 0.006183f
C3665 vdd.n2653 gnd 0.006183f
C3666 vdd.n2654 gnd 0.006183f
C3667 vdd.n2655 gnd 0.006183f
C3668 vdd.n2656 gnd 0.006183f
C3669 vdd.n2658 gnd 0.006183f
C3670 vdd.n2659 gnd 0.006183f
C3671 vdd.n2660 gnd 0.006183f
C3672 vdd.n2661 gnd 0.006183f
C3673 vdd.n2662 gnd 0.006183f
C3674 vdd.n2663 gnd 0.006183f
C3675 vdd.n2665 gnd 0.006183f
C3676 vdd.n2666 gnd 0.006183f
C3677 vdd.n2668 gnd 0.006183f
C3678 vdd.n2669 gnd 0.006183f
C3679 vdd.n2670 gnd 0.014671f
C3680 vdd.n2671 gnd 0.013698f
C3681 vdd.n2672 gnd 0.013698f
C3682 vdd.n2673 gnd 0.91063f
C3683 vdd.n2674 gnd 0.013698f
C3684 vdd.n2675 gnd 0.014671f
C3685 vdd.n2676 gnd 0.013918f
C3686 vdd.n2677 gnd 0.006183f
C3687 vdd.n2678 gnd 0.004774f
C3688 vdd.n2679 gnd 0.006183f
C3689 vdd.n2681 gnd 0.006183f
C3690 vdd.n2682 gnd 0.006183f
C3691 vdd.n2683 gnd 0.006183f
C3692 vdd.n2684 gnd 0.006183f
C3693 vdd.n2685 gnd 0.006183f
C3694 vdd.n2686 gnd 0.006183f
C3695 vdd.n2688 gnd 0.006183f
C3696 vdd.n2689 gnd 0.006183f
C3697 vdd.n2690 gnd 0.006183f
C3698 vdd.n2691 gnd 0.006183f
C3699 vdd.n2692 gnd 0.006183f
C3700 vdd.n2693 gnd 0.006183f
C3701 vdd.n2695 gnd 0.006183f
C3702 vdd.n2696 gnd 0.006183f
C3703 vdd.n2697 gnd 0.006183f
C3704 vdd.n2698 gnd 0.006183f
C3705 vdd.n2699 gnd 0.006183f
C3706 vdd.n2700 gnd 0.006183f
C3707 vdd.n2702 gnd 0.006183f
C3708 vdd.n2703 gnd 0.006183f
C3709 vdd.n2705 gnd 0.006183f
C3710 vdd.n2706 gnd 0.014858f
C3711 vdd.n2707 gnd 0.550295f
C3712 vdd.n2708 gnd 0.00782f
C3713 vdd.n2709 gnd 0.022667f
C3714 vdd.n2710 gnd 0.003476f
C3715 vdd.t82 gnd 0.111862f
C3716 vdd.t83 gnd 0.11955f
C3717 vdd.t81 gnd 0.14609f
C3718 vdd.n2711 gnd 0.187267f
C3719 vdd.n2712 gnd 0.157338f
C3720 vdd.n2713 gnd 0.01127f
C3721 vdd.n2714 gnd 0.009093f
C3722 vdd.n2715 gnd 0.003842f
C3723 vdd.n2716 gnd 0.007318f
C3724 vdd.n2717 gnd 0.009093f
C3725 vdd.n2718 gnd 0.009093f
C3726 vdd.n2719 gnd 0.007318f
C3727 vdd.n2720 gnd 0.007318f
C3728 vdd.n2721 gnd 0.009093f
C3729 vdd.n2722 gnd 0.009093f
C3730 vdd.n2723 gnd 0.007318f
C3731 vdd.n2724 gnd 0.007318f
C3732 vdd.n2725 gnd 0.009093f
C3733 vdd.n2726 gnd 0.009093f
C3734 vdd.n2727 gnd 0.007318f
C3735 vdd.n2728 gnd 0.007318f
C3736 vdd.n2729 gnd 0.009093f
C3737 vdd.n2730 gnd 0.009093f
C3738 vdd.n2731 gnd 0.007318f
C3739 vdd.n2732 gnd 0.007318f
C3740 vdd.n2733 gnd 0.009093f
C3741 vdd.n2734 gnd 0.009093f
C3742 vdd.n2735 gnd 0.007318f
C3743 vdd.n2736 gnd 0.007318f
C3744 vdd.n2737 gnd 0.009093f
C3745 vdd.n2738 gnd 0.009093f
C3746 vdd.n2739 gnd 0.007318f
C3747 vdd.n2740 gnd 0.007318f
C3748 vdd.n2741 gnd 0.009093f
C3749 vdd.n2742 gnd 0.009093f
C3750 vdd.n2743 gnd 0.007318f
C3751 vdd.n2744 gnd 0.007318f
C3752 vdd.n2745 gnd 0.009093f
C3753 vdd.n2746 gnd 0.009093f
C3754 vdd.n2747 gnd 0.007318f
C3755 vdd.n2748 gnd 0.007318f
C3756 vdd.n2749 gnd 0.009093f
C3757 vdd.n2750 gnd 0.009093f
C3758 vdd.n2751 gnd 0.007318f
C3759 vdd.n2752 gnd 0.009093f
C3760 vdd.n2753 gnd 0.009093f
C3761 vdd.n2754 gnd 0.007318f
C3762 vdd.n2755 gnd 0.009093f
C3763 vdd.n2756 gnd 0.009093f
C3764 vdd.n2757 gnd 0.009093f
C3765 vdd.n2758 gnd 0.01493f
C3766 vdd.n2759 gnd 0.009093f
C3767 vdd.n2760 gnd 0.009093f
C3768 vdd.n2761 gnd 0.004977f
C3769 vdd.n2762 gnd 0.007318f
C3770 vdd.n2763 gnd 0.009093f
C3771 vdd.n2764 gnd 0.009093f
C3772 vdd.n2765 gnd 0.007318f
C3773 vdd.n2766 gnd 0.007318f
C3774 vdd.n2767 gnd 0.009093f
C3775 vdd.n2768 gnd 0.009093f
C3776 vdd.n2769 gnd 0.007318f
C3777 vdd.n2770 gnd 0.007318f
C3778 vdd.n2771 gnd 0.009093f
C3779 vdd.n2772 gnd 0.009093f
C3780 vdd.n2773 gnd 0.007318f
C3781 vdd.n2774 gnd 0.007318f
C3782 vdd.n2775 gnd 0.009093f
C3783 vdd.n2776 gnd 0.009093f
C3784 vdd.n2777 gnd 0.007318f
C3785 vdd.n2778 gnd 0.007318f
C3786 vdd.n2779 gnd 0.009093f
C3787 vdd.n2780 gnd 0.009093f
C3788 vdd.n2781 gnd 0.007318f
C3789 vdd.n2782 gnd 0.007318f
C3790 vdd.n2783 gnd 0.009093f
C3791 vdd.n2784 gnd 0.009093f
C3792 vdd.n2785 gnd 0.007318f
C3793 vdd.n2786 gnd 0.007318f
C3794 vdd.n2787 gnd 0.009093f
C3795 vdd.n2788 gnd 0.009093f
C3796 vdd.n2789 gnd 0.007318f
C3797 vdd.n2790 gnd 0.007318f
C3798 vdd.n2791 gnd 0.009093f
C3799 vdd.n2792 gnd 0.009093f
C3800 vdd.n2793 gnd 0.007318f
C3801 vdd.n2794 gnd 0.007318f
C3802 vdd.n2795 gnd 0.009093f
C3803 vdd.n2796 gnd 0.009093f
C3804 vdd.n2797 gnd 0.007318f
C3805 vdd.n2798 gnd 0.009093f
C3806 vdd.n2799 gnd 0.009093f
C3807 vdd.n2800 gnd 0.007318f
C3808 vdd.n2801 gnd 0.009093f
C3809 vdd.n2802 gnd 0.009093f
C3810 vdd.n2803 gnd 0.009093f
C3811 vdd.t19 gnd 0.111862f
C3812 vdd.t20 gnd 0.11955f
C3813 vdd.t18 gnd 0.14609f
C3814 vdd.n2804 gnd 0.187267f
C3815 vdd.n2805 gnd 0.157338f
C3816 vdd.n2806 gnd 0.01493f
C3817 vdd.n2807 gnd 0.009093f
C3818 vdd.n2808 gnd 0.009093f
C3819 vdd.n2809 gnd 0.006111f
C3820 vdd.n2810 gnd 0.007318f
C3821 vdd.n2811 gnd 0.009093f
C3822 vdd.n2812 gnd 0.009093f
C3823 vdd.n2813 gnd 0.007318f
C3824 vdd.n2814 gnd 0.007318f
C3825 vdd.n2815 gnd 0.009093f
C3826 vdd.n2816 gnd 0.009093f
C3827 vdd.n2817 gnd 0.007318f
C3828 vdd.n2818 gnd 0.007318f
C3829 vdd.n2819 gnd 0.009093f
C3830 vdd.n2820 gnd 0.009093f
C3831 vdd.n2821 gnd 0.007318f
C3832 vdd.n2822 gnd 0.007318f
C3833 vdd.n2823 gnd 0.009093f
C3834 vdd.n2824 gnd 0.009093f
C3835 vdd.n2825 gnd 0.007318f
C3836 vdd.n2826 gnd 0.007318f
C3837 vdd.n2827 gnd 0.009093f
C3838 vdd.n2828 gnd 0.009093f
C3839 vdd.n2829 gnd 0.007318f
C3840 vdd.n2830 gnd 0.007318f
C3841 vdd.n2831 gnd 0.009093f
C3842 vdd.n2832 gnd 0.009093f
C3843 vdd.n2833 gnd 0.007318f
C3844 vdd.n2834 gnd 0.007318f
C3845 vdd.n2836 gnd 0.550295f
C3846 vdd.n2838 gnd 0.007318f
C3847 vdd.n2839 gnd 0.009093f
C3848 vdd.n2840 gnd 6.7368f
C3849 vdd.n2842 gnd 0.022667f
C3850 vdd.n2843 gnd 0.006074f
C3851 vdd.n2844 gnd 0.022667f
C3852 vdd.n2845 gnd 0.022159f
C3853 vdd.n2846 gnd 0.009093f
C3854 vdd.n2847 gnd 0.007318f
C3855 vdd.n2848 gnd 0.009093f
C3856 vdd.n2849 gnd 0.580759f
C3857 vdd.n2850 gnd 0.009093f
C3858 vdd.n2851 gnd 0.007318f
C3859 vdd.n2852 gnd 0.009093f
C3860 vdd.n2853 gnd 0.009093f
C3861 vdd.n2854 gnd 0.009093f
C3862 vdd.n2855 gnd 0.007318f
C3863 vdd.n2856 gnd 0.009093f
C3864 vdd.n2857 gnd 0.738725f
C3865 vdd.n2858 gnd 0.929214f
C3866 vdd.n2859 gnd 0.009093f
C3867 vdd.n2860 gnd 0.007318f
C3868 vdd.n2861 gnd 0.009093f
C3869 vdd.n2862 gnd 0.009093f
C3870 vdd.n2863 gnd 0.009093f
C3871 vdd.n2864 gnd 0.007318f
C3872 vdd.n2865 gnd 0.009093f
C3873 vdd.n2866 gnd 0.655096f
C3874 vdd.n2867 gnd 0.009093f
C3875 vdd.n2868 gnd 0.007318f
C3876 vdd.n2869 gnd 0.009093f
C3877 vdd.n2870 gnd 0.009093f
C3878 vdd.n2871 gnd 0.009093f
C3879 vdd.n2872 gnd 0.007318f
C3880 vdd.n2873 gnd 0.009093f
C3881 vdd.t140 gnd 0.464607f
C3882 vdd.n2874 gnd 0.771248f
C3883 vdd.n2875 gnd 0.009093f
C3884 vdd.n2876 gnd 0.007318f
C3885 vdd.n2877 gnd 0.009093f
C3886 vdd.n2878 gnd 0.009093f
C3887 vdd.n2879 gnd 0.009093f
C3888 vdd.n2880 gnd 0.007318f
C3889 vdd.n2881 gnd 0.009093f
C3890 vdd.n2882 gnd 0.729433f
C3891 vdd.n2883 gnd 0.009093f
C3892 vdd.n2884 gnd 0.007318f
C3893 vdd.n2885 gnd 0.009093f
C3894 vdd.n2886 gnd 0.009093f
C3895 vdd.n2887 gnd 0.009093f
C3896 vdd.n2888 gnd 0.007318f
C3897 vdd.n2889 gnd 0.007318f
C3898 vdd.n2890 gnd 0.007318f
C3899 vdd.n2891 gnd 0.009093f
C3900 vdd.n2892 gnd 0.009093f
C3901 vdd.n2893 gnd 0.009093f
C3902 vdd.n2894 gnd 0.007318f
C3903 vdd.n2895 gnd 0.007318f
C3904 vdd.n2896 gnd 0.007318f
C3905 vdd.n2897 gnd 0.009093f
C3906 vdd.n2898 gnd 0.009093f
C3907 vdd.n2899 gnd 0.009093f
C3908 vdd.n2900 gnd 0.007318f
C3909 vdd.n2901 gnd 0.007318f
C3910 vdd.n2902 gnd 0.006074f
C3911 vdd.n2903 gnd 0.022159f
C3912 vdd.n2904 gnd 0.022667f
C3913 vdd.n2906 gnd 0.022667f
C3914 vdd.n2907 gnd 0.003476f
C3915 vdd.t86 gnd 0.111862f
C3916 vdd.t85 gnd 0.11955f
C3917 vdd.t84 gnd 0.14609f
C3918 vdd.n2908 gnd 0.187267f
C3919 vdd.n2909 gnd 0.15807f
C3920 vdd.n2910 gnd 0.012002f
C3921 vdd.n2911 gnd 0.003842f
C3922 vdd.n2912 gnd 0.007318f
C3923 vdd.n2913 gnd 0.009093f
C3924 vdd.n2915 gnd 0.009093f
C3925 vdd.n2916 gnd 0.009093f
C3926 vdd.n2917 gnd 0.007318f
C3927 vdd.n2918 gnd 0.007318f
C3928 vdd.n2919 gnd 0.007318f
C3929 vdd.n2920 gnd 0.009093f
C3930 vdd.n2922 gnd 0.009093f
C3931 vdd.n2923 gnd 0.009093f
C3932 vdd.n2924 gnd 0.007318f
C3933 vdd.n2925 gnd 0.007318f
C3934 vdd.n2926 gnd 0.007318f
C3935 vdd.n2927 gnd 0.009093f
C3936 vdd.n2929 gnd 0.009093f
C3937 vdd.n2930 gnd 0.009093f
C3938 vdd.n2931 gnd 0.007318f
C3939 vdd.n2932 gnd 0.007318f
C3940 vdd.n2933 gnd 0.007318f
C3941 vdd.n2934 gnd 0.009093f
C3942 vdd.n2936 gnd 0.009093f
C3943 vdd.n2937 gnd 0.009093f
C3944 vdd.n2938 gnd 0.007318f
C3945 vdd.n2939 gnd 0.007318f
C3946 vdd.n2940 gnd 0.007318f
C3947 vdd.n2941 gnd 0.009093f
C3948 vdd.n2943 gnd 0.009093f
C3949 vdd.n2944 gnd 0.009093f
C3950 vdd.n2945 gnd 0.007318f
C3951 vdd.n2946 gnd 0.009093f
C3952 vdd.n2947 gnd 0.009093f
C3953 vdd.n2948 gnd 0.009093f
C3954 vdd.n2949 gnd 0.015661f
C3955 vdd.n2950 gnd 0.004977f
C3956 vdd.n2951 gnd 0.007318f
C3957 vdd.n2952 gnd 0.009093f
C3958 vdd.n2954 gnd 0.009093f
C3959 vdd.n2955 gnd 0.009093f
C3960 vdd.n2956 gnd 0.007318f
C3961 vdd.n2957 gnd 0.007318f
C3962 vdd.n2958 gnd 0.007318f
C3963 vdd.n2959 gnd 0.009093f
C3964 vdd.n2961 gnd 0.009093f
C3965 vdd.n2962 gnd 0.009093f
C3966 vdd.n2963 gnd 0.007318f
C3967 vdd.n2964 gnd 0.007318f
C3968 vdd.n2965 gnd 0.007318f
C3969 vdd.n2966 gnd 0.009093f
C3970 vdd.n2968 gnd 0.009093f
C3971 vdd.n2969 gnd 0.009093f
C3972 vdd.n2970 gnd 0.007318f
C3973 vdd.n2971 gnd 0.007318f
C3974 vdd.n2972 gnd 0.007318f
C3975 vdd.n2973 gnd 0.009093f
C3976 vdd.n2975 gnd 0.009093f
C3977 vdd.n2976 gnd 0.009093f
C3978 vdd.n2977 gnd 0.007318f
C3979 vdd.n2978 gnd 0.007318f
C3980 vdd.n2979 gnd 0.007318f
C3981 vdd.n2980 gnd 0.009093f
C3982 vdd.n2982 gnd 0.009093f
C3983 vdd.n2983 gnd 0.009093f
C3984 vdd.n2984 gnd 0.007318f
C3985 vdd.n2985 gnd 0.009093f
C3986 vdd.n2986 gnd 0.009093f
C3987 vdd.n2987 gnd 0.009093f
C3988 vdd.n2988 gnd 0.015661f
C3989 vdd.n2989 gnd 0.006111f
C3990 vdd.n2990 gnd 0.007318f
C3991 vdd.n2991 gnd 0.009093f
C3992 vdd.n2993 gnd 0.009093f
C3993 vdd.n2994 gnd 0.009093f
C3994 vdd.n2995 gnd 0.007318f
C3995 vdd.n2996 gnd 0.007318f
C3996 vdd.n2997 gnd 0.007318f
C3997 vdd.n2998 gnd 0.009093f
C3998 vdd.n3000 gnd 0.009093f
C3999 vdd.n3001 gnd 0.009093f
C4000 vdd.n3002 gnd 0.007318f
C4001 vdd.n3003 gnd 0.007318f
C4002 vdd.n3004 gnd 0.007318f
C4003 vdd.n3005 gnd 0.009093f
C4004 vdd.n3007 gnd 0.009093f
C4005 vdd.n3008 gnd 0.009093f
C4006 vdd.n3009 gnd 0.007318f
C4007 vdd.n3010 gnd 0.007318f
C4008 vdd.n3011 gnd 0.007318f
C4009 vdd.n3012 gnd 0.009093f
C4010 vdd.n3014 gnd 0.009093f
C4011 vdd.n3015 gnd 0.009093f
C4012 vdd.n3017 gnd 0.009093f
C4013 vdd.n3018 gnd 0.007318f
C4014 vdd.n3019 gnd 0.007318f
C4015 vdd.n3020 gnd 0.006074f
C4016 vdd.n3021 gnd 0.022667f
C4017 vdd.n3022 gnd 0.022159f
C4018 vdd.n3023 gnd 0.006074f
C4019 vdd.n3024 gnd 0.022159f
C4020 vdd.n3025 gnd 1.37059f
C4021 vdd.t37 gnd 0.464607f
C4022 vdd.n3026 gnd 0.487837f
C4023 vdd.n3027 gnd 0.929214f
C4024 vdd.n3028 gnd 0.009093f
C4025 vdd.n3029 gnd 0.007318f
C4026 vdd.n3030 gnd 0.007318f
C4027 vdd.n3031 gnd 0.007318f
C4028 vdd.n3032 gnd 0.009093f
C4029 vdd.n3033 gnd 0.831647f
C4030 vdd.t131 gnd 0.464607f
C4031 vdd.n3034 gnd 0.562174f
C4032 vdd.n3035 gnd 0.67368f
C4033 vdd.n3036 gnd 0.009093f
C4034 vdd.n3037 gnd 0.007318f
C4035 vdd.n3038 gnd 0.007318f
C4036 vdd.n3039 gnd 0.007318f
C4037 vdd.n3040 gnd 0.009093f
C4038 vdd.n3041 gnd 0.515714f
C4039 vdd.t153 gnd 0.464607f
C4040 vdd.n3042 gnd 0.771248f
C4041 vdd.t129 gnd 0.464607f
C4042 vdd.n3043 gnd 0.571467f
C4043 vdd.n3044 gnd 0.009093f
C4044 vdd.n3045 gnd 0.007318f
C4045 vdd.n3046 gnd 0.006988f
C4046 vdd.n3047 gnd 0.536312f
C4047 vdd.n3048 gnd 1.84155f
C4048 a_n5644_8799.n0 gnd 0.207505f
C4049 a_n5644_8799.n1 gnd 0.286067f
C4050 a_n5644_8799.n2 gnd 0.217042f
C4051 a_n5644_8799.n3 gnd 0.207505f
C4052 a_n5644_8799.n4 gnd 0.286067f
C4053 a_n5644_8799.n5 gnd 0.217042f
C4054 a_n5644_8799.n6 gnd 0.207505f
C4055 a_n5644_8799.n7 gnd 0.450816f
C4056 a_n5644_8799.n8 gnd 0.217042f
C4057 a_n5644_8799.n9 gnd 0.207505f
C4058 a_n5644_8799.n10 gnd 0.320795f
C4059 a_n5644_8799.n11 gnd 0.182314f
C4060 a_n5644_8799.n12 gnd 0.207505f
C4061 a_n5644_8799.n13 gnd 0.320795f
C4062 a_n5644_8799.n14 gnd 0.182314f
C4063 a_n5644_8799.n15 gnd 0.207505f
C4064 a_n5644_8799.n16 gnd 0.320795f
C4065 a_n5644_8799.n17 gnd 0.347064f
C4066 a_n5644_8799.n18 gnd 2.78717f
C4067 a_n5644_8799.n19 gnd 4.02361f
C4068 a_n5644_8799.n20 gnd 0.362739f
C4069 a_n5644_8799.n21 gnd 3.04009f
C4070 a_n5644_8799.n22 gnd 0.362738f
C4071 a_n5644_8799.n23 gnd 0.854944f
C4072 a_n5644_8799.n24 gnd 0.249816f
C4073 a_n5644_8799.n25 gnd 0.004664f
C4074 a_n5644_8799.n26 gnd 0.010087f
C4075 a_n5644_8799.n27 gnd 0.010087f
C4076 a_n5644_8799.n28 gnd 0.004664f
C4077 a_n5644_8799.n29 gnd 0.249816f
C4078 a_n5644_8799.n30 gnd 0.004664f
C4079 a_n5644_8799.n31 gnd 0.010087f
C4080 a_n5644_8799.n32 gnd 0.010087f
C4081 a_n5644_8799.n33 gnd 0.004664f
C4082 a_n5644_8799.n34 gnd 0.249816f
C4083 a_n5644_8799.n35 gnd 0.004664f
C4084 a_n5644_8799.n36 gnd 0.010087f
C4085 a_n5644_8799.n37 gnd 0.010087f
C4086 a_n5644_8799.n38 gnd 0.004664f
C4087 a_n5644_8799.n39 gnd 0.004664f
C4088 a_n5644_8799.n40 gnd 0.010087f
C4089 a_n5644_8799.n41 gnd 0.010087f
C4090 a_n5644_8799.n42 gnd 0.004664f
C4091 a_n5644_8799.n43 gnd 0.249816f
C4092 a_n5644_8799.n44 gnd 0.004664f
C4093 a_n5644_8799.n45 gnd 0.010087f
C4094 a_n5644_8799.n46 gnd 0.010087f
C4095 a_n5644_8799.n47 gnd 0.004664f
C4096 a_n5644_8799.n48 gnd 0.249816f
C4097 a_n5644_8799.n49 gnd 0.004664f
C4098 a_n5644_8799.n50 gnd 0.010087f
C4099 a_n5644_8799.n51 gnd 0.010087f
C4100 a_n5644_8799.n52 gnd 0.004664f
C4101 a_n5644_8799.n53 gnd 0.249816f
C4102 a_n5644_8799.t19 gnd 0.143928f
C4103 a_n5644_8799.t7 gnd 0.143928f
C4104 a_n5644_8799.t34 gnd 0.143928f
C4105 a_n5644_8799.n54 gnd 1.13518f
C4106 a_n5644_8799.t23 gnd 0.143928f
C4107 a_n5644_8799.t10 gnd 0.143928f
C4108 a_n5644_8799.n55 gnd 1.13331f
C4109 a_n5644_8799.t13 gnd 0.143928f
C4110 a_n5644_8799.t12 gnd 0.143928f
C4111 a_n5644_8799.n56 gnd 1.13331f
C4112 a_n5644_8799.t31 gnd 0.111944f
C4113 a_n5644_8799.t24 gnd 0.111944f
C4114 a_n5644_8799.n57 gnd 0.992092f
C4115 a_n5644_8799.t5 gnd 0.111944f
C4116 a_n5644_8799.t3 gnd 0.111944f
C4117 a_n5644_8799.n58 gnd 0.989175f
C4118 a_n5644_8799.n59 gnd 0.877149f
C4119 a_n5644_8799.t27 gnd 0.111944f
C4120 a_n5644_8799.t17 gnd 0.111944f
C4121 a_n5644_8799.n60 gnd 0.989175f
C4122 a_n5644_8799.t33 gnd 0.111944f
C4123 a_n5644_8799.t9 gnd 0.111944f
C4124 a_n5644_8799.n61 gnd 0.992091f
C4125 a_n5644_8799.t0 gnd 0.111944f
C4126 a_n5644_8799.t28 gnd 0.111944f
C4127 a_n5644_8799.n62 gnd 0.989174f
C4128 a_n5644_8799.n63 gnd 0.877151f
C4129 a_n5644_8799.t26 gnd 0.111944f
C4130 a_n5644_8799.t29 gnd 0.111944f
C4131 a_n5644_8799.n64 gnd 0.989174f
C4132 a_n5644_8799.t16 gnd 0.111944f
C4133 a_n5644_8799.t8 gnd 0.111944f
C4134 a_n5644_8799.n65 gnd 0.992091f
C4135 a_n5644_8799.t11 gnd 0.111944f
C4136 a_n5644_8799.t22 gnd 0.111944f
C4137 a_n5644_8799.n66 gnd 0.989174f
C4138 a_n5644_8799.n67 gnd 0.877151f
C4139 a_n5644_8799.t20 gnd 0.111944f
C4140 a_n5644_8799.t1 gnd 0.111944f
C4141 a_n5644_8799.n68 gnd 0.989174f
C4142 a_n5644_8799.t32 gnd 0.111944f
C4143 a_n5644_8799.t25 gnd 0.111944f
C4144 a_n5644_8799.n69 gnd 0.989175f
C4145 a_n5644_8799.n70 gnd 3.08572f
C4146 a_n5644_8799.t21 gnd 0.111944f
C4147 a_n5644_8799.t35 gnd 0.111944f
C4148 a_n5644_8799.n71 gnd 0.989175f
C4149 a_n5644_8799.n72 gnd 0.431882f
C4150 a_n5644_8799.t30 gnd 0.111944f
C4151 a_n5644_8799.t4 gnd 0.111944f
C4152 a_n5644_8799.n73 gnd 0.989175f
C4153 a_n5644_8799.t75 gnd 0.596792f
C4154 a_n5644_8799.n74 gnd 0.268224f
C4155 a_n5644_8799.t42 gnd 0.596792f
C4156 a_n5644_8799.t62 gnd 0.596792f
C4157 a_n5644_8799.t53 gnd 0.608087f
C4158 a_n5644_8799.n75 gnd 0.250184f
C4159 a_n5644_8799.n76 gnd 0.270608f
C4160 a_n5644_8799.t77 gnd 0.596792f
C4161 a_n5644_8799.n77 gnd 0.268224f
C4162 a_n5644_8799.n78 gnd 0.26382f
C4163 a_n5644_8799.t52 gnd 0.596792f
C4164 a_n5644_8799.n79 gnd 0.26382f
C4165 a_n5644_8799.t41 gnd 0.596792f
C4166 a_n5644_8799.n80 gnd 0.270608f
C4167 a_n5644_8799.t40 gnd 0.608077f
C4168 a_n5644_8799.t79 gnd 0.596792f
C4169 a_n5644_8799.n81 gnd 0.268224f
C4170 a_n5644_8799.t49 gnd 0.596792f
C4171 a_n5644_8799.t68 gnd 0.596792f
C4172 a_n5644_8799.t58 gnd 0.608087f
C4173 a_n5644_8799.n82 gnd 0.250184f
C4174 a_n5644_8799.n83 gnd 0.270608f
C4175 a_n5644_8799.t81 gnd 0.596792f
C4176 a_n5644_8799.n84 gnd 0.268224f
C4177 a_n5644_8799.n85 gnd 0.26382f
C4178 a_n5644_8799.t57 gnd 0.596792f
C4179 a_n5644_8799.n86 gnd 0.26382f
C4180 a_n5644_8799.t45 gnd 0.596792f
C4181 a_n5644_8799.n87 gnd 0.270608f
C4182 a_n5644_8799.t47 gnd 0.608077f
C4183 a_n5644_8799.n88 gnd 0.897554f
C4184 a_n5644_8799.t66 gnd 0.596792f
C4185 a_n5644_8799.n89 gnd 0.268224f
C4186 a_n5644_8799.t74 gnd 0.596792f
C4187 a_n5644_8799.t71 gnd 0.596792f
C4188 a_n5644_8799.t39 gnd 0.608087f
C4189 a_n5644_8799.n90 gnd 0.250184f
C4190 a_n5644_8799.n91 gnd 0.270608f
C4191 a_n5644_8799.t48 gnd 0.596792f
C4192 a_n5644_8799.n92 gnd 0.268224f
C4193 a_n5644_8799.n93 gnd 0.26382f
C4194 a_n5644_8799.t54 gnd 0.596792f
C4195 a_n5644_8799.n94 gnd 0.26382f
C4196 a_n5644_8799.t43 gnd 0.596792f
C4197 a_n5644_8799.n95 gnd 0.270608f
C4198 a_n5644_8799.t83 gnd 0.608077f
C4199 a_n5644_8799.n96 gnd 1.53678f
C4200 a_n5644_8799.t60 gnd 0.608077f
C4201 a_n5644_8799.t59 gnd 0.596792f
C4202 a_n5644_8799.t46 gnd 0.596792f
C4203 a_n5644_8799.n97 gnd 0.268224f
C4204 a_n5644_8799.t76 gnd 0.596792f
C4205 a_n5644_8799.t61 gnd 0.596792f
C4206 a_n5644_8799.t51 gnd 0.596792f
C4207 a_n5644_8799.n98 gnd 0.268224f
C4208 a_n5644_8799.t69 gnd 0.608087f
C4209 a_n5644_8799.n99 gnd 0.250184f
C4210 a_n5644_8799.t78 gnd 0.596792f
C4211 a_n5644_8799.n100 gnd 0.270608f
C4212 a_n5644_8799.n101 gnd 0.26382f
C4213 a_n5644_8799.n102 gnd 0.26382f
C4214 a_n5644_8799.n103 gnd 0.270608f
C4215 a_n5644_8799.t64 gnd 0.608077f
C4216 a_n5644_8799.t63 gnd 0.596792f
C4217 a_n5644_8799.t55 gnd 0.596792f
C4218 a_n5644_8799.n104 gnd 0.268224f
C4219 a_n5644_8799.t80 gnd 0.596792f
C4220 a_n5644_8799.t67 gnd 0.596792f
C4221 a_n5644_8799.t56 gnd 0.596792f
C4222 a_n5644_8799.n105 gnd 0.268224f
C4223 a_n5644_8799.t72 gnd 0.608087f
C4224 a_n5644_8799.n106 gnd 0.250184f
C4225 a_n5644_8799.t36 gnd 0.596792f
C4226 a_n5644_8799.n107 gnd 0.270608f
C4227 a_n5644_8799.n108 gnd 0.26382f
C4228 a_n5644_8799.n109 gnd 0.26382f
C4229 a_n5644_8799.n110 gnd 0.270608f
C4230 a_n5644_8799.n111 gnd 0.897554f
C4231 a_n5644_8799.t82 gnd 0.608077f
C4232 a_n5644_8799.t44 gnd 0.596792f
C4233 a_n5644_8799.t65 gnd 0.596792f
C4234 a_n5644_8799.n112 gnd 0.268224f
C4235 a_n5644_8799.t37 gnd 0.596792f
C4236 a_n5644_8799.t73 gnd 0.596792f
C4237 a_n5644_8799.t50 gnd 0.596792f
C4238 a_n5644_8799.n113 gnd 0.268224f
C4239 a_n5644_8799.t38 gnd 0.608087f
C4240 a_n5644_8799.n114 gnd 0.250184f
C4241 a_n5644_8799.t70 gnd 0.596792f
C4242 a_n5644_8799.n115 gnd 0.270608f
C4243 a_n5644_8799.n116 gnd 0.26382f
C4244 a_n5644_8799.n117 gnd 0.26382f
C4245 a_n5644_8799.n118 gnd 0.270608f
C4246 a_n5644_8799.n119 gnd 1.0844f
C4247 a_n5644_8799.n120 gnd 12.1892f
C4248 a_n5644_8799.n121 gnd 4.36765f
C4249 a_n5644_8799.n122 gnd 5.66677f
C4250 a_n5644_8799.t14 gnd 0.143928f
C4251 a_n5644_8799.t15 gnd 0.143928f
C4252 a_n5644_8799.n123 gnd 1.13331f
C4253 a_n5644_8799.t18 gnd 0.143928f
C4254 a_n5644_8799.t6 gnd 0.143928f
C4255 a_n5644_8799.n124 gnd 1.13331f
C4256 a_n5644_8799.n125 gnd 1.13518f
C4257 a_n5644_8799.t2 gnd 0.143928f
C4258 CSoutput.n0 gnd 0.03724f
C4259 CSoutput.t121 gnd 0.246336f
C4260 CSoutput.n1 gnd 0.111233f
C4261 CSoutput.n2 gnd 0.03724f
C4262 CSoutput.t125 gnd 0.246336f
C4263 CSoutput.n3 gnd 0.029516f
C4264 CSoutput.n4 gnd 0.03724f
C4265 CSoutput.t137 gnd 0.246336f
C4266 CSoutput.n5 gnd 0.025452f
C4267 CSoutput.n6 gnd 0.03724f
C4268 CSoutput.t123 gnd 0.246336f
C4269 CSoutput.t129 gnd 0.246336f
C4270 CSoutput.n7 gnd 0.110021f
C4271 CSoutput.n8 gnd 0.03724f
C4272 CSoutput.t128 gnd 0.246336f
C4273 CSoutput.n9 gnd 0.024267f
C4274 CSoutput.n10 gnd 0.03724f
C4275 CSoutput.t139 gnd 0.246336f
C4276 CSoutput.t126 gnd 0.246336f
C4277 CSoutput.n11 gnd 0.110021f
C4278 CSoutput.n12 gnd 0.03724f
C4279 CSoutput.t124 gnd 0.246336f
C4280 CSoutput.n13 gnd 0.025452f
C4281 CSoutput.n14 gnd 0.03724f
C4282 CSoutput.t138 gnd 0.246336f
C4283 CSoutput.t141 gnd 0.246336f
C4284 CSoutput.n15 gnd 0.110021f
C4285 CSoutput.n16 gnd 0.03724f
C4286 CSoutput.t122 gnd 0.246336f
C4287 CSoutput.n17 gnd 0.027184f
C4288 CSoutput.t133 gnd 0.294378f
C4289 CSoutput.t135 gnd 0.246336f
C4290 CSoutput.n18 gnd 0.140454f
C4291 CSoutput.n19 gnd 0.136289f
C4292 CSoutput.n20 gnd 0.158111f
C4293 CSoutput.n21 gnd 0.03724f
C4294 CSoutput.n22 gnd 0.031081f
C4295 CSoutput.n23 gnd 0.110021f
C4296 CSoutput.n24 gnd 0.029961f
C4297 CSoutput.n25 gnd 0.029516f
C4298 CSoutput.n26 gnd 0.03724f
C4299 CSoutput.n27 gnd 0.03724f
C4300 CSoutput.n28 gnd 0.030842f
C4301 CSoutput.n29 gnd 0.026186f
C4302 CSoutput.n30 gnd 0.11247f
C4303 CSoutput.n31 gnd 0.026546f
C4304 CSoutput.n32 gnd 0.03724f
C4305 CSoutput.n33 gnd 0.03724f
C4306 CSoutput.n34 gnd 0.03724f
C4307 CSoutput.n35 gnd 0.030514f
C4308 CSoutput.n36 gnd 0.110021f
C4309 CSoutput.n37 gnd 0.029182f
C4310 CSoutput.n38 gnd 0.030295f
C4311 CSoutput.n39 gnd 0.03724f
C4312 CSoutput.n40 gnd 0.03724f
C4313 CSoutput.n41 gnd 0.031075f
C4314 CSoutput.n42 gnd 0.028402f
C4315 CSoutput.n43 gnd 0.110021f
C4316 CSoutput.n44 gnd 0.029122f
C4317 CSoutput.n45 gnd 0.03724f
C4318 CSoutput.n46 gnd 0.03724f
C4319 CSoutput.n47 gnd 0.03724f
C4320 CSoutput.n48 gnd 0.029122f
C4321 CSoutput.n49 gnd 0.110021f
C4322 CSoutput.n50 gnd 0.028402f
C4323 CSoutput.n51 gnd 0.031075f
C4324 CSoutput.n52 gnd 0.03724f
C4325 CSoutput.n53 gnd 0.03724f
C4326 CSoutput.n54 gnd 0.030295f
C4327 CSoutput.n55 gnd 0.029182f
C4328 CSoutput.n56 gnd 0.110021f
C4329 CSoutput.n57 gnd 0.030514f
C4330 CSoutput.n58 gnd 0.03724f
C4331 CSoutput.n59 gnd 0.03724f
C4332 CSoutput.n60 gnd 0.03724f
C4333 CSoutput.n61 gnd 0.026546f
C4334 CSoutput.n62 gnd 0.11247f
C4335 CSoutput.n63 gnd 0.026186f
C4336 CSoutput.t132 gnd 0.246336f
C4337 CSoutput.n64 gnd 0.110021f
C4338 CSoutput.n65 gnd 0.030842f
C4339 CSoutput.n66 gnd 0.03724f
C4340 CSoutput.n67 gnd 0.03724f
C4341 CSoutput.n68 gnd 0.03724f
C4342 CSoutput.n69 gnd 0.029961f
C4343 CSoutput.n70 gnd 0.110021f
C4344 CSoutput.n71 gnd 0.031081f
C4345 CSoutput.n72 gnd 0.027184f
C4346 CSoutput.n73 gnd 0.03724f
C4347 CSoutput.n74 gnd 0.03724f
C4348 CSoutput.n75 gnd 0.028191f
C4349 CSoutput.n76 gnd 0.016743f
C4350 CSoutput.t134 gnd 0.276776f
C4351 CSoutput.n77 gnd 0.137491f
C4352 CSoutput.n78 gnd 0.56247f
C4353 CSoutput.t9 gnd 0.046452f
C4354 CSoutput.t110 gnd 0.046452f
C4355 CSoutput.n79 gnd 0.359646f
C4356 CSoutput.t116 gnd 0.046452f
C4357 CSoutput.t117 gnd 0.046452f
C4358 CSoutput.n80 gnd 0.359005f
C4359 CSoutput.n81 gnd 0.364389f
C4360 CSoutput.t7 gnd 0.046452f
C4361 CSoutput.t19 gnd 0.046452f
C4362 CSoutput.n82 gnd 0.359005f
C4363 CSoutput.n83 gnd 0.179556f
C4364 CSoutput.t37 gnd 0.046452f
C4365 CSoutput.t30 gnd 0.046452f
C4366 CSoutput.n84 gnd 0.359005f
C4367 CSoutput.n85 gnd 0.329264f
C4368 CSoutput.t0 gnd 0.046452f
C4369 CSoutput.t5 gnd 0.046452f
C4370 CSoutput.n86 gnd 0.359646f
C4371 CSoutput.t111 gnd 0.046452f
C4372 CSoutput.t21 gnd 0.046452f
C4373 CSoutput.n87 gnd 0.359005f
C4374 CSoutput.n88 gnd 0.364389f
C4375 CSoutput.t118 gnd 0.046452f
C4376 CSoutput.t13 gnd 0.046452f
C4377 CSoutput.n89 gnd 0.359005f
C4378 CSoutput.n90 gnd 0.179556f
C4379 CSoutput.t112 gnd 0.046452f
C4380 CSoutput.t3 gnd 0.046452f
C4381 CSoutput.n91 gnd 0.359005f
C4382 CSoutput.n92 gnd 0.267763f
C4383 CSoutput.n93 gnd 0.337647f
C4384 CSoutput.t4 gnd 0.046452f
C4385 CSoutput.t33 gnd 0.046452f
C4386 CSoutput.n94 gnd 0.359646f
C4387 CSoutput.t18 gnd 0.046452f
C4388 CSoutput.t115 gnd 0.046452f
C4389 CSoutput.n95 gnd 0.359005f
C4390 CSoutput.n96 gnd 0.364389f
C4391 CSoutput.t27 gnd 0.046452f
C4392 CSoutput.t10 gnd 0.046452f
C4393 CSoutput.n97 gnd 0.359005f
C4394 CSoutput.n98 gnd 0.179556f
C4395 CSoutput.t26 gnd 0.046452f
C4396 CSoutput.t8 gnd 0.046452f
C4397 CSoutput.n99 gnd 0.359005f
C4398 CSoutput.n100 gnd 0.267763f
C4399 CSoutput.n101 gnd 0.377403f
C4400 CSoutput.n102 gnd 6.34531f
C4401 CSoutput.n104 gnd 0.658773f
C4402 CSoutput.n105 gnd 0.494079f
C4403 CSoutput.n106 gnd 0.658773f
C4404 CSoutput.n107 gnd 0.658773f
C4405 CSoutput.n108 gnd 1.77362f
C4406 CSoutput.n109 gnd 0.658773f
C4407 CSoutput.n110 gnd 0.658773f
C4408 CSoutput.t140 gnd 0.823466f
C4409 CSoutput.n111 gnd 0.658773f
C4410 CSoutput.n112 gnd 0.658773f
C4411 CSoutput.n116 gnd 0.658773f
C4412 CSoutput.n120 gnd 0.658773f
C4413 CSoutput.n121 gnd 0.658773f
C4414 CSoutput.n123 gnd 0.658773f
C4415 CSoutput.n128 gnd 0.658773f
C4416 CSoutput.n130 gnd 0.658773f
C4417 CSoutput.n131 gnd 0.658773f
C4418 CSoutput.n133 gnd 0.658773f
C4419 CSoutput.n134 gnd 0.658773f
C4420 CSoutput.n136 gnd 0.658773f
C4421 CSoutput.t130 gnd 11.008f
C4422 CSoutput.n138 gnd 0.658773f
C4423 CSoutput.n139 gnd 0.494079f
C4424 CSoutput.n140 gnd 0.658773f
C4425 CSoutput.n141 gnd 0.658773f
C4426 CSoutput.n142 gnd 1.77362f
C4427 CSoutput.n143 gnd 0.658773f
C4428 CSoutput.n144 gnd 0.658773f
C4429 CSoutput.t127 gnd 0.823466f
C4430 CSoutput.n145 gnd 0.658773f
C4431 CSoutput.n146 gnd 0.658773f
C4432 CSoutput.n150 gnd 0.658773f
C4433 CSoutput.n154 gnd 0.658773f
C4434 CSoutput.n155 gnd 0.658773f
C4435 CSoutput.n157 gnd 0.658773f
C4436 CSoutput.n162 gnd 0.658773f
C4437 CSoutput.n164 gnd 0.658773f
C4438 CSoutput.n165 gnd 0.658773f
C4439 CSoutput.n167 gnd 0.658773f
C4440 CSoutput.n168 gnd 0.658773f
C4441 CSoutput.n170 gnd 0.658773f
C4442 CSoutput.n171 gnd 0.494079f
C4443 CSoutput.n173 gnd 0.658773f
C4444 CSoutput.n174 gnd 0.494079f
C4445 CSoutput.n175 gnd 0.658773f
C4446 CSoutput.n176 gnd 0.658773f
C4447 CSoutput.n177 gnd 1.77362f
C4448 CSoutput.n178 gnd 0.658773f
C4449 CSoutput.n179 gnd 0.658773f
C4450 CSoutput.t120 gnd 0.823466f
C4451 CSoutput.n180 gnd 0.658773f
C4452 CSoutput.n181 gnd 1.77362f
C4453 CSoutput.n183 gnd 0.658773f
C4454 CSoutput.n184 gnd 0.658773f
C4455 CSoutput.n186 gnd 0.658773f
C4456 CSoutput.n187 gnd 0.658773f
C4457 CSoutput.t131 gnd 10.8286f
C4458 CSoutput.t136 gnd 11.008f
C4459 CSoutput.n193 gnd 2.06667f
C4460 CSoutput.n194 gnd 8.418849f
C4461 CSoutput.n195 gnd 8.77112f
C4462 CSoutput.n200 gnd 2.23876f
C4463 CSoutput.n206 gnd 0.658773f
C4464 CSoutput.n208 gnd 0.658773f
C4465 CSoutput.n210 gnd 0.658773f
C4466 CSoutput.n212 gnd 0.658773f
C4467 CSoutput.n214 gnd 0.658773f
C4468 CSoutput.n220 gnd 0.658773f
C4469 CSoutput.n227 gnd 1.20859f
C4470 CSoutput.n228 gnd 1.20859f
C4471 CSoutput.n229 gnd 0.658773f
C4472 CSoutput.n230 gnd 0.658773f
C4473 CSoutput.n232 gnd 0.494079f
C4474 CSoutput.n233 gnd 0.423135f
C4475 CSoutput.n235 gnd 0.494079f
C4476 CSoutput.n236 gnd 0.423135f
C4477 CSoutput.n237 gnd 0.494079f
C4478 CSoutput.n239 gnd 0.658773f
C4479 CSoutput.n241 gnd 1.77362f
C4480 CSoutput.n242 gnd 2.06667f
C4481 CSoutput.n243 gnd 7.74317f
C4482 CSoutput.n245 gnd 0.494079f
C4483 CSoutput.n246 gnd 1.2713f
C4484 CSoutput.n247 gnd 0.494079f
C4485 CSoutput.n249 gnd 0.658773f
C4486 CSoutput.n251 gnd 1.77362f
C4487 CSoutput.n252 gnd 3.86323f
C4488 CSoutput.t22 gnd 0.046452f
C4489 CSoutput.t14 gnd 0.046452f
C4490 CSoutput.n253 gnd 0.359646f
C4491 CSoutput.t29 gnd 0.046452f
C4492 CSoutput.t31 gnd 0.046452f
C4493 CSoutput.n254 gnd 0.359005f
C4494 CSoutput.n255 gnd 0.364389f
C4495 CSoutput.t12 gnd 0.046452f
C4496 CSoutput.t1 gnd 0.046452f
C4497 CSoutput.n256 gnd 0.359005f
C4498 CSoutput.n257 gnd 0.179556f
C4499 CSoutput.t25 gnd 0.046452f
C4500 CSoutput.t16 gnd 0.046452f
C4501 CSoutput.n258 gnd 0.359005f
C4502 CSoutput.n259 gnd 0.329264f
C4503 CSoutput.t15 gnd 0.046452f
C4504 CSoutput.t23 gnd 0.046452f
C4505 CSoutput.n260 gnd 0.359646f
C4506 CSoutput.t20 gnd 0.046452f
C4507 CSoutput.t24 gnd 0.046452f
C4508 CSoutput.n261 gnd 0.359005f
C4509 CSoutput.n262 gnd 0.364389f
C4510 CSoutput.t11 gnd 0.046452f
C4511 CSoutput.t36 gnd 0.046452f
C4512 CSoutput.n263 gnd 0.359005f
C4513 CSoutput.n264 gnd 0.179556f
C4514 CSoutput.t113 gnd 0.046452f
C4515 CSoutput.t17 gnd 0.046452f
C4516 CSoutput.n265 gnd 0.359005f
C4517 CSoutput.n266 gnd 0.267763f
C4518 CSoutput.n267 gnd 0.337647f
C4519 CSoutput.t114 gnd 0.046452f
C4520 CSoutput.t6 gnd 0.046452f
C4521 CSoutput.n268 gnd 0.359646f
C4522 CSoutput.t119 gnd 0.046452f
C4523 CSoutput.t34 gnd 0.046452f
C4524 CSoutput.n269 gnd 0.359005f
C4525 CSoutput.n270 gnd 0.364389f
C4526 CSoutput.t32 gnd 0.046452f
C4527 CSoutput.t28 gnd 0.046452f
C4528 CSoutput.n271 gnd 0.359005f
C4529 CSoutput.n272 gnd 0.179556f
C4530 CSoutput.t2 gnd 0.046452f
C4531 CSoutput.t35 gnd 0.046452f
C4532 CSoutput.n273 gnd 0.359004f
C4533 CSoutput.n274 gnd 0.267764f
C4534 CSoutput.n275 gnd 0.377403f
C4535 CSoutput.n276 gnd 9.31949f
C4536 CSoutput.t68 gnd 0.040645f
C4537 CSoutput.t108 gnd 0.040645f
C4538 CSoutput.n277 gnd 0.360359f
C4539 CSoutput.t62 gnd 0.040645f
C4540 CSoutput.t67 gnd 0.040645f
C4541 CSoutput.n278 gnd 0.359157f
C4542 CSoutput.n279 gnd 0.334667f
C4543 CSoutput.t57 gnd 0.040645f
C4544 CSoutput.t71 gnd 0.040645f
C4545 CSoutput.n280 gnd 0.359157f
C4546 CSoutput.n281 gnd 0.164975f
C4547 CSoutput.t80 gnd 0.040645f
C4548 CSoutput.t63 gnd 0.040645f
C4549 CSoutput.n282 gnd 0.359157f
C4550 CSoutput.n283 gnd 0.164975f
C4551 CSoutput.t69 gnd 0.040645f
C4552 CSoutput.t97 gnd 0.040645f
C4553 CSoutput.n284 gnd 0.359157f
C4554 CSoutput.n285 gnd 0.164975f
C4555 CSoutput.t77 gnd 0.040645f
C4556 CSoutput.t84 gnd 0.040645f
C4557 CSoutput.n286 gnd 0.359157f
C4558 CSoutput.n287 gnd 0.304288f
C4559 CSoutput.t105 gnd 0.040645f
C4560 CSoutput.t38 gnd 0.040645f
C4561 CSoutput.n288 gnd 0.360359f
C4562 CSoutput.t47 gnd 0.040645f
C4563 CSoutput.t98 gnd 0.040645f
C4564 CSoutput.n289 gnd 0.359157f
C4565 CSoutput.n290 gnd 0.334667f
C4566 CSoutput.t39 gnd 0.040645f
C4567 CSoutput.t92 gnd 0.040645f
C4568 CSoutput.n291 gnd 0.359157f
C4569 CSoutput.n292 gnd 0.164975f
C4570 CSoutput.t99 gnd 0.040645f
C4571 CSoutput.t40 gnd 0.040645f
C4572 CSoutput.n293 gnd 0.359157f
C4573 CSoutput.n294 gnd 0.164975f
C4574 CSoutput.t86 gnd 0.040645f
C4575 CSoutput.t74 gnd 0.040645f
C4576 CSoutput.n295 gnd 0.359157f
C4577 CSoutput.n296 gnd 0.164975f
C4578 CSoutput.t41 gnd 0.040645f
C4579 CSoutput.t88 gnd 0.040645f
C4580 CSoutput.n297 gnd 0.359157f
C4581 CSoutput.n298 gnd 0.250468f
C4582 CSoutput.n299 gnd 0.315918f
C4583 CSoutput.t48 gnd 0.040645f
C4584 CSoutput.t100 gnd 0.040645f
C4585 CSoutput.n300 gnd 0.360359f
C4586 CSoutput.t61 gnd 0.040645f
C4587 CSoutput.t64 gnd 0.040645f
C4588 CSoutput.n301 gnd 0.359157f
C4589 CSoutput.n302 gnd 0.334667f
C4590 CSoutput.t42 gnd 0.040645f
C4591 CSoutput.t90 gnd 0.040645f
C4592 CSoutput.n303 gnd 0.359157f
C4593 CSoutput.n304 gnd 0.164975f
C4594 CSoutput.t70 gnd 0.040645f
C4595 CSoutput.t49 gnd 0.040645f
C4596 CSoutput.n305 gnd 0.359157f
C4597 CSoutput.n306 gnd 0.164975f
C4598 CSoutput.t54 gnd 0.040645f
C4599 CSoutput.t109 gnd 0.040645f
C4600 CSoutput.n307 gnd 0.359157f
C4601 CSoutput.n308 gnd 0.164975f
C4602 CSoutput.t55 gnd 0.040645f
C4603 CSoutput.t59 gnd 0.040645f
C4604 CSoutput.n309 gnd 0.359157f
C4605 CSoutput.n310 gnd 0.250468f
C4606 CSoutput.n311 gnd 0.339246f
C4607 CSoutput.n312 gnd 9.773809f
C4608 CSoutput.t58 gnd 0.040645f
C4609 CSoutput.t87 gnd 0.040645f
C4610 CSoutput.n313 gnd 0.360359f
C4611 CSoutput.t85 gnd 0.040645f
C4612 CSoutput.t73 gnd 0.040645f
C4613 CSoutput.n314 gnd 0.359157f
C4614 CSoutput.n315 gnd 0.334667f
C4615 CSoutput.t91 gnd 0.040645f
C4616 CSoutput.t65 gnd 0.040645f
C4617 CSoutput.n316 gnd 0.359157f
C4618 CSoutput.n317 gnd 0.164975f
C4619 CSoutput.t78 gnd 0.040645f
C4620 CSoutput.t101 gnd 0.040645f
C4621 CSoutput.n318 gnd 0.359157f
C4622 CSoutput.n319 gnd 0.164975f
C4623 CSoutput.t53 gnd 0.040645f
C4624 CSoutput.t89 gnd 0.040645f
C4625 CSoutput.n320 gnd 0.359157f
C4626 CSoutput.n321 gnd 0.164975f
C4627 CSoutput.t46 gnd 0.040645f
C4628 CSoutput.t93 gnd 0.040645f
C4629 CSoutput.n322 gnd 0.359157f
C4630 CSoutput.n323 gnd 0.304288f
C4631 CSoutput.t50 gnd 0.040645f
C4632 CSoutput.t45 gnd 0.040645f
C4633 CSoutput.n324 gnd 0.360359f
C4634 CSoutput.t43 gnd 0.040645f
C4635 CSoutput.t106 gnd 0.040645f
C4636 CSoutput.n325 gnd 0.359157f
C4637 CSoutput.n326 gnd 0.334667f
C4638 CSoutput.t107 gnd 0.040645f
C4639 CSoutput.t51 gnd 0.040645f
C4640 CSoutput.n327 gnd 0.359157f
C4641 CSoutput.n328 gnd 0.164975f
C4642 CSoutput.t52 gnd 0.040645f
C4643 CSoutput.t81 gnd 0.040645f
C4644 CSoutput.n329 gnd 0.359157f
C4645 CSoutput.n330 gnd 0.164975f
C4646 CSoutput.t82 gnd 0.040645f
C4647 CSoutput.t102 gnd 0.040645f
C4648 CSoutput.n331 gnd 0.359157f
C4649 CSoutput.n332 gnd 0.164975f
C4650 CSoutput.t103 gnd 0.040645f
C4651 CSoutput.t96 gnd 0.040645f
C4652 CSoutput.n333 gnd 0.359157f
C4653 CSoutput.n334 gnd 0.250468f
C4654 CSoutput.n335 gnd 0.315918f
C4655 CSoutput.t76 gnd 0.040645f
C4656 CSoutput.t94 gnd 0.040645f
C4657 CSoutput.n336 gnd 0.360359f
C4658 CSoutput.t56 gnd 0.040645f
C4659 CSoutput.t66 gnd 0.040645f
C4660 CSoutput.n337 gnd 0.359157f
C4661 CSoutput.n338 gnd 0.334667f
C4662 CSoutput.t72 gnd 0.040645f
C4663 CSoutput.t83 gnd 0.040645f
C4664 CSoutput.n339 gnd 0.359157f
C4665 CSoutput.n340 gnd 0.164975f
C4666 CSoutput.t95 gnd 0.040645f
C4667 CSoutput.t75 gnd 0.040645f
C4668 CSoutput.n341 gnd 0.359157f
C4669 CSoutput.n342 gnd 0.164975f
C4670 CSoutput.t79 gnd 0.040645f
C4671 CSoutput.t104 gnd 0.040645f
C4672 CSoutput.n343 gnd 0.359157f
C4673 CSoutput.n344 gnd 0.164975f
C4674 CSoutput.t44 gnd 0.040645f
C4675 CSoutput.t60 gnd 0.040645f
C4676 CSoutput.n345 gnd 0.359157f
C4677 CSoutput.n346 gnd 0.250468f
C4678 CSoutput.n347 gnd 0.339246f
C4679 CSoutput.n348 gnd 5.35614f
C4680 CSoutput.n349 gnd 11.3754f
C4681 commonsourceibias.n0 gnd 0.012292f
C4682 commonsourceibias.t89 gnd 0.186134f
C4683 commonsourceibias.t49 gnd 0.172107f
C4684 commonsourceibias.n1 gnd 0.068671f
C4685 commonsourceibias.n2 gnd 0.009212f
C4686 commonsourceibias.t95 gnd 0.172107f
C4687 commonsourceibias.n3 gnd 0.007452f
C4688 commonsourceibias.n4 gnd 0.009212f
C4689 commonsourceibias.t90 gnd 0.172107f
C4690 commonsourceibias.n5 gnd 0.008893f
C4691 commonsourceibias.n6 gnd 0.009212f
C4692 commonsourceibias.t100 gnd 0.172107f
C4693 commonsourceibias.n7 gnd 0.068671f
C4694 commonsourceibias.t86 gnd 0.172107f
C4695 commonsourceibias.n8 gnd 0.00744f
C4696 commonsourceibias.n9 gnd 0.012292f
C4697 commonsourceibias.t22 gnd 0.186134f
C4698 commonsourceibias.t2 gnd 0.172107f
C4699 commonsourceibias.n10 gnd 0.068671f
C4700 commonsourceibias.n11 gnd 0.009212f
C4701 commonsourceibias.t32 gnd 0.172107f
C4702 commonsourceibias.n12 gnd 0.007452f
C4703 commonsourceibias.n13 gnd 0.009212f
C4704 commonsourceibias.t20 gnd 0.172107f
C4705 commonsourceibias.n14 gnd 0.008893f
C4706 commonsourceibias.n15 gnd 0.009212f
C4707 commonsourceibias.t40 gnd 0.172107f
C4708 commonsourceibias.n16 gnd 0.068671f
C4709 commonsourceibias.t18 gnd 0.172107f
C4710 commonsourceibias.n17 gnd 0.00744f
C4711 commonsourceibias.n18 gnd 0.009212f
C4712 commonsourceibias.t6 gnd 0.172107f
C4713 commonsourceibias.t34 gnd 0.172107f
C4714 commonsourceibias.n19 gnd 0.068671f
C4715 commonsourceibias.n20 gnd 0.009212f
C4716 commonsourceibias.t24 gnd 0.172107f
C4717 commonsourceibias.n21 gnd 0.068671f
C4718 commonsourceibias.n22 gnd 0.009212f
C4719 commonsourceibias.t28 gnd 0.172107f
C4720 commonsourceibias.n23 gnd 0.068671f
C4721 commonsourceibias.n24 gnd 0.046375f
C4722 commonsourceibias.t44 gnd 0.172107f
C4723 commonsourceibias.t8 gnd 0.194203f
C4724 commonsourceibias.n25 gnd 0.079692f
C4725 commonsourceibias.n26 gnd 0.082502f
C4726 commonsourceibias.n27 gnd 0.011354f
C4727 commonsourceibias.n28 gnd 0.012561f
C4728 commonsourceibias.n29 gnd 0.009212f
C4729 commonsourceibias.n30 gnd 0.009212f
C4730 commonsourceibias.n31 gnd 0.012479f
C4731 commonsourceibias.n32 gnd 0.007452f
C4732 commonsourceibias.n33 gnd 0.012633f
C4733 commonsourceibias.n34 gnd 0.009212f
C4734 commonsourceibias.n35 gnd 0.009212f
C4735 commonsourceibias.n36 gnd 0.01271f
C4736 commonsourceibias.n37 gnd 0.01096f
C4737 commonsourceibias.n38 gnd 0.008893f
C4738 commonsourceibias.n39 gnd 0.009212f
C4739 commonsourceibias.n40 gnd 0.009212f
C4740 commonsourceibias.n41 gnd 0.011268f
C4741 commonsourceibias.n42 gnd 0.012647f
C4742 commonsourceibias.n43 gnd 0.068671f
C4743 commonsourceibias.n44 gnd 0.012562f
C4744 commonsourceibias.n45 gnd 0.009212f
C4745 commonsourceibias.n46 gnd 0.009212f
C4746 commonsourceibias.n47 gnd 0.009212f
C4747 commonsourceibias.n48 gnd 0.012562f
C4748 commonsourceibias.n49 gnd 0.068671f
C4749 commonsourceibias.n50 gnd 0.012647f
C4750 commonsourceibias.n51 gnd 0.011268f
C4751 commonsourceibias.n52 gnd 0.009212f
C4752 commonsourceibias.n53 gnd 0.009212f
C4753 commonsourceibias.n54 gnd 0.009212f
C4754 commonsourceibias.n55 gnd 0.01096f
C4755 commonsourceibias.n56 gnd 0.01271f
C4756 commonsourceibias.n57 gnd 0.068671f
C4757 commonsourceibias.n58 gnd 0.012633f
C4758 commonsourceibias.n59 gnd 0.009212f
C4759 commonsourceibias.n60 gnd 0.009212f
C4760 commonsourceibias.n61 gnd 0.009212f
C4761 commonsourceibias.n62 gnd 0.012479f
C4762 commonsourceibias.n63 gnd 0.068671f
C4763 commonsourceibias.n64 gnd 0.012561f
C4764 commonsourceibias.n65 gnd 0.011354f
C4765 commonsourceibias.n66 gnd 0.009212f
C4766 commonsourceibias.n67 gnd 0.009212f
C4767 commonsourceibias.n68 gnd 0.009345f
C4768 commonsourceibias.n69 gnd 0.009661f
C4769 commonsourceibias.n70 gnd 0.082165f
C4770 commonsourceibias.n71 gnd 0.09115f
C4771 commonsourceibias.t23 gnd 0.019878f
C4772 commonsourceibias.t3 gnd 0.019878f
C4773 commonsourceibias.n72 gnd 0.175652f
C4774 commonsourceibias.n73 gnd 0.151777f
C4775 commonsourceibias.t33 gnd 0.019878f
C4776 commonsourceibias.t21 gnd 0.019878f
C4777 commonsourceibias.n74 gnd 0.175652f
C4778 commonsourceibias.n75 gnd 0.080684f
C4779 commonsourceibias.t41 gnd 0.019878f
C4780 commonsourceibias.t19 gnd 0.019878f
C4781 commonsourceibias.n76 gnd 0.175652f
C4782 commonsourceibias.n77 gnd 0.067408f
C4783 commonsourceibias.t45 gnd 0.019878f
C4784 commonsourceibias.t9 gnd 0.019878f
C4785 commonsourceibias.n78 gnd 0.17624f
C4786 commonsourceibias.t25 gnd 0.019878f
C4787 commonsourceibias.t29 gnd 0.019878f
C4788 commonsourceibias.n79 gnd 0.175652f
C4789 commonsourceibias.n80 gnd 0.163675f
C4790 commonsourceibias.t7 gnd 0.019878f
C4791 commonsourceibias.t35 gnd 0.019878f
C4792 commonsourceibias.n81 gnd 0.175652f
C4793 commonsourceibias.n82 gnd 0.067408f
C4794 commonsourceibias.n83 gnd 0.081623f
C4795 commonsourceibias.n84 gnd 0.009212f
C4796 commonsourceibias.t77 gnd 0.172107f
C4797 commonsourceibias.t94 gnd 0.172107f
C4798 commonsourceibias.n85 gnd 0.068671f
C4799 commonsourceibias.n86 gnd 0.009212f
C4800 commonsourceibias.t88 gnd 0.172107f
C4801 commonsourceibias.n87 gnd 0.068671f
C4802 commonsourceibias.n88 gnd 0.009212f
C4803 commonsourceibias.t60 gnd 0.172107f
C4804 commonsourceibias.n89 gnd 0.068671f
C4805 commonsourceibias.n90 gnd 0.046375f
C4806 commonsourceibias.t80 gnd 0.172107f
C4807 commonsourceibias.t73 gnd 0.194203f
C4808 commonsourceibias.n91 gnd 0.079692f
C4809 commonsourceibias.n92 gnd 0.082502f
C4810 commonsourceibias.n93 gnd 0.011354f
C4811 commonsourceibias.n94 gnd 0.012561f
C4812 commonsourceibias.n95 gnd 0.009212f
C4813 commonsourceibias.n96 gnd 0.009212f
C4814 commonsourceibias.n97 gnd 0.012479f
C4815 commonsourceibias.n98 gnd 0.007452f
C4816 commonsourceibias.n99 gnd 0.012633f
C4817 commonsourceibias.n100 gnd 0.009212f
C4818 commonsourceibias.n101 gnd 0.009212f
C4819 commonsourceibias.n102 gnd 0.01271f
C4820 commonsourceibias.n103 gnd 0.01096f
C4821 commonsourceibias.n104 gnd 0.008893f
C4822 commonsourceibias.n105 gnd 0.009212f
C4823 commonsourceibias.n106 gnd 0.009212f
C4824 commonsourceibias.n107 gnd 0.011268f
C4825 commonsourceibias.n108 gnd 0.012647f
C4826 commonsourceibias.n109 gnd 0.068671f
C4827 commonsourceibias.n110 gnd 0.012562f
C4828 commonsourceibias.n111 gnd 0.009168f
C4829 commonsourceibias.n112 gnd 0.066591f
C4830 commonsourceibias.n113 gnd 0.009168f
C4831 commonsourceibias.n114 gnd 0.012562f
C4832 commonsourceibias.n115 gnd 0.068671f
C4833 commonsourceibias.n116 gnd 0.012647f
C4834 commonsourceibias.n117 gnd 0.011268f
C4835 commonsourceibias.n118 gnd 0.009212f
C4836 commonsourceibias.n119 gnd 0.009212f
C4837 commonsourceibias.n120 gnd 0.009212f
C4838 commonsourceibias.n121 gnd 0.01096f
C4839 commonsourceibias.n122 gnd 0.01271f
C4840 commonsourceibias.n123 gnd 0.068671f
C4841 commonsourceibias.n124 gnd 0.012633f
C4842 commonsourceibias.n125 gnd 0.009212f
C4843 commonsourceibias.n126 gnd 0.009212f
C4844 commonsourceibias.n127 gnd 0.009212f
C4845 commonsourceibias.n128 gnd 0.012479f
C4846 commonsourceibias.n129 gnd 0.068671f
C4847 commonsourceibias.n130 gnd 0.012561f
C4848 commonsourceibias.n131 gnd 0.011354f
C4849 commonsourceibias.n132 gnd 0.009212f
C4850 commonsourceibias.n133 gnd 0.009212f
C4851 commonsourceibias.n134 gnd 0.009345f
C4852 commonsourceibias.n135 gnd 0.009661f
C4853 commonsourceibias.n136 gnd 0.082165f
C4854 commonsourceibias.n137 gnd 0.053193f
C4855 commonsourceibias.n138 gnd 0.012292f
C4856 commonsourceibias.t52 gnd 0.186134f
C4857 commonsourceibias.t119 gnd 0.172107f
C4858 commonsourceibias.n139 gnd 0.068671f
C4859 commonsourceibias.n140 gnd 0.009212f
C4860 commonsourceibias.t110 gnd 0.172107f
C4861 commonsourceibias.n141 gnd 0.007452f
C4862 commonsourceibias.n142 gnd 0.009212f
C4863 commonsourceibias.t59 gnd 0.172107f
C4864 commonsourceibias.n143 gnd 0.008893f
C4865 commonsourceibias.n144 gnd 0.009212f
C4866 commonsourceibias.t118 gnd 0.172107f
C4867 commonsourceibias.n145 gnd 0.068671f
C4868 commonsourceibias.t65 gnd 0.172107f
C4869 commonsourceibias.n146 gnd 0.00744f
C4870 commonsourceibias.n147 gnd 0.009212f
C4871 commonsourceibias.t58 gnd 0.172107f
C4872 commonsourceibias.t117 gnd 0.172107f
C4873 commonsourceibias.n148 gnd 0.068671f
C4874 commonsourceibias.n149 gnd 0.009212f
C4875 commonsourceibias.t71 gnd 0.172107f
C4876 commonsourceibias.n150 gnd 0.068671f
C4877 commonsourceibias.n151 gnd 0.009212f
C4878 commonsourceibias.t83 gnd 0.172107f
C4879 commonsourceibias.n152 gnd 0.068671f
C4880 commonsourceibias.n153 gnd 0.046375f
C4881 commonsourceibias.t116 gnd 0.172107f
C4882 commonsourceibias.t69 gnd 0.194203f
C4883 commonsourceibias.n154 gnd 0.079692f
C4884 commonsourceibias.n155 gnd 0.082502f
C4885 commonsourceibias.n156 gnd 0.011354f
C4886 commonsourceibias.n157 gnd 0.012561f
C4887 commonsourceibias.n158 gnd 0.009212f
C4888 commonsourceibias.n159 gnd 0.009212f
C4889 commonsourceibias.n160 gnd 0.012479f
C4890 commonsourceibias.n161 gnd 0.007452f
C4891 commonsourceibias.n162 gnd 0.012633f
C4892 commonsourceibias.n163 gnd 0.009212f
C4893 commonsourceibias.n164 gnd 0.009212f
C4894 commonsourceibias.n165 gnd 0.01271f
C4895 commonsourceibias.n166 gnd 0.01096f
C4896 commonsourceibias.n167 gnd 0.008893f
C4897 commonsourceibias.n168 gnd 0.009212f
C4898 commonsourceibias.n169 gnd 0.009212f
C4899 commonsourceibias.n170 gnd 0.011268f
C4900 commonsourceibias.n171 gnd 0.012647f
C4901 commonsourceibias.n172 gnd 0.068671f
C4902 commonsourceibias.n173 gnd 0.012562f
C4903 commonsourceibias.n174 gnd 0.009212f
C4904 commonsourceibias.n175 gnd 0.009212f
C4905 commonsourceibias.n176 gnd 0.009212f
C4906 commonsourceibias.n177 gnd 0.012562f
C4907 commonsourceibias.n178 gnd 0.068671f
C4908 commonsourceibias.n179 gnd 0.012647f
C4909 commonsourceibias.n180 gnd 0.011268f
C4910 commonsourceibias.n181 gnd 0.009212f
C4911 commonsourceibias.n182 gnd 0.009212f
C4912 commonsourceibias.n183 gnd 0.009212f
C4913 commonsourceibias.n184 gnd 0.01096f
C4914 commonsourceibias.n185 gnd 0.01271f
C4915 commonsourceibias.n186 gnd 0.068671f
C4916 commonsourceibias.n187 gnd 0.012633f
C4917 commonsourceibias.n188 gnd 0.009212f
C4918 commonsourceibias.n189 gnd 0.009212f
C4919 commonsourceibias.n190 gnd 0.009212f
C4920 commonsourceibias.n191 gnd 0.012479f
C4921 commonsourceibias.n192 gnd 0.068671f
C4922 commonsourceibias.n193 gnd 0.012561f
C4923 commonsourceibias.n194 gnd 0.011354f
C4924 commonsourceibias.n195 gnd 0.009212f
C4925 commonsourceibias.n196 gnd 0.009212f
C4926 commonsourceibias.n197 gnd 0.009345f
C4927 commonsourceibias.n198 gnd 0.009661f
C4928 commonsourceibias.n199 gnd 0.082165f
C4929 commonsourceibias.n200 gnd 0.027962f
C4930 commonsourceibias.n201 gnd 0.146988f
C4931 commonsourceibias.n202 gnd 0.012292f
C4932 commonsourceibias.t57 gnd 0.172107f
C4933 commonsourceibias.n203 gnd 0.068671f
C4934 commonsourceibias.n204 gnd 0.009212f
C4935 commonsourceibias.t96 gnd 0.172107f
C4936 commonsourceibias.n205 gnd 0.007452f
C4937 commonsourceibias.n206 gnd 0.009212f
C4938 commonsourceibias.t93 gnd 0.172107f
C4939 commonsourceibias.n207 gnd 0.008893f
C4940 commonsourceibias.n208 gnd 0.009212f
C4941 commonsourceibias.t115 gnd 0.172107f
C4942 commonsourceibias.n209 gnd 0.068671f
C4943 commonsourceibias.t67 gnd 0.172107f
C4944 commonsourceibias.n210 gnd 0.00744f
C4945 commonsourceibias.n211 gnd 0.009212f
C4946 commonsourceibias.t87 gnd 0.172107f
C4947 commonsourceibias.t108 gnd 0.172107f
C4948 commonsourceibias.n212 gnd 0.068671f
C4949 commonsourceibias.n213 gnd 0.009212f
C4950 commonsourceibias.t103 gnd 0.172107f
C4951 commonsourceibias.n214 gnd 0.068671f
C4952 commonsourceibias.n215 gnd 0.009212f
C4953 commonsourceibias.t48 gnd 0.172107f
C4954 commonsourceibias.n216 gnd 0.068671f
C4955 commonsourceibias.n217 gnd 0.046375f
C4956 commonsourceibias.t102 gnd 0.172107f
C4957 commonsourceibias.t98 gnd 0.194203f
C4958 commonsourceibias.n218 gnd 0.079692f
C4959 commonsourceibias.n219 gnd 0.082502f
C4960 commonsourceibias.n220 gnd 0.011354f
C4961 commonsourceibias.n221 gnd 0.012561f
C4962 commonsourceibias.n222 gnd 0.009212f
C4963 commonsourceibias.n223 gnd 0.009212f
C4964 commonsourceibias.n224 gnd 0.012479f
C4965 commonsourceibias.n225 gnd 0.007452f
C4966 commonsourceibias.n226 gnd 0.012633f
C4967 commonsourceibias.n227 gnd 0.009212f
C4968 commonsourceibias.n228 gnd 0.009212f
C4969 commonsourceibias.n229 gnd 0.01271f
C4970 commonsourceibias.n230 gnd 0.01096f
C4971 commonsourceibias.n231 gnd 0.008893f
C4972 commonsourceibias.n232 gnd 0.009212f
C4973 commonsourceibias.n233 gnd 0.009212f
C4974 commonsourceibias.n234 gnd 0.011268f
C4975 commonsourceibias.n235 gnd 0.012647f
C4976 commonsourceibias.n236 gnd 0.068671f
C4977 commonsourceibias.n237 gnd 0.012562f
C4978 commonsourceibias.n238 gnd 0.009212f
C4979 commonsourceibias.n239 gnd 0.009212f
C4980 commonsourceibias.n240 gnd 0.009212f
C4981 commonsourceibias.n241 gnd 0.012562f
C4982 commonsourceibias.n242 gnd 0.068671f
C4983 commonsourceibias.n243 gnd 0.012647f
C4984 commonsourceibias.n244 gnd 0.011268f
C4985 commonsourceibias.n245 gnd 0.009212f
C4986 commonsourceibias.n246 gnd 0.009212f
C4987 commonsourceibias.n247 gnd 0.009212f
C4988 commonsourceibias.n248 gnd 0.01096f
C4989 commonsourceibias.n249 gnd 0.01271f
C4990 commonsourceibias.n250 gnd 0.068671f
C4991 commonsourceibias.n251 gnd 0.012633f
C4992 commonsourceibias.n252 gnd 0.009212f
C4993 commonsourceibias.n253 gnd 0.009212f
C4994 commonsourceibias.n254 gnd 0.009212f
C4995 commonsourceibias.n255 gnd 0.012479f
C4996 commonsourceibias.n256 gnd 0.068671f
C4997 commonsourceibias.n257 gnd 0.012561f
C4998 commonsourceibias.n258 gnd 0.011354f
C4999 commonsourceibias.n259 gnd 0.009212f
C5000 commonsourceibias.n260 gnd 0.009212f
C5001 commonsourceibias.n261 gnd 0.009345f
C5002 commonsourceibias.n262 gnd 0.009661f
C5003 commonsourceibias.t109 gnd 0.186134f
C5004 commonsourceibias.n263 gnd 0.082165f
C5005 commonsourceibias.n264 gnd 0.027962f
C5006 commonsourceibias.n265 gnd 0.437625f
C5007 commonsourceibias.n266 gnd 0.012292f
C5008 commonsourceibias.t70 gnd 0.186134f
C5009 commonsourceibias.t99 gnd 0.172107f
C5010 commonsourceibias.n267 gnd 0.068671f
C5011 commonsourceibias.n268 gnd 0.009212f
C5012 commonsourceibias.t84 gnd 0.172107f
C5013 commonsourceibias.n269 gnd 0.007452f
C5014 commonsourceibias.n270 gnd 0.009212f
C5015 commonsourceibias.t72 gnd 0.172107f
C5016 commonsourceibias.n271 gnd 0.008893f
C5017 commonsourceibias.n272 gnd 0.009212f
C5018 commonsourceibias.t66 gnd 0.172107f
C5019 commonsourceibias.n273 gnd 0.00744f
C5020 commonsourceibias.n274 gnd 0.009212f
C5021 commonsourceibias.t56 gnd 0.172107f
C5022 commonsourceibias.t79 gnd 0.172107f
C5023 commonsourceibias.n275 gnd 0.068671f
C5024 commonsourceibias.n276 gnd 0.009212f
C5025 commonsourceibias.t68 gnd 0.172107f
C5026 commonsourceibias.n277 gnd 0.068671f
C5027 commonsourceibias.n278 gnd 0.009212f
C5028 commonsourceibias.t104 gnd 0.172107f
C5029 commonsourceibias.n279 gnd 0.068671f
C5030 commonsourceibias.n280 gnd 0.046375f
C5031 commonsourceibias.t64 gnd 0.172107f
C5032 commonsourceibias.t111 gnd 0.194203f
C5033 commonsourceibias.n281 gnd 0.079692f
C5034 commonsourceibias.n282 gnd 0.082502f
C5035 commonsourceibias.n283 gnd 0.011354f
C5036 commonsourceibias.n284 gnd 0.012561f
C5037 commonsourceibias.n285 gnd 0.009212f
C5038 commonsourceibias.n286 gnd 0.009212f
C5039 commonsourceibias.n287 gnd 0.012479f
C5040 commonsourceibias.n288 gnd 0.007452f
C5041 commonsourceibias.n289 gnd 0.012633f
C5042 commonsourceibias.n290 gnd 0.009212f
C5043 commonsourceibias.n291 gnd 0.009212f
C5044 commonsourceibias.n292 gnd 0.01271f
C5045 commonsourceibias.n293 gnd 0.01096f
C5046 commonsourceibias.n294 gnd 0.008893f
C5047 commonsourceibias.n295 gnd 0.009212f
C5048 commonsourceibias.n296 gnd 0.009212f
C5049 commonsourceibias.n297 gnd 0.011268f
C5050 commonsourceibias.n298 gnd 0.012647f
C5051 commonsourceibias.n299 gnd 0.068671f
C5052 commonsourceibias.n300 gnd 0.012562f
C5053 commonsourceibias.n301 gnd 0.009168f
C5054 commonsourceibias.t5 gnd 0.019878f
C5055 commonsourceibias.t27 gnd 0.019878f
C5056 commonsourceibias.n302 gnd 0.17624f
C5057 commonsourceibias.t39 gnd 0.019878f
C5058 commonsourceibias.t15 gnd 0.019878f
C5059 commonsourceibias.n303 gnd 0.175652f
C5060 commonsourceibias.n304 gnd 0.163675f
C5061 commonsourceibias.t47 gnd 0.019878f
C5062 commonsourceibias.t31 gnd 0.019878f
C5063 commonsourceibias.n305 gnd 0.175652f
C5064 commonsourceibias.n306 gnd 0.067408f
C5065 commonsourceibias.n307 gnd 0.012292f
C5066 commonsourceibias.t0 gnd 0.172107f
C5067 commonsourceibias.n308 gnd 0.068671f
C5068 commonsourceibias.n309 gnd 0.009212f
C5069 commonsourceibias.t42 gnd 0.172107f
C5070 commonsourceibias.n310 gnd 0.007452f
C5071 commonsourceibias.n311 gnd 0.009212f
C5072 commonsourceibias.t10 gnd 0.172107f
C5073 commonsourceibias.n312 gnd 0.008893f
C5074 commonsourceibias.n313 gnd 0.009212f
C5075 commonsourceibias.t16 gnd 0.172107f
C5076 commonsourceibias.n314 gnd 0.00744f
C5077 commonsourceibias.n315 gnd 0.009212f
C5078 commonsourceibias.t30 gnd 0.172107f
C5079 commonsourceibias.t46 gnd 0.172107f
C5080 commonsourceibias.n316 gnd 0.068671f
C5081 commonsourceibias.n317 gnd 0.009212f
C5082 commonsourceibias.t14 gnd 0.172107f
C5083 commonsourceibias.n318 gnd 0.068671f
C5084 commonsourceibias.n319 gnd 0.009212f
C5085 commonsourceibias.t38 gnd 0.172107f
C5086 commonsourceibias.n320 gnd 0.068671f
C5087 commonsourceibias.n321 gnd 0.046375f
C5088 commonsourceibias.t26 gnd 0.172107f
C5089 commonsourceibias.t4 gnd 0.194203f
C5090 commonsourceibias.n322 gnd 0.079692f
C5091 commonsourceibias.n323 gnd 0.082502f
C5092 commonsourceibias.n324 gnd 0.011354f
C5093 commonsourceibias.n325 gnd 0.012561f
C5094 commonsourceibias.n326 gnd 0.009212f
C5095 commonsourceibias.n327 gnd 0.009212f
C5096 commonsourceibias.n328 gnd 0.012479f
C5097 commonsourceibias.n329 gnd 0.007452f
C5098 commonsourceibias.n330 gnd 0.012633f
C5099 commonsourceibias.n331 gnd 0.009212f
C5100 commonsourceibias.n332 gnd 0.009212f
C5101 commonsourceibias.n333 gnd 0.01271f
C5102 commonsourceibias.n334 gnd 0.01096f
C5103 commonsourceibias.n335 gnd 0.008893f
C5104 commonsourceibias.n336 gnd 0.009212f
C5105 commonsourceibias.n337 gnd 0.009212f
C5106 commonsourceibias.n338 gnd 0.011268f
C5107 commonsourceibias.n339 gnd 0.012647f
C5108 commonsourceibias.n340 gnd 0.068671f
C5109 commonsourceibias.n341 gnd 0.012562f
C5110 commonsourceibias.n342 gnd 0.009212f
C5111 commonsourceibias.n343 gnd 0.009212f
C5112 commonsourceibias.n344 gnd 0.009212f
C5113 commonsourceibias.n345 gnd 0.012562f
C5114 commonsourceibias.n346 gnd 0.068671f
C5115 commonsourceibias.n347 gnd 0.012647f
C5116 commonsourceibias.t36 gnd 0.172107f
C5117 commonsourceibias.n348 gnd 0.068671f
C5118 commonsourceibias.n349 gnd 0.011268f
C5119 commonsourceibias.n350 gnd 0.009212f
C5120 commonsourceibias.n351 gnd 0.009212f
C5121 commonsourceibias.n352 gnd 0.009212f
C5122 commonsourceibias.n353 gnd 0.01096f
C5123 commonsourceibias.n354 gnd 0.01271f
C5124 commonsourceibias.n355 gnd 0.068671f
C5125 commonsourceibias.n356 gnd 0.012633f
C5126 commonsourceibias.n357 gnd 0.009212f
C5127 commonsourceibias.n358 gnd 0.009212f
C5128 commonsourceibias.n359 gnd 0.009212f
C5129 commonsourceibias.n360 gnd 0.012479f
C5130 commonsourceibias.n361 gnd 0.068671f
C5131 commonsourceibias.n362 gnd 0.012561f
C5132 commonsourceibias.n363 gnd 0.011354f
C5133 commonsourceibias.n364 gnd 0.009212f
C5134 commonsourceibias.n365 gnd 0.009212f
C5135 commonsourceibias.n366 gnd 0.009345f
C5136 commonsourceibias.n367 gnd 0.009661f
C5137 commonsourceibias.t12 gnd 0.186134f
C5138 commonsourceibias.n368 gnd 0.082165f
C5139 commonsourceibias.n369 gnd 0.09115f
C5140 commonsourceibias.t1 gnd 0.019878f
C5141 commonsourceibias.t13 gnd 0.019878f
C5142 commonsourceibias.n370 gnd 0.175652f
C5143 commonsourceibias.n371 gnd 0.151777f
C5144 commonsourceibias.t11 gnd 0.019878f
C5145 commonsourceibias.t43 gnd 0.019878f
C5146 commonsourceibias.n372 gnd 0.175652f
C5147 commonsourceibias.n373 gnd 0.080684f
C5148 commonsourceibias.t17 gnd 0.019878f
C5149 commonsourceibias.t37 gnd 0.019878f
C5150 commonsourceibias.n374 gnd 0.175652f
C5151 commonsourceibias.n375 gnd 0.067408f
C5152 commonsourceibias.n376 gnd 0.081623f
C5153 commonsourceibias.n377 gnd 0.066591f
C5154 commonsourceibias.n378 gnd 0.009168f
C5155 commonsourceibias.n379 gnd 0.012562f
C5156 commonsourceibias.n380 gnd 0.068671f
C5157 commonsourceibias.n381 gnd 0.012647f
C5158 commonsourceibias.t92 gnd 0.172107f
C5159 commonsourceibias.n382 gnd 0.068671f
C5160 commonsourceibias.n383 gnd 0.011268f
C5161 commonsourceibias.n384 gnd 0.009212f
C5162 commonsourceibias.n385 gnd 0.009212f
C5163 commonsourceibias.n386 gnd 0.009212f
C5164 commonsourceibias.n387 gnd 0.01096f
C5165 commonsourceibias.n388 gnd 0.01271f
C5166 commonsourceibias.n389 gnd 0.068671f
C5167 commonsourceibias.n390 gnd 0.012633f
C5168 commonsourceibias.n391 gnd 0.009212f
C5169 commonsourceibias.n392 gnd 0.009212f
C5170 commonsourceibias.n393 gnd 0.009212f
C5171 commonsourceibias.n394 gnd 0.012479f
C5172 commonsourceibias.n395 gnd 0.068671f
C5173 commonsourceibias.n396 gnd 0.012561f
C5174 commonsourceibias.n397 gnd 0.011354f
C5175 commonsourceibias.n398 gnd 0.009212f
C5176 commonsourceibias.n399 gnd 0.009212f
C5177 commonsourceibias.n400 gnd 0.009345f
C5178 commonsourceibias.n401 gnd 0.009661f
C5179 commonsourceibias.n402 gnd 0.082165f
C5180 commonsourceibias.n403 gnd 0.053193f
C5181 commonsourceibias.n404 gnd 0.012292f
C5182 commonsourceibias.t107 gnd 0.172107f
C5183 commonsourceibias.n405 gnd 0.068671f
C5184 commonsourceibias.n406 gnd 0.009212f
C5185 commonsourceibias.t51 gnd 0.172107f
C5186 commonsourceibias.n407 gnd 0.007452f
C5187 commonsourceibias.n408 gnd 0.009212f
C5188 commonsourceibias.t114 gnd 0.172107f
C5189 commonsourceibias.n409 gnd 0.008893f
C5190 commonsourceibias.n410 gnd 0.009212f
C5191 commonsourceibias.t50 gnd 0.172107f
C5192 commonsourceibias.n411 gnd 0.00744f
C5193 commonsourceibias.n412 gnd 0.009212f
C5194 commonsourceibias.t76 gnd 0.172107f
C5195 commonsourceibias.t105 gnd 0.172107f
C5196 commonsourceibias.n413 gnd 0.068671f
C5197 commonsourceibias.n414 gnd 0.009212f
C5198 commonsourceibias.t55 gnd 0.172107f
C5199 commonsourceibias.n415 gnd 0.068671f
C5200 commonsourceibias.n416 gnd 0.009212f
C5201 commonsourceibias.t75 gnd 0.172107f
C5202 commonsourceibias.n417 gnd 0.068671f
C5203 commonsourceibias.n418 gnd 0.046375f
C5204 commonsourceibias.t61 gnd 0.172107f
C5205 commonsourceibias.t54 gnd 0.194203f
C5206 commonsourceibias.n419 gnd 0.079692f
C5207 commonsourceibias.n420 gnd 0.082502f
C5208 commonsourceibias.n421 gnd 0.011354f
C5209 commonsourceibias.n422 gnd 0.012561f
C5210 commonsourceibias.n423 gnd 0.009212f
C5211 commonsourceibias.n424 gnd 0.009212f
C5212 commonsourceibias.n425 gnd 0.012479f
C5213 commonsourceibias.n426 gnd 0.007452f
C5214 commonsourceibias.n427 gnd 0.012633f
C5215 commonsourceibias.n428 gnd 0.009212f
C5216 commonsourceibias.n429 gnd 0.009212f
C5217 commonsourceibias.n430 gnd 0.01271f
C5218 commonsourceibias.n431 gnd 0.01096f
C5219 commonsourceibias.n432 gnd 0.008893f
C5220 commonsourceibias.n433 gnd 0.009212f
C5221 commonsourceibias.n434 gnd 0.009212f
C5222 commonsourceibias.n435 gnd 0.011268f
C5223 commonsourceibias.n436 gnd 0.012647f
C5224 commonsourceibias.n437 gnd 0.068671f
C5225 commonsourceibias.n438 gnd 0.012562f
C5226 commonsourceibias.n439 gnd 0.009212f
C5227 commonsourceibias.n440 gnd 0.009212f
C5228 commonsourceibias.n441 gnd 0.009212f
C5229 commonsourceibias.n442 gnd 0.012562f
C5230 commonsourceibias.n443 gnd 0.068671f
C5231 commonsourceibias.n444 gnd 0.012647f
C5232 commonsourceibias.t106 gnd 0.172107f
C5233 commonsourceibias.n445 gnd 0.068671f
C5234 commonsourceibias.n446 gnd 0.011268f
C5235 commonsourceibias.n447 gnd 0.009212f
C5236 commonsourceibias.n448 gnd 0.009212f
C5237 commonsourceibias.n449 gnd 0.009212f
C5238 commonsourceibias.n450 gnd 0.01096f
C5239 commonsourceibias.n451 gnd 0.01271f
C5240 commonsourceibias.n452 gnd 0.068671f
C5241 commonsourceibias.n453 gnd 0.012633f
C5242 commonsourceibias.n454 gnd 0.009212f
C5243 commonsourceibias.n455 gnd 0.009212f
C5244 commonsourceibias.n456 gnd 0.009212f
C5245 commonsourceibias.n457 gnd 0.012479f
C5246 commonsourceibias.n458 gnd 0.068671f
C5247 commonsourceibias.n459 gnd 0.012561f
C5248 commonsourceibias.n460 gnd 0.011354f
C5249 commonsourceibias.n461 gnd 0.009212f
C5250 commonsourceibias.n462 gnd 0.009212f
C5251 commonsourceibias.n463 gnd 0.009345f
C5252 commonsourceibias.n464 gnd 0.009661f
C5253 commonsourceibias.t112 gnd 0.186134f
C5254 commonsourceibias.n465 gnd 0.082165f
C5255 commonsourceibias.n466 gnd 0.027962f
C5256 commonsourceibias.n467 gnd 0.146988f
C5257 commonsourceibias.n468 gnd 0.012292f
C5258 commonsourceibias.t81 gnd 0.172107f
C5259 commonsourceibias.n469 gnd 0.068671f
C5260 commonsourceibias.n470 gnd 0.009212f
C5261 commonsourceibias.t91 gnd 0.172107f
C5262 commonsourceibias.n471 gnd 0.007452f
C5263 commonsourceibias.n472 gnd 0.009212f
C5264 commonsourceibias.t101 gnd 0.172107f
C5265 commonsourceibias.n473 gnd 0.008893f
C5266 commonsourceibias.n474 gnd 0.009212f
C5267 commonsourceibias.t85 gnd 0.172107f
C5268 commonsourceibias.n475 gnd 0.00744f
C5269 commonsourceibias.n476 gnd 0.009212f
C5270 commonsourceibias.t82 gnd 0.172107f
C5271 commonsourceibias.t62 gnd 0.172107f
C5272 commonsourceibias.n477 gnd 0.068671f
C5273 commonsourceibias.n478 gnd 0.009212f
C5274 commonsourceibias.t53 gnd 0.172107f
C5275 commonsourceibias.n479 gnd 0.068671f
C5276 commonsourceibias.n480 gnd 0.009212f
C5277 commonsourceibias.t78 gnd 0.172107f
C5278 commonsourceibias.n481 gnd 0.068671f
C5279 commonsourceibias.n482 gnd 0.046375f
C5280 commonsourceibias.t97 gnd 0.172107f
C5281 commonsourceibias.t113 gnd 0.194203f
C5282 commonsourceibias.n483 gnd 0.079692f
C5283 commonsourceibias.n484 gnd 0.082502f
C5284 commonsourceibias.n485 gnd 0.011354f
C5285 commonsourceibias.n486 gnd 0.012561f
C5286 commonsourceibias.n487 gnd 0.009212f
C5287 commonsourceibias.n488 gnd 0.009212f
C5288 commonsourceibias.n489 gnd 0.012479f
C5289 commonsourceibias.n490 gnd 0.007452f
C5290 commonsourceibias.n491 gnd 0.012633f
C5291 commonsourceibias.n492 gnd 0.009212f
C5292 commonsourceibias.n493 gnd 0.009212f
C5293 commonsourceibias.n494 gnd 0.01271f
C5294 commonsourceibias.n495 gnd 0.01096f
C5295 commonsourceibias.n496 gnd 0.008893f
C5296 commonsourceibias.n497 gnd 0.009212f
C5297 commonsourceibias.n498 gnd 0.009212f
C5298 commonsourceibias.n499 gnd 0.011268f
C5299 commonsourceibias.n500 gnd 0.012647f
C5300 commonsourceibias.n501 gnd 0.068671f
C5301 commonsourceibias.n502 gnd 0.012562f
C5302 commonsourceibias.n503 gnd 0.009212f
C5303 commonsourceibias.n504 gnd 0.009212f
C5304 commonsourceibias.n505 gnd 0.009212f
C5305 commonsourceibias.n506 gnd 0.012562f
C5306 commonsourceibias.n507 gnd 0.068671f
C5307 commonsourceibias.n508 gnd 0.012647f
C5308 commonsourceibias.t74 gnd 0.172107f
C5309 commonsourceibias.n509 gnd 0.068671f
C5310 commonsourceibias.n510 gnd 0.011268f
C5311 commonsourceibias.n511 gnd 0.009212f
C5312 commonsourceibias.n512 gnd 0.009212f
C5313 commonsourceibias.n513 gnd 0.009212f
C5314 commonsourceibias.n514 gnd 0.01096f
C5315 commonsourceibias.n515 gnd 0.01271f
C5316 commonsourceibias.n516 gnd 0.068671f
C5317 commonsourceibias.n517 gnd 0.012633f
C5318 commonsourceibias.n518 gnd 0.009212f
C5319 commonsourceibias.n519 gnd 0.009212f
C5320 commonsourceibias.n520 gnd 0.009212f
C5321 commonsourceibias.n521 gnd 0.012479f
C5322 commonsourceibias.n522 gnd 0.068671f
C5323 commonsourceibias.n523 gnd 0.012561f
C5324 commonsourceibias.n524 gnd 0.011354f
C5325 commonsourceibias.n525 gnd 0.009212f
C5326 commonsourceibias.n526 gnd 0.009212f
C5327 commonsourceibias.n527 gnd 0.009345f
C5328 commonsourceibias.n528 gnd 0.009661f
C5329 commonsourceibias.t63 gnd 0.186134f
C5330 commonsourceibias.n529 gnd 0.082165f
C5331 commonsourceibias.n530 gnd 0.027962f
C5332 commonsourceibias.n531 gnd 0.194173f
C5333 commonsourceibias.n532 gnd 4.69557f
.ends

