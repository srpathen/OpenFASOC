* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t31 plus.t0 drain_left.t8 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X1 source.t14 minus.t0 drain_right.t15 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X2 a_n3110_n1488# a_n3110_n1488# a_n3110_n1488# a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=1
X3 drain_left.t1 plus.t1 source.t30 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X4 drain_left.t9 plus.t2 source.t29 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X5 drain_left.t2 plus.t3 source.t28 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X6 drain_right.t14 minus.t1 source.t2 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X7 source.t15 minus.t2 drain_right.t13 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
X8 drain_left.t3 plus.t4 source.t27 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X9 source.t26 plus.t5 drain_left.t0 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X10 source.t25 plus.t6 drain_left.t4 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X11 drain_right.t12 minus.t3 source.t1 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X12 drain_left.t10 plus.t7 source.t24 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X13 source.t23 plus.t8 drain_left.t13 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X14 drain_left.t14 plus.t9 source.t22 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X15 a_n3110_n1488# a_n3110_n1488# a_n3110_n1488# a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1
X16 drain_right.t11 minus.t4 source.t13 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X17 source.t10 minus.t5 drain_right.t10 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X18 source.t21 plus.t10 drain_left.t15 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X19 drain_right.t9 minus.t6 source.t6 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X20 source.t9 minus.t7 drain_right.t8 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X21 drain_right.t7 minus.t8 source.t12 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X22 a_n3110_n1488# a_n3110_n1488# a_n3110_n1488# a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1
X23 drain_left.t5 plus.t11 source.t20 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X24 source.t19 plus.t12 drain_left.t11 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
X25 drain_right.t6 minus.t9 source.t4 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X26 a_n3110_n1488# a_n3110_n1488# a_n3110_n1488# a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1
X27 drain_left.t6 plus.t13 source.t18 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X28 source.t11 minus.t10 drain_right.t5 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X29 source.t17 plus.t14 drain_left.t12 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X30 source.t5 minus.t11 drain_right.t4 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X31 source.t16 plus.t15 drain_left.t7 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
X32 source.t7 minus.t12 drain_right.t3 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X33 drain_right.t2 minus.t13 source.t8 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X34 drain_right.t1 minus.t14 source.t3 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X35 source.t0 minus.t15 drain_right.t0 a_n3110_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
R0 plus.n10 plus.n7 161.3
R1 plus.n12 plus.n11 161.3
R2 plus.n13 plus.n6 161.3
R3 plus.n16 plus.n15 161.3
R4 plus.n17 plus.n5 161.3
R5 plus.n19 plus.n18 161.3
R6 plus.n21 plus.n4 161.3
R7 plus.n24 plus.n23 161.3
R8 plus.n25 plus.n3 161.3
R9 plus.n27 plus.n26 161.3
R10 plus.n28 plus.n2 161.3
R11 plus.n31 plus.n30 161.3
R12 plus.n32 plus.n1 161.3
R13 plus.n34 plus.n33 161.3
R14 plus.n36 plus.n0 161.3
R15 plus.n50 plus.n47 161.3
R16 plus.n52 plus.n51 161.3
R17 plus.n53 plus.n46 161.3
R18 plus.n56 plus.n55 161.3
R19 plus.n57 plus.n45 161.3
R20 plus.n59 plus.n58 161.3
R21 plus.n61 plus.n43 161.3
R22 plus.n63 plus.n62 161.3
R23 plus.n64 plus.n42 161.3
R24 plus.n66 plus.n65 161.3
R25 plus.n67 plus.n41 161.3
R26 plus.n70 plus.n69 161.3
R27 plus.n71 plus.n40 161.3
R28 plus.n73 plus.n72 161.3
R29 plus.n75 plus.n39 161.3
R30 plus.n9 plus.t15 125.856
R31 plus.n49 plus.t9 125.856
R32 plus.n37 plus.t7 111.584
R33 plus.n76 plus.t12 111.584
R34 plus.n38 plus.n37 80.6037
R35 plus.n77 plus.n76 80.6037
R36 plus.n35 plus.t10 72.3005
R37 plus.n29 plus.t4 72.3005
R38 plus.n22 plus.t8 72.3005
R39 plus.n20 plus.t2 72.3005
R40 plus.n14 plus.t0 72.3005
R41 plus.n8 plus.t1 72.3005
R42 plus.n74 plus.t3 72.3005
R43 plus.n68 plus.t6 72.3005
R44 plus.n44 plus.t13 72.3005
R45 plus.n60 plus.t14 72.3005
R46 plus.n54 plus.t11 72.3005
R47 plus.n48 plus.t5 72.3005
R48 plus.n23 plus.n21 56.5617
R49 plus.n62 plus.n61 56.5617
R50 plus.n37 plus.n36 51.8893
R51 plus.n76 plus.n75 51.8893
R52 plus.n9 plus.n8 49.3649
R53 plus.n49 plus.n48 49.3649
R54 plus.n30 plus.n1 49.296
R55 plus.n13 plus.n12 49.296
R56 plus.n69 plus.n40 49.296
R57 plus.n53 plus.n52 49.296
R58 plus.n28 plus.n27 48.3272
R59 plus.n15 plus.n5 48.3272
R60 plus.n67 plus.n66 48.3272
R61 plus.n55 plus.n45 48.3272
R62 plus.n10 plus.n9 44.557
R63 plus.n50 plus.n49 44.557
R64 plus.n27 plus.n3 32.8269
R65 plus.n19 plus.n5 32.8269
R66 plus.n66 plus.n42 32.8269
R67 plus.n59 plus.n45 32.8269
R68 plus.n34 plus.n1 31.8581
R69 plus.n12 plus.n7 31.8581
R70 plus.n73 plus.n40 31.8581
R71 plus.n52 plus.n47 31.8581
R72 plus plus.n77 31.7192
R73 plus.n36 plus.n35 20.9036
R74 plus.n75 plus.n74 20.9036
R75 plus.n23 plus.n22 20.4117
R76 plus.n21 plus.n20 20.4117
R77 plus.n62 plus.n44 20.4117
R78 plus.n61 plus.n60 20.4117
R79 plus.n30 plus.n29 12.5423
R80 plus.n14 plus.n13 12.5423
R81 plus.n69 plus.n68 12.5423
R82 plus.n54 plus.n53 12.5423
R83 plus.n29 plus.n28 12.0505
R84 plus.n15 plus.n14 12.0505
R85 plus.n68 plus.n67 12.0505
R86 plus.n55 plus.n54 12.0505
R87 plus plus.n38 9.08049
R88 plus.n22 plus.n3 4.18111
R89 plus.n20 plus.n19 4.18111
R90 plus.n44 plus.n42 4.18111
R91 plus.n60 plus.n59 4.18111
R92 plus.n35 plus.n34 3.68928
R93 plus.n8 plus.n7 3.68928
R94 plus.n74 plus.n73 3.68928
R95 plus.n48 plus.n47 3.68928
R96 plus.n38 plus.n0 0.285035
R97 plus.n77 plus.n39 0.285035
R98 plus.n11 plus.n10 0.189894
R99 plus.n11 plus.n6 0.189894
R100 plus.n16 plus.n6 0.189894
R101 plus.n17 plus.n16 0.189894
R102 plus.n18 plus.n17 0.189894
R103 plus.n18 plus.n4 0.189894
R104 plus.n24 plus.n4 0.189894
R105 plus.n25 plus.n24 0.189894
R106 plus.n26 plus.n25 0.189894
R107 plus.n26 plus.n2 0.189894
R108 plus.n31 plus.n2 0.189894
R109 plus.n32 plus.n31 0.189894
R110 plus.n33 plus.n32 0.189894
R111 plus.n33 plus.n0 0.189894
R112 plus.n72 plus.n39 0.189894
R113 plus.n72 plus.n71 0.189894
R114 plus.n71 plus.n70 0.189894
R115 plus.n70 plus.n41 0.189894
R116 plus.n65 plus.n41 0.189894
R117 plus.n65 plus.n64 0.189894
R118 plus.n64 plus.n63 0.189894
R119 plus.n63 plus.n43 0.189894
R120 plus.n58 plus.n43 0.189894
R121 plus.n58 plus.n57 0.189894
R122 plus.n57 plus.n56 0.189894
R123 plus.n56 plus.n46 0.189894
R124 plus.n51 plus.n46 0.189894
R125 plus.n51 plus.n50 0.189894
R126 drain_left.n9 drain_left.n7 80.9197
R127 drain_left.n5 drain_left.n3 80.9196
R128 drain_left.n2 drain_left.n0 80.9196
R129 drain_left.n13 drain_left.n12 79.7731
R130 drain_left.n11 drain_left.n10 79.7731
R131 drain_left.n9 drain_left.n8 79.7731
R132 drain_left.n5 drain_left.n4 79.773
R133 drain_left.n2 drain_left.n1 79.773
R134 drain_left drain_left.n6 28.0015
R135 drain_left drain_left.n13 6.79977
R136 drain_left.n3 drain_left.t0 6.6005
R137 drain_left.n3 drain_left.t14 6.6005
R138 drain_left.n4 drain_left.t12 6.6005
R139 drain_left.n4 drain_left.t5 6.6005
R140 drain_left.n1 drain_left.t4 6.6005
R141 drain_left.n1 drain_left.t6 6.6005
R142 drain_left.n0 drain_left.t11 6.6005
R143 drain_left.n0 drain_left.t2 6.6005
R144 drain_left.n12 drain_left.t15 6.6005
R145 drain_left.n12 drain_left.t10 6.6005
R146 drain_left.n10 drain_left.t13 6.6005
R147 drain_left.n10 drain_left.t3 6.6005
R148 drain_left.n8 drain_left.t8 6.6005
R149 drain_left.n8 drain_left.t9 6.6005
R150 drain_left.n7 drain_left.t7 6.6005
R151 drain_left.n7 drain_left.t1 6.6005
R152 drain_left.n11 drain_left.n9 1.14705
R153 drain_left.n13 drain_left.n11 1.14705
R154 drain_left.n6 drain_left.n5 0.51843
R155 drain_left.n6 drain_left.n2 0.51843
R156 source.n0 source.t24 69.6943
R157 source.n7 source.t16 69.6943
R158 source.n8 source.t12 69.6943
R159 source.n15 source.t15 69.6943
R160 source.n31 source.t6 69.6942
R161 source.n24 source.t0 69.6942
R162 source.n23 source.t22 69.6942
R163 source.n16 source.t19 69.6942
R164 source.n2 source.n1 63.0943
R165 source.n4 source.n3 63.0943
R166 source.n6 source.n5 63.0943
R167 source.n10 source.n9 63.0943
R168 source.n12 source.n11 63.0943
R169 source.n14 source.n13 63.0943
R170 source.n30 source.n29 63.0942
R171 source.n28 source.n27 63.0942
R172 source.n26 source.n25 63.0942
R173 source.n22 source.n21 63.0942
R174 source.n20 source.n19 63.0942
R175 source.n18 source.n17 63.0942
R176 source.n16 source.n15 15.6161
R177 source.n32 source.n0 9.77989
R178 source.n29 source.t3 6.6005
R179 source.n29 source.t7 6.6005
R180 source.n27 source.t13 6.6005
R181 source.n27 source.t9 6.6005
R182 source.n25 source.t8 6.6005
R183 source.n25 source.t10 6.6005
R184 source.n21 source.t20 6.6005
R185 source.n21 source.t26 6.6005
R186 source.n19 source.t18 6.6005
R187 source.n19 source.t17 6.6005
R188 source.n17 source.t28 6.6005
R189 source.n17 source.t25 6.6005
R190 source.n1 source.t27 6.6005
R191 source.n1 source.t21 6.6005
R192 source.n3 source.t29 6.6005
R193 source.n3 source.t23 6.6005
R194 source.n5 source.t30 6.6005
R195 source.n5 source.t31 6.6005
R196 source.n9 source.t4 6.6005
R197 source.n9 source.t11 6.6005
R198 source.n11 source.t2 6.6005
R199 source.n11 source.t5 6.6005
R200 source.n13 source.t1 6.6005
R201 source.n13 source.t14 6.6005
R202 source.n32 source.n31 5.83671
R203 source.n15 source.n14 1.14705
R204 source.n14 source.n12 1.14705
R205 source.n12 source.n10 1.14705
R206 source.n10 source.n8 1.14705
R207 source.n7 source.n6 1.14705
R208 source.n6 source.n4 1.14705
R209 source.n4 source.n2 1.14705
R210 source.n2 source.n0 1.14705
R211 source.n18 source.n16 1.14705
R212 source.n20 source.n18 1.14705
R213 source.n22 source.n20 1.14705
R214 source.n23 source.n22 1.14705
R215 source.n26 source.n24 1.14705
R216 source.n28 source.n26 1.14705
R217 source.n30 source.n28 1.14705
R218 source.n31 source.n30 1.14705
R219 source.n8 source.n7 0.470328
R220 source.n24 source.n23 0.470328
R221 source source.n32 0.188
R222 minus.n36 minus.n0 161.3
R223 minus.n34 minus.n33 161.3
R224 minus.n32 minus.n1 161.3
R225 minus.n31 minus.n30 161.3
R226 minus.n28 minus.n2 161.3
R227 minus.n27 minus.n26 161.3
R228 minus.n25 minus.n3 161.3
R229 minus.n24 minus.n23 161.3
R230 minus.n22 minus.n4 161.3
R231 minus.n20 minus.n19 161.3
R232 minus.n18 minus.n6 161.3
R233 minus.n17 minus.n16 161.3
R234 minus.n14 minus.n7 161.3
R235 minus.n13 minus.n12 161.3
R236 minus.n11 minus.n8 161.3
R237 minus.n75 minus.n39 161.3
R238 minus.n73 minus.n72 161.3
R239 minus.n71 minus.n40 161.3
R240 minus.n70 minus.n69 161.3
R241 minus.n67 minus.n41 161.3
R242 minus.n66 minus.n65 161.3
R243 minus.n64 minus.n42 161.3
R244 minus.n63 minus.n62 161.3
R245 minus.n60 minus.n43 161.3
R246 minus.n58 minus.n57 161.3
R247 minus.n56 minus.n44 161.3
R248 minus.n55 minus.n54 161.3
R249 minus.n52 minus.n45 161.3
R250 minus.n51 minus.n50 161.3
R251 minus.n49 minus.n46 161.3
R252 minus.n10 minus.t8 125.856
R253 minus.n48 minus.t15 125.856
R254 minus.n37 minus.t2 111.584
R255 minus.n76 minus.t6 111.584
R256 minus.n38 minus.n37 80.6037
R257 minus.n77 minus.n76 80.6037
R258 minus.n9 minus.t10 72.3005
R259 minus.n15 minus.t9 72.3005
R260 minus.n21 minus.t11 72.3005
R261 minus.n5 minus.t1 72.3005
R262 minus.n29 minus.t0 72.3005
R263 minus.n35 minus.t3 72.3005
R264 minus.n47 minus.t13 72.3005
R265 minus.n53 minus.t5 72.3005
R266 minus.n59 minus.t4 72.3005
R267 minus.n61 minus.t7 72.3005
R268 minus.n68 minus.t14 72.3005
R269 minus.n74 minus.t12 72.3005
R270 minus.n23 minus.n22 56.5617
R271 minus.n62 minus.n60 56.5617
R272 minus.n37 minus.n36 51.8893
R273 minus.n76 minus.n75 51.8893
R274 minus.n10 minus.n9 49.3649
R275 minus.n48 minus.n47 49.3649
R276 minus.n14 minus.n13 49.296
R277 minus.n30 minus.n1 49.296
R278 minus.n52 minus.n51 49.296
R279 minus.n69 minus.n40 49.296
R280 minus.n16 minus.n6 48.3272
R281 minus.n28 minus.n27 48.3272
R282 minus.n54 minus.n44 48.3272
R283 minus.n67 minus.n66 48.3272
R284 minus.n11 minus.n10 44.557
R285 minus.n49 minus.n48 44.557
R286 minus.n78 minus.n38 34.429
R287 minus.n20 minus.n6 32.8269
R288 minus.n27 minus.n3 32.8269
R289 minus.n58 minus.n44 32.8269
R290 minus.n66 minus.n42 32.8269
R291 minus.n13 minus.n8 31.8581
R292 minus.n34 minus.n1 31.8581
R293 minus.n51 minus.n46 31.8581
R294 minus.n73 minus.n40 31.8581
R295 minus.n36 minus.n35 20.9036
R296 minus.n75 minus.n74 20.9036
R297 minus.n22 minus.n21 20.4117
R298 minus.n23 minus.n5 20.4117
R299 minus.n60 minus.n59 20.4117
R300 minus.n62 minus.n61 20.4117
R301 minus.n15 minus.n14 12.5423
R302 minus.n30 minus.n29 12.5423
R303 minus.n53 minus.n52 12.5423
R304 minus.n69 minus.n68 12.5423
R305 minus.n16 minus.n15 12.0505
R306 minus.n29 minus.n28 12.0505
R307 minus.n54 minus.n53 12.0505
R308 minus.n68 minus.n67 12.0505
R309 minus.n78 minus.n77 6.84564
R310 minus.n21 minus.n20 4.18111
R311 minus.n5 minus.n3 4.18111
R312 minus.n59 minus.n58 4.18111
R313 minus.n61 minus.n42 4.18111
R314 minus.n9 minus.n8 3.68928
R315 minus.n35 minus.n34 3.68928
R316 minus.n47 minus.n46 3.68928
R317 minus.n74 minus.n73 3.68928
R318 minus.n38 minus.n0 0.285035
R319 minus.n77 minus.n39 0.285035
R320 minus.n33 minus.n0 0.189894
R321 minus.n33 minus.n32 0.189894
R322 minus.n32 minus.n31 0.189894
R323 minus.n31 minus.n2 0.189894
R324 minus.n26 minus.n2 0.189894
R325 minus.n26 minus.n25 0.189894
R326 minus.n25 minus.n24 0.189894
R327 minus.n24 minus.n4 0.189894
R328 minus.n19 minus.n4 0.189894
R329 minus.n19 minus.n18 0.189894
R330 minus.n18 minus.n17 0.189894
R331 minus.n17 minus.n7 0.189894
R332 minus.n12 minus.n7 0.189894
R333 minus.n12 minus.n11 0.189894
R334 minus.n50 minus.n49 0.189894
R335 minus.n50 minus.n45 0.189894
R336 minus.n55 minus.n45 0.189894
R337 minus.n56 minus.n55 0.189894
R338 minus.n57 minus.n56 0.189894
R339 minus.n57 minus.n43 0.189894
R340 minus.n63 minus.n43 0.189894
R341 minus.n64 minus.n63 0.189894
R342 minus.n65 minus.n64 0.189894
R343 minus.n65 minus.n41 0.189894
R344 minus.n70 minus.n41 0.189894
R345 minus.n71 minus.n70 0.189894
R346 minus.n72 minus.n71 0.189894
R347 minus.n72 minus.n39 0.189894
R348 minus minus.n78 0.188
R349 drain_right.n9 drain_right.n7 80.9197
R350 drain_right.n5 drain_right.n3 80.9196
R351 drain_right.n2 drain_right.n0 80.9196
R352 drain_right.n9 drain_right.n8 79.7731
R353 drain_right.n11 drain_right.n10 79.7731
R354 drain_right.n13 drain_right.n12 79.7731
R355 drain_right.n5 drain_right.n4 79.773
R356 drain_right.n2 drain_right.n1 79.773
R357 drain_right drain_right.n6 27.4483
R358 drain_right drain_right.n13 6.79977
R359 drain_right.n3 drain_right.t3 6.6005
R360 drain_right.n3 drain_right.t9 6.6005
R361 drain_right.n4 drain_right.t8 6.6005
R362 drain_right.n4 drain_right.t1 6.6005
R363 drain_right.n1 drain_right.t10 6.6005
R364 drain_right.n1 drain_right.t11 6.6005
R365 drain_right.n0 drain_right.t0 6.6005
R366 drain_right.n0 drain_right.t2 6.6005
R367 drain_right.n7 drain_right.t5 6.6005
R368 drain_right.n7 drain_right.t7 6.6005
R369 drain_right.n8 drain_right.t4 6.6005
R370 drain_right.n8 drain_right.t6 6.6005
R371 drain_right.n10 drain_right.t15 6.6005
R372 drain_right.n10 drain_right.t14 6.6005
R373 drain_right.n12 drain_right.t13 6.6005
R374 drain_right.n12 drain_right.t12 6.6005
R375 drain_right.n13 drain_right.n11 1.14705
R376 drain_right.n11 drain_right.n9 1.14705
R377 drain_right.n6 drain_right.n5 0.51843
R378 drain_right.n6 drain_right.n2 0.51843
C0 drain_right minus 3.52274f
C1 source drain_left 7.19295f
C2 drain_left plus 3.83344f
C3 drain_left drain_right 1.64323f
C4 drain_left minus 0.179283f
C5 source plus 4.31017f
C6 source drain_right 7.19684f
C7 source minus 4.29618f
C8 plus drain_right 0.474553f
C9 plus minus 5.35961f
C10 drain_right a_n3110_n1488# 5.58845f
C11 drain_left a_n3110_n1488# 6.03491f
C12 source a_n3110_n1488# 4.162623f
C13 minus a_n3110_n1488# 11.742491f
C14 plus a_n3110_n1488# 13.05495f
C15 drain_right.t0 a_n3110_n1488# 0.060461f
C16 drain_right.t2 a_n3110_n1488# 0.060461f
C17 drain_right.n0 a_n3110_n1488# 0.441744f
C18 drain_right.t10 a_n3110_n1488# 0.060461f
C19 drain_right.t11 a_n3110_n1488# 0.060461f
C20 drain_right.n1 a_n3110_n1488# 0.436036f
C21 drain_right.n2 a_n3110_n1488# 0.739232f
C22 drain_right.t3 a_n3110_n1488# 0.060461f
C23 drain_right.t9 a_n3110_n1488# 0.060461f
C24 drain_right.n3 a_n3110_n1488# 0.441744f
C25 drain_right.t8 a_n3110_n1488# 0.060461f
C26 drain_right.t1 a_n3110_n1488# 0.060461f
C27 drain_right.n4 a_n3110_n1488# 0.436036f
C28 drain_right.n5 a_n3110_n1488# 0.739232f
C29 drain_right.n6 a_n3110_n1488# 1.08547f
C30 drain_right.t5 a_n3110_n1488# 0.060461f
C31 drain_right.t7 a_n3110_n1488# 0.060461f
C32 drain_right.n7 a_n3110_n1488# 0.441746f
C33 drain_right.t4 a_n3110_n1488# 0.060461f
C34 drain_right.t6 a_n3110_n1488# 0.060461f
C35 drain_right.n8 a_n3110_n1488# 0.436038f
C36 drain_right.n9 a_n3110_n1488# 0.789745f
C37 drain_right.t15 a_n3110_n1488# 0.060461f
C38 drain_right.t14 a_n3110_n1488# 0.060461f
C39 drain_right.n10 a_n3110_n1488# 0.436038f
C40 drain_right.n11 a_n3110_n1488# 0.392591f
C41 drain_right.t13 a_n3110_n1488# 0.060461f
C42 drain_right.t12 a_n3110_n1488# 0.060461f
C43 drain_right.n12 a_n3110_n1488# 0.436038f
C44 drain_right.n13 a_n3110_n1488# 0.627258f
C45 minus.n0 a_n3110_n1488# 0.050579f
C46 minus.t3 a_n3110_n1488# 0.283269f
C47 minus.n1 a_n3110_n1488# 0.034717f
C48 minus.n2 a_n3110_n1488# 0.037904f
C49 minus.t0 a_n3110_n1488# 0.283269f
C50 minus.n3 a_n3110_n1488# 0.047234f
C51 minus.n4 a_n3110_n1488# 0.037904f
C52 minus.t1 a_n3110_n1488# 0.283269f
C53 minus.n5 a_n3110_n1488# 0.140926f
C54 minus.t11 a_n3110_n1488# 0.283269f
C55 minus.n6 a_n3110_n1488# 0.033824f
C56 minus.n7 a_n3110_n1488# 0.037904f
C57 minus.t9 a_n3110_n1488# 0.283269f
C58 minus.n8 a_n3110_n1488# 0.046335f
C59 minus.t8 a_n3110_n1488# 0.363436f
C60 minus.t10 a_n3110_n1488# 0.283269f
C61 minus.n9 a_n3110_n1488# 0.168364f
C62 minus.n10 a_n3110_n1488# 0.196181f
C63 minus.n11 a_n3110_n1488# 0.158101f
C64 minus.n12 a_n3110_n1488# 0.037904f
C65 minus.n13 a_n3110_n1488# 0.034717f
C66 minus.n14 a_n3110_n1488# 0.052939f
C67 minus.n15 a_n3110_n1488# 0.140926f
C68 minus.n16 a_n3110_n1488# 0.052934f
C69 minus.n17 a_n3110_n1488# 0.037904f
C70 minus.n18 a_n3110_n1488# 0.037904f
C71 minus.n19 a_n3110_n1488# 0.037904f
C72 minus.n20 a_n3110_n1488# 0.047234f
C73 minus.n21 a_n3110_n1488# 0.140926f
C74 minus.n22 a_n3110_n1488# 0.049201f
C75 minus.n23 a_n3110_n1488# 0.049201f
C76 minus.n24 a_n3110_n1488# 0.037904f
C77 minus.n25 a_n3110_n1488# 0.037904f
C78 minus.n26 a_n3110_n1488# 0.037904f
C79 minus.n27 a_n3110_n1488# 0.033824f
C80 minus.n28 a_n3110_n1488# 0.052934f
C81 minus.n29 a_n3110_n1488# 0.140926f
C82 minus.n30 a_n3110_n1488# 0.052939f
C83 minus.n31 a_n3110_n1488# 0.037904f
C84 minus.n32 a_n3110_n1488# 0.037904f
C85 minus.n33 a_n3110_n1488# 0.037904f
C86 minus.n34 a_n3110_n1488# 0.046335f
C87 minus.n35 a_n3110_n1488# 0.140926f
C88 minus.n36 a_n3110_n1488# 0.047589f
C89 minus.t2 a_n3110_n1488# 0.340985f
C90 minus.n37 a_n3110_n1488# 0.19772f
C91 minus.n38 a_n3110_n1488# 1.26186f
C92 minus.n39 a_n3110_n1488# 0.050579f
C93 minus.t12 a_n3110_n1488# 0.283269f
C94 minus.n40 a_n3110_n1488# 0.034717f
C95 minus.n41 a_n3110_n1488# 0.037904f
C96 minus.t14 a_n3110_n1488# 0.283269f
C97 minus.n42 a_n3110_n1488# 0.047234f
C98 minus.n43 a_n3110_n1488# 0.037904f
C99 minus.t4 a_n3110_n1488# 0.283269f
C100 minus.n44 a_n3110_n1488# 0.033824f
C101 minus.n45 a_n3110_n1488# 0.037904f
C102 minus.t5 a_n3110_n1488# 0.283269f
C103 minus.n46 a_n3110_n1488# 0.046335f
C104 minus.t15 a_n3110_n1488# 0.363436f
C105 minus.t13 a_n3110_n1488# 0.283269f
C106 minus.n47 a_n3110_n1488# 0.168364f
C107 minus.n48 a_n3110_n1488# 0.196181f
C108 minus.n49 a_n3110_n1488# 0.158101f
C109 minus.n50 a_n3110_n1488# 0.037904f
C110 minus.n51 a_n3110_n1488# 0.034717f
C111 minus.n52 a_n3110_n1488# 0.052939f
C112 minus.n53 a_n3110_n1488# 0.140926f
C113 minus.n54 a_n3110_n1488# 0.052934f
C114 minus.n55 a_n3110_n1488# 0.037904f
C115 minus.n56 a_n3110_n1488# 0.037904f
C116 minus.n57 a_n3110_n1488# 0.037904f
C117 minus.n58 a_n3110_n1488# 0.047234f
C118 minus.n59 a_n3110_n1488# 0.140926f
C119 minus.n60 a_n3110_n1488# 0.049201f
C120 minus.t7 a_n3110_n1488# 0.283269f
C121 minus.n61 a_n3110_n1488# 0.140926f
C122 minus.n62 a_n3110_n1488# 0.049201f
C123 minus.n63 a_n3110_n1488# 0.037904f
C124 minus.n64 a_n3110_n1488# 0.037904f
C125 minus.n65 a_n3110_n1488# 0.037904f
C126 minus.n66 a_n3110_n1488# 0.033824f
C127 minus.n67 a_n3110_n1488# 0.052934f
C128 minus.n68 a_n3110_n1488# 0.140926f
C129 minus.n69 a_n3110_n1488# 0.052939f
C130 minus.n70 a_n3110_n1488# 0.037904f
C131 minus.n71 a_n3110_n1488# 0.037904f
C132 minus.n72 a_n3110_n1488# 0.037904f
C133 minus.n73 a_n3110_n1488# 0.046335f
C134 minus.n74 a_n3110_n1488# 0.140926f
C135 minus.n75 a_n3110_n1488# 0.047589f
C136 minus.t6 a_n3110_n1488# 0.340985f
C137 minus.n76 a_n3110_n1488# 0.19772f
C138 minus.n77 a_n3110_n1488# 0.2914f
C139 minus.n78 a_n3110_n1488# 1.51321f
C140 source.t24 a_n3110_n1488# 0.553537f
C141 source.n0 a_n3110_n1488# 0.851063f
C142 source.t27 a_n3110_n1488# 0.066661f
C143 source.t21 a_n3110_n1488# 0.066661f
C144 source.n1 a_n3110_n1488# 0.422666f
C145 source.n2 a_n3110_n1488# 0.452714f
C146 source.t29 a_n3110_n1488# 0.066661f
C147 source.t23 a_n3110_n1488# 0.066661f
C148 source.n3 a_n3110_n1488# 0.422666f
C149 source.n4 a_n3110_n1488# 0.452714f
C150 source.t30 a_n3110_n1488# 0.066661f
C151 source.t31 a_n3110_n1488# 0.066661f
C152 source.n5 a_n3110_n1488# 0.422666f
C153 source.n6 a_n3110_n1488# 0.452714f
C154 source.t16 a_n3110_n1488# 0.553537f
C155 source.n7 a_n3110_n1488# 0.442331f
C156 source.t12 a_n3110_n1488# 0.553537f
C157 source.n8 a_n3110_n1488# 0.442331f
C158 source.t4 a_n3110_n1488# 0.066661f
C159 source.t11 a_n3110_n1488# 0.066661f
C160 source.n9 a_n3110_n1488# 0.422666f
C161 source.n10 a_n3110_n1488# 0.452714f
C162 source.t2 a_n3110_n1488# 0.066661f
C163 source.t5 a_n3110_n1488# 0.066661f
C164 source.n11 a_n3110_n1488# 0.422666f
C165 source.n12 a_n3110_n1488# 0.452714f
C166 source.t1 a_n3110_n1488# 0.066661f
C167 source.t14 a_n3110_n1488# 0.066661f
C168 source.n13 a_n3110_n1488# 0.422666f
C169 source.n14 a_n3110_n1488# 0.452714f
C170 source.t15 a_n3110_n1488# 0.553537f
C171 source.n15 a_n3110_n1488# 1.15766f
C172 source.t19 a_n3110_n1488# 0.553534f
C173 source.n16 a_n3110_n1488# 1.15766f
C174 source.t28 a_n3110_n1488# 0.066661f
C175 source.t25 a_n3110_n1488# 0.066661f
C176 source.n17 a_n3110_n1488# 0.422663f
C177 source.n18 a_n3110_n1488# 0.452717f
C178 source.t18 a_n3110_n1488# 0.066661f
C179 source.t17 a_n3110_n1488# 0.066661f
C180 source.n19 a_n3110_n1488# 0.422663f
C181 source.n20 a_n3110_n1488# 0.452717f
C182 source.t20 a_n3110_n1488# 0.066661f
C183 source.t26 a_n3110_n1488# 0.066661f
C184 source.n21 a_n3110_n1488# 0.422663f
C185 source.n22 a_n3110_n1488# 0.452717f
C186 source.t22 a_n3110_n1488# 0.553534f
C187 source.n23 a_n3110_n1488# 0.442333f
C188 source.t0 a_n3110_n1488# 0.553534f
C189 source.n24 a_n3110_n1488# 0.442333f
C190 source.t8 a_n3110_n1488# 0.066661f
C191 source.t10 a_n3110_n1488# 0.066661f
C192 source.n25 a_n3110_n1488# 0.422663f
C193 source.n26 a_n3110_n1488# 0.452717f
C194 source.t13 a_n3110_n1488# 0.066661f
C195 source.t9 a_n3110_n1488# 0.066661f
C196 source.n27 a_n3110_n1488# 0.422663f
C197 source.n28 a_n3110_n1488# 0.452717f
C198 source.t3 a_n3110_n1488# 0.066661f
C199 source.t7 a_n3110_n1488# 0.066661f
C200 source.n29 a_n3110_n1488# 0.422663f
C201 source.n30 a_n3110_n1488# 0.452717f
C202 source.t6 a_n3110_n1488# 0.553534f
C203 source.n31 a_n3110_n1488# 0.643918f
C204 source.n32 a_n3110_n1488# 0.840339f
C205 drain_left.t11 a_n3110_n1488# 0.061582f
C206 drain_left.t2 a_n3110_n1488# 0.061582f
C207 drain_left.n0 a_n3110_n1488# 0.449935f
C208 drain_left.t4 a_n3110_n1488# 0.061582f
C209 drain_left.t6 a_n3110_n1488# 0.061582f
C210 drain_left.n1 a_n3110_n1488# 0.444121f
C211 drain_left.n2 a_n3110_n1488# 0.752938f
C212 drain_left.t0 a_n3110_n1488# 0.061582f
C213 drain_left.t14 a_n3110_n1488# 0.061582f
C214 drain_left.n3 a_n3110_n1488# 0.449935f
C215 drain_left.t12 a_n3110_n1488# 0.061582f
C216 drain_left.t5 a_n3110_n1488# 0.061582f
C217 drain_left.n4 a_n3110_n1488# 0.444121f
C218 drain_left.n5 a_n3110_n1488# 0.752938f
C219 drain_left.n6 a_n3110_n1488# 1.15634f
C220 drain_left.t7 a_n3110_n1488# 0.061582f
C221 drain_left.t1 a_n3110_n1488# 0.061582f
C222 drain_left.n7 a_n3110_n1488# 0.449937f
C223 drain_left.t8 a_n3110_n1488# 0.061582f
C224 drain_left.t9 a_n3110_n1488# 0.061582f
C225 drain_left.n8 a_n3110_n1488# 0.444123f
C226 drain_left.n9 a_n3110_n1488# 0.804387f
C227 drain_left.t13 a_n3110_n1488# 0.061582f
C228 drain_left.t3 a_n3110_n1488# 0.061582f
C229 drain_left.n10 a_n3110_n1488# 0.444123f
C230 drain_left.n11 a_n3110_n1488# 0.399869f
C231 drain_left.t15 a_n3110_n1488# 0.061582f
C232 drain_left.t10 a_n3110_n1488# 0.061582f
C233 drain_left.n12 a_n3110_n1488# 0.444123f
C234 drain_left.n13 a_n3110_n1488# 0.638888f
C235 plus.n0 a_n3110_n1488# 0.05203f
C236 plus.t7 a_n3110_n1488# 0.350771f
C237 plus.t10 a_n3110_n1488# 0.291399f
C238 plus.n1 a_n3110_n1488# 0.035714f
C239 plus.n2 a_n3110_n1488# 0.038992f
C240 plus.t4 a_n3110_n1488# 0.291399f
C241 plus.n3 a_n3110_n1488# 0.048589f
C242 plus.n4 a_n3110_n1488# 0.038992f
C243 plus.t2 a_n3110_n1488# 0.291399f
C244 plus.n5 a_n3110_n1488# 0.034794f
C245 plus.n6 a_n3110_n1488# 0.038992f
C246 plus.t0 a_n3110_n1488# 0.291399f
C247 plus.n7 a_n3110_n1488# 0.047665f
C248 plus.t1 a_n3110_n1488# 0.291399f
C249 plus.n8 a_n3110_n1488# 0.173196f
C250 plus.t15 a_n3110_n1488# 0.373866f
C251 plus.n9 a_n3110_n1488# 0.201812f
C252 plus.n10 a_n3110_n1488# 0.162639f
C253 plus.n11 a_n3110_n1488# 0.038992f
C254 plus.n12 a_n3110_n1488# 0.035714f
C255 plus.n13 a_n3110_n1488# 0.054459f
C256 plus.n14 a_n3110_n1488# 0.144971f
C257 plus.n15 a_n3110_n1488# 0.054453f
C258 plus.n16 a_n3110_n1488# 0.038992f
C259 plus.n17 a_n3110_n1488# 0.038992f
C260 plus.n18 a_n3110_n1488# 0.038992f
C261 plus.n19 a_n3110_n1488# 0.048589f
C262 plus.n20 a_n3110_n1488# 0.144971f
C263 plus.n21 a_n3110_n1488# 0.050613f
C264 plus.t8 a_n3110_n1488# 0.291399f
C265 plus.n22 a_n3110_n1488# 0.144971f
C266 plus.n23 a_n3110_n1488# 0.050613f
C267 plus.n24 a_n3110_n1488# 0.038992f
C268 plus.n25 a_n3110_n1488# 0.038992f
C269 plus.n26 a_n3110_n1488# 0.038992f
C270 plus.n27 a_n3110_n1488# 0.034794f
C271 plus.n28 a_n3110_n1488# 0.054453f
C272 plus.n29 a_n3110_n1488# 0.144971f
C273 plus.n30 a_n3110_n1488# 0.054459f
C274 plus.n31 a_n3110_n1488# 0.038992f
C275 plus.n32 a_n3110_n1488# 0.038992f
C276 plus.n33 a_n3110_n1488# 0.038992f
C277 plus.n34 a_n3110_n1488# 0.047665f
C278 plus.n35 a_n3110_n1488# 0.144971f
C279 plus.n36 a_n3110_n1488# 0.048954f
C280 plus.n37 a_n3110_n1488# 0.203395f
C281 plus.n38 a_n3110_n1488# 0.337904f
C282 plus.n39 a_n3110_n1488# 0.05203f
C283 plus.t12 a_n3110_n1488# 0.350771f
C284 plus.t3 a_n3110_n1488# 0.291399f
C285 plus.n40 a_n3110_n1488# 0.035714f
C286 plus.n41 a_n3110_n1488# 0.038992f
C287 plus.t6 a_n3110_n1488# 0.291399f
C288 plus.n42 a_n3110_n1488# 0.048589f
C289 plus.n43 a_n3110_n1488# 0.038992f
C290 plus.t13 a_n3110_n1488# 0.291399f
C291 plus.n44 a_n3110_n1488# 0.144971f
C292 plus.t14 a_n3110_n1488# 0.291399f
C293 plus.n45 a_n3110_n1488# 0.034794f
C294 plus.n46 a_n3110_n1488# 0.038992f
C295 plus.t11 a_n3110_n1488# 0.291399f
C296 plus.n47 a_n3110_n1488# 0.047665f
C297 plus.t9 a_n3110_n1488# 0.373866f
C298 plus.t5 a_n3110_n1488# 0.291399f
C299 plus.n48 a_n3110_n1488# 0.173196f
C300 plus.n49 a_n3110_n1488# 0.201812f
C301 plus.n50 a_n3110_n1488# 0.162639f
C302 plus.n51 a_n3110_n1488# 0.038992f
C303 plus.n52 a_n3110_n1488# 0.035714f
C304 plus.n53 a_n3110_n1488# 0.054459f
C305 plus.n54 a_n3110_n1488# 0.144971f
C306 plus.n55 a_n3110_n1488# 0.054453f
C307 plus.n56 a_n3110_n1488# 0.038992f
C308 plus.n57 a_n3110_n1488# 0.038992f
C309 plus.n58 a_n3110_n1488# 0.038992f
C310 plus.n59 a_n3110_n1488# 0.048589f
C311 plus.n60 a_n3110_n1488# 0.144971f
C312 plus.n61 a_n3110_n1488# 0.050613f
C313 plus.n62 a_n3110_n1488# 0.050613f
C314 plus.n63 a_n3110_n1488# 0.038992f
C315 plus.n64 a_n3110_n1488# 0.038992f
C316 plus.n65 a_n3110_n1488# 0.038992f
C317 plus.n66 a_n3110_n1488# 0.034794f
C318 plus.n67 a_n3110_n1488# 0.054453f
C319 plus.n68 a_n3110_n1488# 0.144971f
C320 plus.n69 a_n3110_n1488# 0.054459f
C321 plus.n70 a_n3110_n1488# 0.038992f
C322 plus.n71 a_n3110_n1488# 0.038992f
C323 plus.n72 a_n3110_n1488# 0.038992f
C324 plus.n73 a_n3110_n1488# 0.047665f
C325 plus.n74 a_n3110_n1488# 0.144971f
C326 plus.n75 a_n3110_n1488# 0.048954f
C327 plus.n76 a_n3110_n1488# 0.203395f
C328 plus.n77 a_n3110_n1488# 1.22047f
.ends

