* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t28 plus.t0 drain_left.t1 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X1 source.t0 minus.t0 drain_right.t15 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X2 drain_left.t10 plus.t1 source.t27 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X3 drain_left.t13 plus.t2 source.t26 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X4 drain_left.t7 plus.t3 source.t25 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X5 drain_right.t14 minus.t1 source.t11 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X6 drain_right.t13 minus.t2 source.t3 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X7 source.t1 minus.t3 drain_right.t12 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X8 drain_left.t6 plus.t4 source.t24 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X9 drain_right.t11 minus.t4 source.t7 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X10 drain_left.t5 plus.t5 source.t23 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X11 source.t22 plus.t6 drain_left.t4 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X12 drain_left.t14 plus.t7 source.t21 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X13 a_n3110_n2088# a_n3110_n2088# a_n3110_n2088# a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=1
X14 source.t20 plus.t8 drain_left.t8 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X15 source.t4 minus.t5 drain_right.t10 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X16 source.t19 plus.t9 drain_left.t3 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X17 source.t18 plus.t10 drain_left.t9 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X18 source.t17 plus.t11 drain_left.t11 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X19 drain_right.t9 minus.t6 source.t6 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X20 drain_left.t12 plus.t12 source.t16 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X21 source.t9 minus.t7 drain_right.t8 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X22 drain_right.t7 minus.t8 source.t31 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X23 a_n3110_n2088# a_n3110_n2088# a_n3110_n2088# a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X24 a_n3110_n2088# a_n3110_n2088# a_n3110_n2088# a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X25 source.t30 minus.t9 drain_right.t6 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X26 drain_right.t5 minus.t10 source.t12 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X27 drain_right.t4 minus.t11 source.t5 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X28 drain_right.t3 minus.t12 source.t8 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X29 drain_left.t0 plus.t13 source.t15 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X30 a_n3110_n2088# a_n3110_n2088# a_n3110_n2088# a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X31 source.t29 minus.t13 drain_right.t2 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X32 source.t10 minus.t14 drain_right.t1 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X33 source.t14 plus.t14 drain_left.t15 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X34 source.t2 minus.t15 drain_right.t0 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X35 source.t13 plus.t15 drain_left.t2 a_n3110_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
R0 plus.n9 plus.t15 198.156
R1 plus.n49 plus.t12 198.156
R2 plus.n37 plus.t5 183.883
R3 plus.n76 plus.t14 183.883
R4 plus.n10 plus.n7 161.3
R5 plus.n12 plus.n11 161.3
R6 plus.n13 plus.n6 161.3
R7 plus.n16 plus.n15 161.3
R8 plus.n17 plus.n5 161.3
R9 plus.n19 plus.n18 161.3
R10 plus.n21 plus.n4 161.3
R11 plus.n24 plus.n23 161.3
R12 plus.n25 plus.n3 161.3
R13 plus.n27 plus.n26 161.3
R14 plus.n28 plus.n2 161.3
R15 plus.n31 plus.n30 161.3
R16 plus.n32 plus.n1 161.3
R17 plus.n34 plus.n33 161.3
R18 plus.n36 plus.n0 161.3
R19 plus.n50 plus.n47 161.3
R20 plus.n52 plus.n51 161.3
R21 plus.n53 plus.n46 161.3
R22 plus.n56 plus.n55 161.3
R23 plus.n57 plus.n45 161.3
R24 plus.n59 plus.n58 161.3
R25 plus.n61 plus.n43 161.3
R26 plus.n63 plus.n62 161.3
R27 plus.n64 plus.n42 161.3
R28 plus.n66 plus.n65 161.3
R29 plus.n67 plus.n41 161.3
R30 plus.n70 plus.n69 161.3
R31 plus.n71 plus.n40 161.3
R32 plus.n73 plus.n72 161.3
R33 plus.n75 plus.n39 161.3
R34 plus.n35 plus.t8 144.601
R35 plus.n29 plus.t4 144.601
R36 plus.n22 plus.t6 144.601
R37 plus.n20 plus.t3 144.601
R38 plus.n14 plus.t0 144.601
R39 plus.n8 plus.t1 144.601
R40 plus.n74 plus.t7 144.601
R41 plus.n68 plus.t11 144.601
R42 plus.n44 plus.t2 144.601
R43 plus.n60 plus.t9 144.601
R44 plus.n54 plus.t13 144.601
R45 plus.n48 plus.t10 144.601
R46 plus.n38 plus.n37 80.6037
R47 plus.n77 plus.n76 80.6037
R48 plus.n23 plus.n21 56.5617
R49 plus.n62 plus.n61 56.5617
R50 plus.n37 plus.n36 51.8893
R51 plus.n76 plus.n75 51.8893
R52 plus.n9 plus.n8 49.3649
R53 plus.n49 plus.n48 49.3649
R54 plus.n30 plus.n1 49.296
R55 plus.n13 plus.n12 49.296
R56 plus.n69 plus.n40 49.296
R57 plus.n53 plus.n52 49.296
R58 plus.n28 plus.n27 48.3272
R59 plus.n15 plus.n5 48.3272
R60 plus.n67 plus.n66 48.3272
R61 plus.n55 plus.n45 48.3272
R62 plus.n10 plus.n9 44.557
R63 plus.n50 plus.n49 44.557
R64 plus plus.n77 32.8555
R65 plus.n27 plus.n3 32.8269
R66 plus.n19 plus.n5 32.8269
R67 plus.n66 plus.n42 32.8269
R68 plus.n59 plus.n45 32.8269
R69 plus.n34 plus.n1 31.8581
R70 plus.n12 plus.n7 31.8581
R71 plus.n73 plus.n40 31.8581
R72 plus.n52 plus.n47 31.8581
R73 plus.n36 plus.n35 20.9036
R74 plus.n75 plus.n74 20.9036
R75 plus.n23 plus.n22 20.4117
R76 plus.n21 plus.n20 20.4117
R77 plus.n62 plus.n44 20.4117
R78 plus.n61 plus.n60 20.4117
R79 plus.n30 plus.n29 12.5423
R80 plus.n14 plus.n13 12.5423
R81 plus.n69 plus.n68 12.5423
R82 plus.n54 plus.n53 12.5423
R83 plus.n29 plus.n28 12.0505
R84 plus.n15 plus.n14 12.0505
R85 plus.n68 plus.n67 12.0505
R86 plus.n55 plus.n54 12.0505
R87 plus plus.n38 10.2169
R88 plus.n22 plus.n3 4.18111
R89 plus.n20 plus.n19 4.18111
R90 plus.n44 plus.n42 4.18111
R91 plus.n60 plus.n59 4.18111
R92 plus.n35 plus.n34 3.68928
R93 plus.n8 plus.n7 3.68928
R94 plus.n74 plus.n73 3.68928
R95 plus.n48 plus.n47 3.68928
R96 plus.n38 plus.n0 0.285035
R97 plus.n77 plus.n39 0.285035
R98 plus.n11 plus.n10 0.189894
R99 plus.n11 plus.n6 0.189894
R100 plus.n16 plus.n6 0.189894
R101 plus.n17 plus.n16 0.189894
R102 plus.n18 plus.n17 0.189894
R103 plus.n18 plus.n4 0.189894
R104 plus.n24 plus.n4 0.189894
R105 plus.n25 plus.n24 0.189894
R106 plus.n26 plus.n25 0.189894
R107 plus.n26 plus.n2 0.189894
R108 plus.n31 plus.n2 0.189894
R109 plus.n32 plus.n31 0.189894
R110 plus.n33 plus.n32 0.189894
R111 plus.n33 plus.n0 0.189894
R112 plus.n72 plus.n39 0.189894
R113 plus.n72 plus.n71 0.189894
R114 plus.n71 plus.n70 0.189894
R115 plus.n70 plus.n41 0.189894
R116 plus.n65 plus.n41 0.189894
R117 plus.n65 plus.n64 0.189894
R118 plus.n64 plus.n63 0.189894
R119 plus.n63 plus.n43 0.189894
R120 plus.n58 plus.n43 0.189894
R121 plus.n58 plus.n57 0.189894
R122 plus.n57 plus.n56 0.189894
R123 plus.n56 plus.n46 0.189894
R124 plus.n51 plus.n46 0.189894
R125 plus.n51 plus.n50 0.189894
R126 drain_left.n9 drain_left.n7 68.3374
R127 drain_left.n5 drain_left.n3 68.3372
R128 drain_left.n2 drain_left.n0 68.3372
R129 drain_left.n11 drain_left.n10 67.1908
R130 drain_left.n9 drain_left.n8 67.1908
R131 drain_left.n13 drain_left.n12 67.1907
R132 drain_left.n5 drain_left.n4 67.1907
R133 drain_left.n2 drain_left.n1 67.1907
R134 drain_left drain_left.n6 30.2742
R135 drain_left drain_left.n13 6.79977
R136 drain_left.n3 drain_left.t9 3.3005
R137 drain_left.n3 drain_left.t12 3.3005
R138 drain_left.n4 drain_left.t3 3.3005
R139 drain_left.n4 drain_left.t0 3.3005
R140 drain_left.n1 drain_left.t11 3.3005
R141 drain_left.n1 drain_left.t13 3.3005
R142 drain_left.n0 drain_left.t15 3.3005
R143 drain_left.n0 drain_left.t14 3.3005
R144 drain_left.n12 drain_left.t8 3.3005
R145 drain_left.n12 drain_left.t5 3.3005
R146 drain_left.n10 drain_left.t4 3.3005
R147 drain_left.n10 drain_left.t6 3.3005
R148 drain_left.n8 drain_left.t1 3.3005
R149 drain_left.n8 drain_left.t7 3.3005
R150 drain_left.n7 drain_left.t2 3.3005
R151 drain_left.n7 drain_left.t10 3.3005
R152 drain_left.n11 drain_left.n9 1.14705
R153 drain_left.n13 drain_left.n11 1.14705
R154 drain_left.n6 drain_left.n5 0.51843
R155 drain_left.n6 drain_left.n2 0.51843
R156 source.n274 source.n248 289.615
R157 source.n236 source.n210 289.615
R158 source.n204 source.n178 289.615
R159 source.n166 source.n140 289.615
R160 source.n26 source.n0 289.615
R161 source.n64 source.n38 289.615
R162 source.n96 source.n70 289.615
R163 source.n134 source.n108 289.615
R164 source.n259 source.n258 185
R165 source.n256 source.n255 185
R166 source.n265 source.n264 185
R167 source.n267 source.n266 185
R168 source.n252 source.n251 185
R169 source.n273 source.n272 185
R170 source.n275 source.n274 185
R171 source.n221 source.n220 185
R172 source.n218 source.n217 185
R173 source.n227 source.n226 185
R174 source.n229 source.n228 185
R175 source.n214 source.n213 185
R176 source.n235 source.n234 185
R177 source.n237 source.n236 185
R178 source.n189 source.n188 185
R179 source.n186 source.n185 185
R180 source.n195 source.n194 185
R181 source.n197 source.n196 185
R182 source.n182 source.n181 185
R183 source.n203 source.n202 185
R184 source.n205 source.n204 185
R185 source.n151 source.n150 185
R186 source.n148 source.n147 185
R187 source.n157 source.n156 185
R188 source.n159 source.n158 185
R189 source.n144 source.n143 185
R190 source.n165 source.n164 185
R191 source.n167 source.n166 185
R192 source.n27 source.n26 185
R193 source.n25 source.n24 185
R194 source.n4 source.n3 185
R195 source.n19 source.n18 185
R196 source.n17 source.n16 185
R197 source.n8 source.n7 185
R198 source.n11 source.n10 185
R199 source.n65 source.n64 185
R200 source.n63 source.n62 185
R201 source.n42 source.n41 185
R202 source.n57 source.n56 185
R203 source.n55 source.n54 185
R204 source.n46 source.n45 185
R205 source.n49 source.n48 185
R206 source.n97 source.n96 185
R207 source.n95 source.n94 185
R208 source.n74 source.n73 185
R209 source.n89 source.n88 185
R210 source.n87 source.n86 185
R211 source.n78 source.n77 185
R212 source.n81 source.n80 185
R213 source.n135 source.n134 185
R214 source.n133 source.n132 185
R215 source.n112 source.n111 185
R216 source.n127 source.n126 185
R217 source.n125 source.n124 185
R218 source.n116 source.n115 185
R219 source.n119 source.n118 185
R220 source.t11 source.n257 147.661
R221 source.t30 source.n219 147.661
R222 source.t16 source.n187 147.661
R223 source.t14 source.n149 147.661
R224 source.t23 source.n9 147.661
R225 source.t13 source.n47 147.661
R226 source.t31 source.n79 147.661
R227 source.t1 source.n117 147.661
R228 source.n258 source.n255 104.615
R229 source.n265 source.n255 104.615
R230 source.n266 source.n265 104.615
R231 source.n266 source.n251 104.615
R232 source.n273 source.n251 104.615
R233 source.n274 source.n273 104.615
R234 source.n220 source.n217 104.615
R235 source.n227 source.n217 104.615
R236 source.n228 source.n227 104.615
R237 source.n228 source.n213 104.615
R238 source.n235 source.n213 104.615
R239 source.n236 source.n235 104.615
R240 source.n188 source.n185 104.615
R241 source.n195 source.n185 104.615
R242 source.n196 source.n195 104.615
R243 source.n196 source.n181 104.615
R244 source.n203 source.n181 104.615
R245 source.n204 source.n203 104.615
R246 source.n150 source.n147 104.615
R247 source.n157 source.n147 104.615
R248 source.n158 source.n157 104.615
R249 source.n158 source.n143 104.615
R250 source.n165 source.n143 104.615
R251 source.n166 source.n165 104.615
R252 source.n26 source.n25 104.615
R253 source.n25 source.n3 104.615
R254 source.n18 source.n3 104.615
R255 source.n18 source.n17 104.615
R256 source.n17 source.n7 104.615
R257 source.n10 source.n7 104.615
R258 source.n64 source.n63 104.615
R259 source.n63 source.n41 104.615
R260 source.n56 source.n41 104.615
R261 source.n56 source.n55 104.615
R262 source.n55 source.n45 104.615
R263 source.n48 source.n45 104.615
R264 source.n96 source.n95 104.615
R265 source.n95 source.n73 104.615
R266 source.n88 source.n73 104.615
R267 source.n88 source.n87 104.615
R268 source.n87 source.n77 104.615
R269 source.n80 source.n77 104.615
R270 source.n134 source.n133 104.615
R271 source.n133 source.n111 104.615
R272 source.n126 source.n111 104.615
R273 source.n126 source.n125 104.615
R274 source.n125 source.n115 104.615
R275 source.n118 source.n115 104.615
R276 source.n258 source.t11 52.3082
R277 source.n220 source.t30 52.3082
R278 source.n188 source.t16 52.3082
R279 source.n150 source.t14 52.3082
R280 source.n10 source.t23 52.3082
R281 source.n48 source.t13 52.3082
R282 source.n80 source.t31 52.3082
R283 source.n118 source.t1 52.3082
R284 source.n33 source.n32 50.512
R285 source.n35 source.n34 50.512
R286 source.n37 source.n36 50.512
R287 source.n103 source.n102 50.512
R288 source.n105 source.n104 50.512
R289 source.n107 source.n106 50.512
R290 source.n247 source.n246 50.5119
R291 source.n245 source.n244 50.5119
R292 source.n243 source.n242 50.5119
R293 source.n177 source.n176 50.5119
R294 source.n175 source.n174 50.5119
R295 source.n173 source.n172 50.5119
R296 source.n279 source.n278 32.1853
R297 source.n241 source.n240 32.1853
R298 source.n209 source.n208 32.1853
R299 source.n171 source.n170 32.1853
R300 source.n31 source.n30 32.1853
R301 source.n69 source.n68 32.1853
R302 source.n101 source.n100 32.1853
R303 source.n139 source.n138 32.1853
R304 source.n171 source.n139 17.8888
R305 source.n259 source.n257 15.6674
R306 source.n221 source.n219 15.6674
R307 source.n189 source.n187 15.6674
R308 source.n151 source.n149 15.6674
R309 source.n11 source.n9 15.6674
R310 source.n49 source.n47 15.6674
R311 source.n81 source.n79 15.6674
R312 source.n119 source.n117 15.6674
R313 source.n260 source.n256 12.8005
R314 source.n222 source.n218 12.8005
R315 source.n190 source.n186 12.8005
R316 source.n152 source.n148 12.8005
R317 source.n12 source.n8 12.8005
R318 source.n50 source.n46 12.8005
R319 source.n82 source.n78 12.8005
R320 source.n120 source.n116 12.8005
R321 source.n280 source.n31 12.0526
R322 source.n264 source.n263 12.0247
R323 source.n226 source.n225 12.0247
R324 source.n194 source.n193 12.0247
R325 source.n156 source.n155 12.0247
R326 source.n16 source.n15 12.0247
R327 source.n54 source.n53 12.0247
R328 source.n86 source.n85 12.0247
R329 source.n124 source.n123 12.0247
R330 source.n267 source.n254 11.249
R331 source.n229 source.n216 11.249
R332 source.n197 source.n184 11.249
R333 source.n159 source.n146 11.249
R334 source.n19 source.n6 11.249
R335 source.n57 source.n44 11.249
R336 source.n89 source.n76 11.249
R337 source.n127 source.n114 11.249
R338 source.n268 source.n252 10.4732
R339 source.n230 source.n214 10.4732
R340 source.n198 source.n182 10.4732
R341 source.n160 source.n144 10.4732
R342 source.n20 source.n4 10.4732
R343 source.n58 source.n42 10.4732
R344 source.n90 source.n74 10.4732
R345 source.n128 source.n112 10.4732
R346 source.n272 source.n271 9.69747
R347 source.n234 source.n233 9.69747
R348 source.n202 source.n201 9.69747
R349 source.n164 source.n163 9.69747
R350 source.n24 source.n23 9.69747
R351 source.n62 source.n61 9.69747
R352 source.n94 source.n93 9.69747
R353 source.n132 source.n131 9.69747
R354 source.n278 source.n277 9.45567
R355 source.n240 source.n239 9.45567
R356 source.n208 source.n207 9.45567
R357 source.n170 source.n169 9.45567
R358 source.n30 source.n29 9.45567
R359 source.n68 source.n67 9.45567
R360 source.n100 source.n99 9.45567
R361 source.n138 source.n137 9.45567
R362 source.n277 source.n276 9.3005
R363 source.n250 source.n249 9.3005
R364 source.n271 source.n270 9.3005
R365 source.n269 source.n268 9.3005
R366 source.n254 source.n253 9.3005
R367 source.n263 source.n262 9.3005
R368 source.n261 source.n260 9.3005
R369 source.n239 source.n238 9.3005
R370 source.n212 source.n211 9.3005
R371 source.n233 source.n232 9.3005
R372 source.n231 source.n230 9.3005
R373 source.n216 source.n215 9.3005
R374 source.n225 source.n224 9.3005
R375 source.n223 source.n222 9.3005
R376 source.n207 source.n206 9.3005
R377 source.n180 source.n179 9.3005
R378 source.n201 source.n200 9.3005
R379 source.n199 source.n198 9.3005
R380 source.n184 source.n183 9.3005
R381 source.n193 source.n192 9.3005
R382 source.n191 source.n190 9.3005
R383 source.n169 source.n168 9.3005
R384 source.n142 source.n141 9.3005
R385 source.n163 source.n162 9.3005
R386 source.n161 source.n160 9.3005
R387 source.n146 source.n145 9.3005
R388 source.n155 source.n154 9.3005
R389 source.n153 source.n152 9.3005
R390 source.n29 source.n28 9.3005
R391 source.n2 source.n1 9.3005
R392 source.n23 source.n22 9.3005
R393 source.n21 source.n20 9.3005
R394 source.n6 source.n5 9.3005
R395 source.n15 source.n14 9.3005
R396 source.n13 source.n12 9.3005
R397 source.n67 source.n66 9.3005
R398 source.n40 source.n39 9.3005
R399 source.n61 source.n60 9.3005
R400 source.n59 source.n58 9.3005
R401 source.n44 source.n43 9.3005
R402 source.n53 source.n52 9.3005
R403 source.n51 source.n50 9.3005
R404 source.n99 source.n98 9.3005
R405 source.n72 source.n71 9.3005
R406 source.n93 source.n92 9.3005
R407 source.n91 source.n90 9.3005
R408 source.n76 source.n75 9.3005
R409 source.n85 source.n84 9.3005
R410 source.n83 source.n82 9.3005
R411 source.n137 source.n136 9.3005
R412 source.n110 source.n109 9.3005
R413 source.n131 source.n130 9.3005
R414 source.n129 source.n128 9.3005
R415 source.n114 source.n113 9.3005
R416 source.n123 source.n122 9.3005
R417 source.n121 source.n120 9.3005
R418 source.n275 source.n250 8.92171
R419 source.n237 source.n212 8.92171
R420 source.n205 source.n180 8.92171
R421 source.n167 source.n142 8.92171
R422 source.n27 source.n2 8.92171
R423 source.n65 source.n40 8.92171
R424 source.n97 source.n72 8.92171
R425 source.n135 source.n110 8.92171
R426 source.n276 source.n248 8.14595
R427 source.n238 source.n210 8.14595
R428 source.n206 source.n178 8.14595
R429 source.n168 source.n140 8.14595
R430 source.n28 source.n0 8.14595
R431 source.n66 source.n38 8.14595
R432 source.n98 source.n70 8.14595
R433 source.n136 source.n108 8.14595
R434 source.n280 source.n279 5.83671
R435 source.n278 source.n248 5.81868
R436 source.n240 source.n210 5.81868
R437 source.n208 source.n178 5.81868
R438 source.n170 source.n140 5.81868
R439 source.n30 source.n0 5.81868
R440 source.n68 source.n38 5.81868
R441 source.n100 source.n70 5.81868
R442 source.n138 source.n108 5.81868
R443 source.n276 source.n275 5.04292
R444 source.n238 source.n237 5.04292
R445 source.n206 source.n205 5.04292
R446 source.n168 source.n167 5.04292
R447 source.n28 source.n27 5.04292
R448 source.n66 source.n65 5.04292
R449 source.n98 source.n97 5.04292
R450 source.n136 source.n135 5.04292
R451 source.n261 source.n257 4.38594
R452 source.n223 source.n219 4.38594
R453 source.n191 source.n187 4.38594
R454 source.n153 source.n149 4.38594
R455 source.n13 source.n9 4.38594
R456 source.n51 source.n47 4.38594
R457 source.n83 source.n79 4.38594
R458 source.n121 source.n117 4.38594
R459 source.n272 source.n250 4.26717
R460 source.n234 source.n212 4.26717
R461 source.n202 source.n180 4.26717
R462 source.n164 source.n142 4.26717
R463 source.n24 source.n2 4.26717
R464 source.n62 source.n40 4.26717
R465 source.n94 source.n72 4.26717
R466 source.n132 source.n110 4.26717
R467 source.n271 source.n252 3.49141
R468 source.n233 source.n214 3.49141
R469 source.n201 source.n182 3.49141
R470 source.n163 source.n144 3.49141
R471 source.n23 source.n4 3.49141
R472 source.n61 source.n42 3.49141
R473 source.n93 source.n74 3.49141
R474 source.n131 source.n112 3.49141
R475 source.n246 source.t12 3.3005
R476 source.n246 source.t9 3.3005
R477 source.n244 source.t8 3.3005
R478 source.n244 source.t4 3.3005
R479 source.n242 source.t6 3.3005
R480 source.n242 source.t10 3.3005
R481 source.n176 source.t15 3.3005
R482 source.n176 source.t18 3.3005
R483 source.n174 source.t26 3.3005
R484 source.n174 source.t19 3.3005
R485 source.n172 source.t21 3.3005
R486 source.n172 source.t17 3.3005
R487 source.n32 source.t24 3.3005
R488 source.n32 source.t20 3.3005
R489 source.n34 source.t25 3.3005
R490 source.n34 source.t22 3.3005
R491 source.n36 source.t27 3.3005
R492 source.n36 source.t28 3.3005
R493 source.n102 source.t5 3.3005
R494 source.n102 source.t29 3.3005
R495 source.n104 source.t3 3.3005
R496 source.n104 source.t2 3.3005
R497 source.n106 source.t7 3.3005
R498 source.n106 source.t0 3.3005
R499 source.n268 source.n267 2.71565
R500 source.n230 source.n229 2.71565
R501 source.n198 source.n197 2.71565
R502 source.n160 source.n159 2.71565
R503 source.n20 source.n19 2.71565
R504 source.n58 source.n57 2.71565
R505 source.n90 source.n89 2.71565
R506 source.n128 source.n127 2.71565
R507 source.n264 source.n254 1.93989
R508 source.n226 source.n216 1.93989
R509 source.n194 source.n184 1.93989
R510 source.n156 source.n146 1.93989
R511 source.n16 source.n6 1.93989
R512 source.n54 source.n44 1.93989
R513 source.n86 source.n76 1.93989
R514 source.n124 source.n114 1.93989
R515 source.n263 source.n256 1.16414
R516 source.n225 source.n218 1.16414
R517 source.n193 source.n186 1.16414
R518 source.n155 source.n148 1.16414
R519 source.n15 source.n8 1.16414
R520 source.n53 source.n46 1.16414
R521 source.n85 source.n78 1.16414
R522 source.n123 source.n116 1.16414
R523 source.n139 source.n107 1.14705
R524 source.n107 source.n105 1.14705
R525 source.n105 source.n103 1.14705
R526 source.n103 source.n101 1.14705
R527 source.n69 source.n37 1.14705
R528 source.n37 source.n35 1.14705
R529 source.n35 source.n33 1.14705
R530 source.n33 source.n31 1.14705
R531 source.n173 source.n171 1.14705
R532 source.n175 source.n173 1.14705
R533 source.n177 source.n175 1.14705
R534 source.n209 source.n177 1.14705
R535 source.n243 source.n241 1.14705
R536 source.n245 source.n243 1.14705
R537 source.n247 source.n245 1.14705
R538 source.n279 source.n247 1.14705
R539 source.n101 source.n69 0.470328
R540 source.n241 source.n209 0.470328
R541 source.n260 source.n259 0.388379
R542 source.n222 source.n221 0.388379
R543 source.n190 source.n189 0.388379
R544 source.n152 source.n151 0.388379
R545 source.n12 source.n11 0.388379
R546 source.n50 source.n49 0.388379
R547 source.n82 source.n81 0.388379
R548 source.n120 source.n119 0.388379
R549 source source.n280 0.188
R550 source.n262 source.n261 0.155672
R551 source.n262 source.n253 0.155672
R552 source.n269 source.n253 0.155672
R553 source.n270 source.n269 0.155672
R554 source.n270 source.n249 0.155672
R555 source.n277 source.n249 0.155672
R556 source.n224 source.n223 0.155672
R557 source.n224 source.n215 0.155672
R558 source.n231 source.n215 0.155672
R559 source.n232 source.n231 0.155672
R560 source.n232 source.n211 0.155672
R561 source.n239 source.n211 0.155672
R562 source.n192 source.n191 0.155672
R563 source.n192 source.n183 0.155672
R564 source.n199 source.n183 0.155672
R565 source.n200 source.n199 0.155672
R566 source.n200 source.n179 0.155672
R567 source.n207 source.n179 0.155672
R568 source.n154 source.n153 0.155672
R569 source.n154 source.n145 0.155672
R570 source.n161 source.n145 0.155672
R571 source.n162 source.n161 0.155672
R572 source.n162 source.n141 0.155672
R573 source.n169 source.n141 0.155672
R574 source.n29 source.n1 0.155672
R575 source.n22 source.n1 0.155672
R576 source.n22 source.n21 0.155672
R577 source.n21 source.n5 0.155672
R578 source.n14 source.n5 0.155672
R579 source.n14 source.n13 0.155672
R580 source.n67 source.n39 0.155672
R581 source.n60 source.n39 0.155672
R582 source.n60 source.n59 0.155672
R583 source.n59 source.n43 0.155672
R584 source.n52 source.n43 0.155672
R585 source.n52 source.n51 0.155672
R586 source.n99 source.n71 0.155672
R587 source.n92 source.n71 0.155672
R588 source.n92 source.n91 0.155672
R589 source.n91 source.n75 0.155672
R590 source.n84 source.n75 0.155672
R591 source.n84 source.n83 0.155672
R592 source.n137 source.n109 0.155672
R593 source.n130 source.n109 0.155672
R594 source.n130 source.n129 0.155672
R595 source.n129 source.n113 0.155672
R596 source.n122 source.n113 0.155672
R597 source.n122 source.n121 0.155672
R598 minus.n10 minus.t8 198.156
R599 minus.n48 minus.t9 198.156
R600 minus.n37 minus.t3 183.883
R601 minus.n76 minus.t1 183.883
R602 minus.n36 minus.n0 161.3
R603 minus.n34 minus.n33 161.3
R604 minus.n32 minus.n1 161.3
R605 minus.n31 minus.n30 161.3
R606 minus.n28 minus.n2 161.3
R607 minus.n27 minus.n26 161.3
R608 minus.n25 minus.n3 161.3
R609 minus.n24 minus.n23 161.3
R610 minus.n22 minus.n4 161.3
R611 minus.n20 minus.n19 161.3
R612 minus.n18 minus.n6 161.3
R613 minus.n17 minus.n16 161.3
R614 minus.n14 minus.n7 161.3
R615 minus.n13 minus.n12 161.3
R616 minus.n11 minus.n8 161.3
R617 minus.n75 minus.n39 161.3
R618 minus.n73 minus.n72 161.3
R619 minus.n71 minus.n40 161.3
R620 minus.n70 minus.n69 161.3
R621 minus.n67 minus.n41 161.3
R622 minus.n66 minus.n65 161.3
R623 minus.n64 minus.n42 161.3
R624 minus.n63 minus.n62 161.3
R625 minus.n60 minus.n43 161.3
R626 minus.n58 minus.n57 161.3
R627 minus.n56 minus.n44 161.3
R628 minus.n55 minus.n54 161.3
R629 minus.n52 minus.n45 161.3
R630 minus.n51 minus.n50 161.3
R631 minus.n49 minus.n46 161.3
R632 minus.n9 minus.t13 144.601
R633 minus.n15 minus.t11 144.601
R634 minus.n21 minus.t15 144.601
R635 minus.n5 minus.t2 144.601
R636 minus.n29 minus.t0 144.601
R637 minus.n35 minus.t4 144.601
R638 minus.n47 minus.t6 144.601
R639 minus.n53 minus.t14 144.601
R640 minus.n59 minus.t12 144.601
R641 minus.n61 minus.t5 144.601
R642 minus.n68 minus.t10 144.601
R643 minus.n74 minus.t7 144.601
R644 minus.n38 minus.n37 80.6037
R645 minus.n77 minus.n76 80.6037
R646 minus.n23 minus.n22 56.5617
R647 minus.n62 minus.n60 56.5617
R648 minus.n37 minus.n36 51.8893
R649 minus.n76 minus.n75 51.8893
R650 minus.n10 minus.n9 49.3649
R651 minus.n48 minus.n47 49.3649
R652 minus.n14 minus.n13 49.296
R653 minus.n30 minus.n1 49.296
R654 minus.n52 minus.n51 49.296
R655 minus.n69 minus.n40 49.296
R656 minus.n16 minus.n6 48.3272
R657 minus.n28 minus.n27 48.3272
R658 minus.n54 minus.n44 48.3272
R659 minus.n67 minus.n66 48.3272
R660 minus.n11 minus.n10 44.557
R661 minus.n49 minus.n48 44.557
R662 minus.n78 minus.n38 36.7017
R663 minus.n20 minus.n6 32.8269
R664 minus.n27 minus.n3 32.8269
R665 minus.n58 minus.n44 32.8269
R666 minus.n66 minus.n42 32.8269
R667 minus.n13 minus.n8 31.8581
R668 minus.n34 minus.n1 31.8581
R669 minus.n51 minus.n46 31.8581
R670 minus.n73 minus.n40 31.8581
R671 minus.n36 minus.n35 20.9036
R672 minus.n75 minus.n74 20.9036
R673 minus.n22 minus.n21 20.4117
R674 minus.n23 minus.n5 20.4117
R675 minus.n60 minus.n59 20.4117
R676 minus.n62 minus.n61 20.4117
R677 minus.n15 minus.n14 12.5423
R678 minus.n30 minus.n29 12.5423
R679 minus.n53 minus.n52 12.5423
R680 minus.n69 minus.n68 12.5423
R681 minus.n16 minus.n15 12.0505
R682 minus.n29 minus.n28 12.0505
R683 minus.n54 minus.n53 12.0505
R684 minus.n68 minus.n67 12.0505
R685 minus.n78 minus.n77 6.84564
R686 minus.n21 minus.n20 4.18111
R687 minus.n5 minus.n3 4.18111
R688 minus.n59 minus.n58 4.18111
R689 minus.n61 minus.n42 4.18111
R690 minus.n9 minus.n8 3.68928
R691 minus.n35 minus.n34 3.68928
R692 minus.n47 minus.n46 3.68928
R693 minus.n74 minus.n73 3.68928
R694 minus.n38 minus.n0 0.285035
R695 minus.n77 minus.n39 0.285035
R696 minus.n33 minus.n0 0.189894
R697 minus.n33 minus.n32 0.189894
R698 minus.n32 minus.n31 0.189894
R699 minus.n31 minus.n2 0.189894
R700 minus.n26 minus.n2 0.189894
R701 minus.n26 minus.n25 0.189894
R702 minus.n25 minus.n24 0.189894
R703 minus.n24 minus.n4 0.189894
R704 minus.n19 minus.n4 0.189894
R705 minus.n19 minus.n18 0.189894
R706 minus.n18 minus.n17 0.189894
R707 minus.n17 minus.n7 0.189894
R708 minus.n12 minus.n7 0.189894
R709 minus.n12 minus.n11 0.189894
R710 minus.n50 minus.n49 0.189894
R711 minus.n50 minus.n45 0.189894
R712 minus.n55 minus.n45 0.189894
R713 minus.n56 minus.n55 0.189894
R714 minus.n57 minus.n56 0.189894
R715 minus.n57 minus.n43 0.189894
R716 minus.n63 minus.n43 0.189894
R717 minus.n64 minus.n63 0.189894
R718 minus.n65 minus.n64 0.189894
R719 minus.n65 minus.n41 0.189894
R720 minus.n70 minus.n41 0.189894
R721 minus.n71 minus.n70 0.189894
R722 minus.n72 minus.n71 0.189894
R723 minus.n72 minus.n39 0.189894
R724 minus minus.n78 0.188
R725 drain_right.n5 drain_right.n3 68.3372
R726 drain_right.n2 drain_right.n0 68.3372
R727 drain_right.n9 drain_right.n7 68.3372
R728 drain_right.n9 drain_right.n8 67.1908
R729 drain_right.n11 drain_right.n10 67.1908
R730 drain_right.n13 drain_right.n12 67.1908
R731 drain_right.n5 drain_right.n4 67.1907
R732 drain_right.n2 drain_right.n1 67.1907
R733 drain_right drain_right.n6 29.721
R734 drain_right drain_right.n13 6.79977
R735 drain_right.n3 drain_right.t8 3.3005
R736 drain_right.n3 drain_right.t14 3.3005
R737 drain_right.n4 drain_right.t10 3.3005
R738 drain_right.n4 drain_right.t5 3.3005
R739 drain_right.n1 drain_right.t1 3.3005
R740 drain_right.n1 drain_right.t3 3.3005
R741 drain_right.n0 drain_right.t6 3.3005
R742 drain_right.n0 drain_right.t9 3.3005
R743 drain_right.n7 drain_right.t2 3.3005
R744 drain_right.n7 drain_right.t7 3.3005
R745 drain_right.n8 drain_right.t0 3.3005
R746 drain_right.n8 drain_right.t4 3.3005
R747 drain_right.n10 drain_right.t15 3.3005
R748 drain_right.n10 drain_right.t13 3.3005
R749 drain_right.n12 drain_right.t12 3.3005
R750 drain_right.n12 drain_right.t11 3.3005
R751 drain_right.n13 drain_right.n11 1.14705
R752 drain_right.n11 drain_right.n9 1.14705
R753 drain_right.n6 drain_right.n5 0.51843
R754 drain_right.n6 drain_right.n2 0.51843
C0 source minus 7.03926f
C1 drain_left minus 0.174261f
C2 source drain_right 10.3801f
C3 plus minus 5.90846f
C4 drain_left drain_right 1.64323f
C5 plus drain_right 0.468824f
C6 drain_right minus 6.42775f
C7 source drain_left 10.3762f
C8 source plus 7.05328f
C9 plus drain_left 6.7386f
C10 drain_right a_n3110_n2088# 6.16579f
C11 drain_left a_n3110_n2088# 6.60225f
C12 source a_n3110_n2088# 5.921499f
C13 minus a_n3110_n2088# 11.975189f
C14 plus a_n3110_n2088# 13.37842f
C15 drain_right.t6 a_n3110_n2088# 0.121258f
C16 drain_right.t9 a_n3110_n2088# 0.121258f
C17 drain_right.n0 a_n3110_n2088# 1.01812f
C18 drain_right.t1 a_n3110_n2088# 0.121258f
C19 drain_right.t3 a_n3110_n2088# 0.121258f
C20 drain_right.n1 a_n3110_n2088# 1.01129f
C21 drain_right.n2 a_n3110_n2088# 0.74589f
C22 drain_right.t8 a_n3110_n2088# 0.121258f
C23 drain_right.t14 a_n3110_n2088# 0.121258f
C24 drain_right.n3 a_n3110_n2088# 1.01812f
C25 drain_right.t10 a_n3110_n2088# 0.121258f
C26 drain_right.t5 a_n3110_n2088# 0.121258f
C27 drain_right.n4 a_n3110_n2088# 1.01129f
C28 drain_right.n5 a_n3110_n2088# 0.74589f
C29 drain_right.n6 a_n3110_n2088# 1.23911f
C30 drain_right.t2 a_n3110_n2088# 0.121258f
C31 drain_right.t7 a_n3110_n2088# 0.121258f
C32 drain_right.n7 a_n3110_n2088# 1.01812f
C33 drain_right.t0 a_n3110_n2088# 0.121258f
C34 drain_right.t4 a_n3110_n2088# 0.121258f
C35 drain_right.n8 a_n3110_n2088# 1.01129f
C36 drain_right.n9 a_n3110_n2088# 0.796543f
C37 drain_right.t15 a_n3110_n2088# 0.121258f
C38 drain_right.t13 a_n3110_n2088# 0.121258f
C39 drain_right.n10 a_n3110_n2088# 1.01129f
C40 drain_right.n11 a_n3110_n2088# 0.396532f
C41 drain_right.t12 a_n3110_n2088# 0.121258f
C42 drain_right.t11 a_n3110_n2088# 0.121258f
C43 drain_right.n12 a_n3110_n2088# 1.01129f
C44 drain_right.n13 a_n3110_n2088# 0.631852f
C45 minus.n0 a_n3110_n2088# 0.048137f
C46 minus.t4 a_n3110_n2088# 0.57289f
C47 minus.n1 a_n3110_n2088# 0.033042f
C48 minus.n2 a_n3110_n2088# 0.036075f
C49 minus.t0 a_n3110_n2088# 0.57289f
C50 minus.n3 a_n3110_n2088# 0.044954f
C51 minus.n4 a_n3110_n2088# 0.036075f
C52 minus.t2 a_n3110_n2088# 0.57289f
C53 minus.n5 a_n3110_n2088# 0.235222f
C54 minus.t15 a_n3110_n2088# 0.57289f
C55 minus.n6 a_n3110_n2088# 0.032191f
C56 minus.n7 a_n3110_n2088# 0.036075f
C57 minus.t11 a_n3110_n2088# 0.57289f
C58 minus.n8 a_n3110_n2088# 0.044098f
C59 minus.t8 a_n3110_n2088# 0.648673f
C60 minus.t13 a_n3110_n2088# 0.57289f
C61 minus.n9 a_n3110_n2088# 0.261335f
C62 minus.n10 a_n3110_n2088# 0.288324f
C63 minus.n11 a_n3110_n2088# 0.15047f
C64 minus.n12 a_n3110_n2088# 0.036075f
C65 minus.n13 a_n3110_n2088# 0.033042f
C66 minus.n14 a_n3110_n2088# 0.050384f
C67 minus.n15 a_n3110_n2088# 0.235222f
C68 minus.n16 a_n3110_n2088# 0.050379f
C69 minus.n17 a_n3110_n2088# 0.036075f
C70 minus.n18 a_n3110_n2088# 0.036075f
C71 minus.n19 a_n3110_n2088# 0.036075f
C72 minus.n20 a_n3110_n2088# 0.044954f
C73 minus.n21 a_n3110_n2088# 0.235222f
C74 minus.n22 a_n3110_n2088# 0.046826f
C75 minus.n23 a_n3110_n2088# 0.046826f
C76 minus.n24 a_n3110_n2088# 0.036075f
C77 minus.n25 a_n3110_n2088# 0.036075f
C78 minus.n26 a_n3110_n2088# 0.036075f
C79 minus.n27 a_n3110_n2088# 0.032191f
C80 minus.n28 a_n3110_n2088# 0.050379f
C81 minus.n29 a_n3110_n2088# 0.235222f
C82 minus.n30 a_n3110_n2088# 0.050384f
C83 minus.n31 a_n3110_n2088# 0.036075f
C84 minus.n32 a_n3110_n2088# 0.036075f
C85 minus.n33 a_n3110_n2088# 0.036075f
C86 minus.n34 a_n3110_n2088# 0.044098f
C87 minus.n35 a_n3110_n2088# 0.235222f
C88 minus.n36 a_n3110_n2088# 0.045291f
C89 minus.t3 a_n3110_n2088# 0.62782f
C90 minus.n37 a_n3110_n2088# 0.289274f
C91 minus.n38 a_n3110_n2088# 1.32519f
C92 minus.n39 a_n3110_n2088# 0.048137f
C93 minus.t7 a_n3110_n2088# 0.57289f
C94 minus.n40 a_n3110_n2088# 0.033042f
C95 minus.n41 a_n3110_n2088# 0.036075f
C96 minus.t10 a_n3110_n2088# 0.57289f
C97 minus.n42 a_n3110_n2088# 0.044954f
C98 minus.n43 a_n3110_n2088# 0.036075f
C99 minus.t12 a_n3110_n2088# 0.57289f
C100 minus.n44 a_n3110_n2088# 0.032191f
C101 minus.n45 a_n3110_n2088# 0.036075f
C102 minus.t14 a_n3110_n2088# 0.57289f
C103 minus.n46 a_n3110_n2088# 0.044098f
C104 minus.t9 a_n3110_n2088# 0.648673f
C105 minus.t6 a_n3110_n2088# 0.57289f
C106 minus.n47 a_n3110_n2088# 0.261335f
C107 minus.n48 a_n3110_n2088# 0.288324f
C108 minus.n49 a_n3110_n2088# 0.15047f
C109 minus.n50 a_n3110_n2088# 0.036075f
C110 minus.n51 a_n3110_n2088# 0.033042f
C111 minus.n52 a_n3110_n2088# 0.050384f
C112 minus.n53 a_n3110_n2088# 0.235222f
C113 minus.n54 a_n3110_n2088# 0.050379f
C114 minus.n55 a_n3110_n2088# 0.036075f
C115 minus.n56 a_n3110_n2088# 0.036075f
C116 minus.n57 a_n3110_n2088# 0.036075f
C117 minus.n58 a_n3110_n2088# 0.044954f
C118 minus.n59 a_n3110_n2088# 0.235222f
C119 minus.n60 a_n3110_n2088# 0.046826f
C120 minus.t5 a_n3110_n2088# 0.57289f
C121 minus.n61 a_n3110_n2088# 0.235222f
C122 minus.n62 a_n3110_n2088# 0.046826f
C123 minus.n63 a_n3110_n2088# 0.036075f
C124 minus.n64 a_n3110_n2088# 0.036075f
C125 minus.n65 a_n3110_n2088# 0.036075f
C126 minus.n66 a_n3110_n2088# 0.032191f
C127 minus.n67 a_n3110_n2088# 0.050379f
C128 minus.n68 a_n3110_n2088# 0.235222f
C129 minus.n69 a_n3110_n2088# 0.050384f
C130 minus.n70 a_n3110_n2088# 0.036075f
C131 minus.n71 a_n3110_n2088# 0.036075f
C132 minus.n72 a_n3110_n2088# 0.036075f
C133 minus.n73 a_n3110_n2088# 0.044098f
C134 minus.n74 a_n3110_n2088# 0.235222f
C135 minus.n75 a_n3110_n2088# 0.045291f
C136 minus.t1 a_n3110_n2088# 0.62782f
C137 minus.n76 a_n3110_n2088# 0.289274f
C138 minus.n77 a_n3110_n2088# 0.277334f
C139 minus.n78 a_n3110_n2088# 1.58282f
C140 source.n0 a_n3110_n2088# 0.034652f
C141 source.n1 a_n3110_n2088# 0.024653f
C142 source.n2 a_n3110_n2088# 0.013247f
C143 source.n3 a_n3110_n2088# 0.031312f
C144 source.n4 a_n3110_n2088# 0.014027f
C145 source.n5 a_n3110_n2088# 0.024653f
C146 source.n6 a_n3110_n2088# 0.013247f
C147 source.n7 a_n3110_n2088# 0.031312f
C148 source.n8 a_n3110_n2088# 0.014027f
C149 source.n9 a_n3110_n2088# 0.105496f
C150 source.t23 a_n3110_n2088# 0.051034f
C151 source.n10 a_n3110_n2088# 0.023484f
C152 source.n11 a_n3110_n2088# 0.018496f
C153 source.n12 a_n3110_n2088# 0.013247f
C154 source.n13 a_n3110_n2088# 0.586587f
C155 source.n14 a_n3110_n2088# 0.024653f
C156 source.n15 a_n3110_n2088# 0.013247f
C157 source.n16 a_n3110_n2088# 0.014027f
C158 source.n17 a_n3110_n2088# 0.031312f
C159 source.n18 a_n3110_n2088# 0.031312f
C160 source.n19 a_n3110_n2088# 0.014027f
C161 source.n20 a_n3110_n2088# 0.013247f
C162 source.n21 a_n3110_n2088# 0.024653f
C163 source.n22 a_n3110_n2088# 0.024653f
C164 source.n23 a_n3110_n2088# 0.013247f
C165 source.n24 a_n3110_n2088# 0.014027f
C166 source.n25 a_n3110_n2088# 0.031312f
C167 source.n26 a_n3110_n2088# 0.067785f
C168 source.n27 a_n3110_n2088# 0.014027f
C169 source.n28 a_n3110_n2088# 0.013247f
C170 source.n29 a_n3110_n2088# 0.056984f
C171 source.n30 a_n3110_n2088# 0.037928f
C172 source.n31 a_n3110_n2088# 0.679068f
C173 source.t24 a_n3110_n2088# 0.116888f
C174 source.t20 a_n3110_n2088# 0.116888f
C175 source.n32 a_n3110_n2088# 0.910333f
C176 source.n33 a_n3110_n2088# 0.413252f
C177 source.t25 a_n3110_n2088# 0.116888f
C178 source.t22 a_n3110_n2088# 0.116888f
C179 source.n34 a_n3110_n2088# 0.910333f
C180 source.n35 a_n3110_n2088# 0.413252f
C181 source.t27 a_n3110_n2088# 0.116888f
C182 source.t28 a_n3110_n2088# 0.116888f
C183 source.n36 a_n3110_n2088# 0.910333f
C184 source.n37 a_n3110_n2088# 0.413252f
C185 source.n38 a_n3110_n2088# 0.034652f
C186 source.n39 a_n3110_n2088# 0.024653f
C187 source.n40 a_n3110_n2088# 0.013247f
C188 source.n41 a_n3110_n2088# 0.031312f
C189 source.n42 a_n3110_n2088# 0.014027f
C190 source.n43 a_n3110_n2088# 0.024653f
C191 source.n44 a_n3110_n2088# 0.013247f
C192 source.n45 a_n3110_n2088# 0.031312f
C193 source.n46 a_n3110_n2088# 0.014027f
C194 source.n47 a_n3110_n2088# 0.105496f
C195 source.t13 a_n3110_n2088# 0.051034f
C196 source.n48 a_n3110_n2088# 0.023484f
C197 source.n49 a_n3110_n2088# 0.018496f
C198 source.n50 a_n3110_n2088# 0.013247f
C199 source.n51 a_n3110_n2088# 0.586587f
C200 source.n52 a_n3110_n2088# 0.024653f
C201 source.n53 a_n3110_n2088# 0.013247f
C202 source.n54 a_n3110_n2088# 0.014027f
C203 source.n55 a_n3110_n2088# 0.031312f
C204 source.n56 a_n3110_n2088# 0.031312f
C205 source.n57 a_n3110_n2088# 0.014027f
C206 source.n58 a_n3110_n2088# 0.013247f
C207 source.n59 a_n3110_n2088# 0.024653f
C208 source.n60 a_n3110_n2088# 0.024653f
C209 source.n61 a_n3110_n2088# 0.013247f
C210 source.n62 a_n3110_n2088# 0.014027f
C211 source.n63 a_n3110_n2088# 0.031312f
C212 source.n64 a_n3110_n2088# 0.067785f
C213 source.n65 a_n3110_n2088# 0.014027f
C214 source.n66 a_n3110_n2088# 0.013247f
C215 source.n67 a_n3110_n2088# 0.056984f
C216 source.n68 a_n3110_n2088# 0.037928f
C217 source.n69 a_n3110_n2088# 0.149455f
C218 source.n70 a_n3110_n2088# 0.034652f
C219 source.n71 a_n3110_n2088# 0.024653f
C220 source.n72 a_n3110_n2088# 0.013247f
C221 source.n73 a_n3110_n2088# 0.031312f
C222 source.n74 a_n3110_n2088# 0.014027f
C223 source.n75 a_n3110_n2088# 0.024653f
C224 source.n76 a_n3110_n2088# 0.013247f
C225 source.n77 a_n3110_n2088# 0.031312f
C226 source.n78 a_n3110_n2088# 0.014027f
C227 source.n79 a_n3110_n2088# 0.105496f
C228 source.t31 a_n3110_n2088# 0.051034f
C229 source.n80 a_n3110_n2088# 0.023484f
C230 source.n81 a_n3110_n2088# 0.018496f
C231 source.n82 a_n3110_n2088# 0.013247f
C232 source.n83 a_n3110_n2088# 0.586587f
C233 source.n84 a_n3110_n2088# 0.024653f
C234 source.n85 a_n3110_n2088# 0.013247f
C235 source.n86 a_n3110_n2088# 0.014027f
C236 source.n87 a_n3110_n2088# 0.031312f
C237 source.n88 a_n3110_n2088# 0.031312f
C238 source.n89 a_n3110_n2088# 0.014027f
C239 source.n90 a_n3110_n2088# 0.013247f
C240 source.n91 a_n3110_n2088# 0.024653f
C241 source.n92 a_n3110_n2088# 0.024653f
C242 source.n93 a_n3110_n2088# 0.013247f
C243 source.n94 a_n3110_n2088# 0.014027f
C244 source.n95 a_n3110_n2088# 0.031312f
C245 source.n96 a_n3110_n2088# 0.067785f
C246 source.n97 a_n3110_n2088# 0.014027f
C247 source.n98 a_n3110_n2088# 0.013247f
C248 source.n99 a_n3110_n2088# 0.056984f
C249 source.n100 a_n3110_n2088# 0.037928f
C250 source.n101 a_n3110_n2088# 0.149455f
C251 source.t5 a_n3110_n2088# 0.116888f
C252 source.t29 a_n3110_n2088# 0.116888f
C253 source.n102 a_n3110_n2088# 0.910333f
C254 source.n103 a_n3110_n2088# 0.413252f
C255 source.t3 a_n3110_n2088# 0.116888f
C256 source.t2 a_n3110_n2088# 0.116888f
C257 source.n104 a_n3110_n2088# 0.910333f
C258 source.n105 a_n3110_n2088# 0.413252f
C259 source.t7 a_n3110_n2088# 0.116888f
C260 source.t0 a_n3110_n2088# 0.116888f
C261 source.n106 a_n3110_n2088# 0.910333f
C262 source.n107 a_n3110_n2088# 0.413252f
C263 source.n108 a_n3110_n2088# 0.034652f
C264 source.n109 a_n3110_n2088# 0.024653f
C265 source.n110 a_n3110_n2088# 0.013247f
C266 source.n111 a_n3110_n2088# 0.031312f
C267 source.n112 a_n3110_n2088# 0.014027f
C268 source.n113 a_n3110_n2088# 0.024653f
C269 source.n114 a_n3110_n2088# 0.013247f
C270 source.n115 a_n3110_n2088# 0.031312f
C271 source.n116 a_n3110_n2088# 0.014027f
C272 source.n117 a_n3110_n2088# 0.105496f
C273 source.t1 a_n3110_n2088# 0.051034f
C274 source.n118 a_n3110_n2088# 0.023484f
C275 source.n119 a_n3110_n2088# 0.018496f
C276 source.n120 a_n3110_n2088# 0.013247f
C277 source.n121 a_n3110_n2088# 0.586587f
C278 source.n122 a_n3110_n2088# 0.024653f
C279 source.n123 a_n3110_n2088# 0.013247f
C280 source.n124 a_n3110_n2088# 0.014027f
C281 source.n125 a_n3110_n2088# 0.031312f
C282 source.n126 a_n3110_n2088# 0.031312f
C283 source.n127 a_n3110_n2088# 0.014027f
C284 source.n128 a_n3110_n2088# 0.013247f
C285 source.n129 a_n3110_n2088# 0.024653f
C286 source.n130 a_n3110_n2088# 0.024653f
C287 source.n131 a_n3110_n2088# 0.013247f
C288 source.n132 a_n3110_n2088# 0.014027f
C289 source.n133 a_n3110_n2088# 0.031312f
C290 source.n134 a_n3110_n2088# 0.067785f
C291 source.n135 a_n3110_n2088# 0.014027f
C292 source.n136 a_n3110_n2088# 0.013247f
C293 source.n137 a_n3110_n2088# 0.056984f
C294 source.n138 a_n3110_n2088# 0.037928f
C295 source.n139 a_n3110_n2088# 1.01039f
C296 source.n140 a_n3110_n2088# 0.034652f
C297 source.n141 a_n3110_n2088# 0.024653f
C298 source.n142 a_n3110_n2088# 0.013247f
C299 source.n143 a_n3110_n2088# 0.031312f
C300 source.n144 a_n3110_n2088# 0.014027f
C301 source.n145 a_n3110_n2088# 0.024653f
C302 source.n146 a_n3110_n2088# 0.013247f
C303 source.n147 a_n3110_n2088# 0.031312f
C304 source.n148 a_n3110_n2088# 0.014027f
C305 source.n149 a_n3110_n2088# 0.105496f
C306 source.t14 a_n3110_n2088# 0.051034f
C307 source.n150 a_n3110_n2088# 0.023484f
C308 source.n151 a_n3110_n2088# 0.018496f
C309 source.n152 a_n3110_n2088# 0.013247f
C310 source.n153 a_n3110_n2088# 0.586587f
C311 source.n154 a_n3110_n2088# 0.024653f
C312 source.n155 a_n3110_n2088# 0.013247f
C313 source.n156 a_n3110_n2088# 0.014027f
C314 source.n157 a_n3110_n2088# 0.031312f
C315 source.n158 a_n3110_n2088# 0.031312f
C316 source.n159 a_n3110_n2088# 0.014027f
C317 source.n160 a_n3110_n2088# 0.013247f
C318 source.n161 a_n3110_n2088# 0.024653f
C319 source.n162 a_n3110_n2088# 0.024653f
C320 source.n163 a_n3110_n2088# 0.013247f
C321 source.n164 a_n3110_n2088# 0.014027f
C322 source.n165 a_n3110_n2088# 0.031312f
C323 source.n166 a_n3110_n2088# 0.067785f
C324 source.n167 a_n3110_n2088# 0.014027f
C325 source.n168 a_n3110_n2088# 0.013247f
C326 source.n169 a_n3110_n2088# 0.056984f
C327 source.n170 a_n3110_n2088# 0.037928f
C328 source.n171 a_n3110_n2088# 1.01039f
C329 source.t21 a_n3110_n2088# 0.116888f
C330 source.t17 a_n3110_n2088# 0.116888f
C331 source.n172 a_n3110_n2088# 0.910327f
C332 source.n173 a_n3110_n2088# 0.413258f
C333 source.t26 a_n3110_n2088# 0.116888f
C334 source.t19 a_n3110_n2088# 0.116888f
C335 source.n174 a_n3110_n2088# 0.910327f
C336 source.n175 a_n3110_n2088# 0.413258f
C337 source.t15 a_n3110_n2088# 0.116888f
C338 source.t18 a_n3110_n2088# 0.116888f
C339 source.n176 a_n3110_n2088# 0.910327f
C340 source.n177 a_n3110_n2088# 0.413258f
C341 source.n178 a_n3110_n2088# 0.034652f
C342 source.n179 a_n3110_n2088# 0.024653f
C343 source.n180 a_n3110_n2088# 0.013247f
C344 source.n181 a_n3110_n2088# 0.031312f
C345 source.n182 a_n3110_n2088# 0.014027f
C346 source.n183 a_n3110_n2088# 0.024653f
C347 source.n184 a_n3110_n2088# 0.013247f
C348 source.n185 a_n3110_n2088# 0.031312f
C349 source.n186 a_n3110_n2088# 0.014027f
C350 source.n187 a_n3110_n2088# 0.105496f
C351 source.t16 a_n3110_n2088# 0.051034f
C352 source.n188 a_n3110_n2088# 0.023484f
C353 source.n189 a_n3110_n2088# 0.018496f
C354 source.n190 a_n3110_n2088# 0.013247f
C355 source.n191 a_n3110_n2088# 0.586587f
C356 source.n192 a_n3110_n2088# 0.024653f
C357 source.n193 a_n3110_n2088# 0.013247f
C358 source.n194 a_n3110_n2088# 0.014027f
C359 source.n195 a_n3110_n2088# 0.031312f
C360 source.n196 a_n3110_n2088# 0.031312f
C361 source.n197 a_n3110_n2088# 0.014027f
C362 source.n198 a_n3110_n2088# 0.013247f
C363 source.n199 a_n3110_n2088# 0.024653f
C364 source.n200 a_n3110_n2088# 0.024653f
C365 source.n201 a_n3110_n2088# 0.013247f
C366 source.n202 a_n3110_n2088# 0.014027f
C367 source.n203 a_n3110_n2088# 0.031312f
C368 source.n204 a_n3110_n2088# 0.067785f
C369 source.n205 a_n3110_n2088# 0.014027f
C370 source.n206 a_n3110_n2088# 0.013247f
C371 source.n207 a_n3110_n2088# 0.056984f
C372 source.n208 a_n3110_n2088# 0.037928f
C373 source.n209 a_n3110_n2088# 0.149455f
C374 source.n210 a_n3110_n2088# 0.034652f
C375 source.n211 a_n3110_n2088# 0.024653f
C376 source.n212 a_n3110_n2088# 0.013247f
C377 source.n213 a_n3110_n2088# 0.031312f
C378 source.n214 a_n3110_n2088# 0.014027f
C379 source.n215 a_n3110_n2088# 0.024653f
C380 source.n216 a_n3110_n2088# 0.013247f
C381 source.n217 a_n3110_n2088# 0.031312f
C382 source.n218 a_n3110_n2088# 0.014027f
C383 source.n219 a_n3110_n2088# 0.105496f
C384 source.t30 a_n3110_n2088# 0.051034f
C385 source.n220 a_n3110_n2088# 0.023484f
C386 source.n221 a_n3110_n2088# 0.018496f
C387 source.n222 a_n3110_n2088# 0.013247f
C388 source.n223 a_n3110_n2088# 0.586587f
C389 source.n224 a_n3110_n2088# 0.024653f
C390 source.n225 a_n3110_n2088# 0.013247f
C391 source.n226 a_n3110_n2088# 0.014027f
C392 source.n227 a_n3110_n2088# 0.031312f
C393 source.n228 a_n3110_n2088# 0.031312f
C394 source.n229 a_n3110_n2088# 0.014027f
C395 source.n230 a_n3110_n2088# 0.013247f
C396 source.n231 a_n3110_n2088# 0.024653f
C397 source.n232 a_n3110_n2088# 0.024653f
C398 source.n233 a_n3110_n2088# 0.013247f
C399 source.n234 a_n3110_n2088# 0.014027f
C400 source.n235 a_n3110_n2088# 0.031312f
C401 source.n236 a_n3110_n2088# 0.067785f
C402 source.n237 a_n3110_n2088# 0.014027f
C403 source.n238 a_n3110_n2088# 0.013247f
C404 source.n239 a_n3110_n2088# 0.056984f
C405 source.n240 a_n3110_n2088# 0.037928f
C406 source.n241 a_n3110_n2088# 0.149455f
C407 source.t6 a_n3110_n2088# 0.116888f
C408 source.t10 a_n3110_n2088# 0.116888f
C409 source.n242 a_n3110_n2088# 0.910327f
C410 source.n243 a_n3110_n2088# 0.413258f
C411 source.t8 a_n3110_n2088# 0.116888f
C412 source.t4 a_n3110_n2088# 0.116888f
C413 source.n244 a_n3110_n2088# 0.910327f
C414 source.n245 a_n3110_n2088# 0.413258f
C415 source.t12 a_n3110_n2088# 0.116888f
C416 source.t9 a_n3110_n2088# 0.116888f
C417 source.n246 a_n3110_n2088# 0.910327f
C418 source.n247 a_n3110_n2088# 0.413258f
C419 source.n248 a_n3110_n2088# 0.034652f
C420 source.n249 a_n3110_n2088# 0.024653f
C421 source.n250 a_n3110_n2088# 0.013247f
C422 source.n251 a_n3110_n2088# 0.031312f
C423 source.n252 a_n3110_n2088# 0.014027f
C424 source.n253 a_n3110_n2088# 0.024653f
C425 source.n254 a_n3110_n2088# 0.013247f
C426 source.n255 a_n3110_n2088# 0.031312f
C427 source.n256 a_n3110_n2088# 0.014027f
C428 source.n257 a_n3110_n2088# 0.105496f
C429 source.t11 a_n3110_n2088# 0.051034f
C430 source.n258 a_n3110_n2088# 0.023484f
C431 source.n259 a_n3110_n2088# 0.018496f
C432 source.n260 a_n3110_n2088# 0.013247f
C433 source.n261 a_n3110_n2088# 0.586587f
C434 source.n262 a_n3110_n2088# 0.024653f
C435 source.n263 a_n3110_n2088# 0.013247f
C436 source.n264 a_n3110_n2088# 0.014027f
C437 source.n265 a_n3110_n2088# 0.031312f
C438 source.n266 a_n3110_n2088# 0.031312f
C439 source.n267 a_n3110_n2088# 0.014027f
C440 source.n268 a_n3110_n2088# 0.013247f
C441 source.n269 a_n3110_n2088# 0.024653f
C442 source.n270 a_n3110_n2088# 0.024653f
C443 source.n271 a_n3110_n2088# 0.013247f
C444 source.n272 a_n3110_n2088# 0.014027f
C445 source.n273 a_n3110_n2088# 0.031312f
C446 source.n274 a_n3110_n2088# 0.067785f
C447 source.n275 a_n3110_n2088# 0.014027f
C448 source.n276 a_n3110_n2088# 0.013247f
C449 source.n277 a_n3110_n2088# 0.056984f
C450 source.n278 a_n3110_n2088# 0.037928f
C451 source.n279 a_n3110_n2088# 0.326192f
C452 source.n280 a_n3110_n2088# 1.03305f
C453 drain_left.t15 a_n3110_n2088# 0.122692f
C454 drain_left.t14 a_n3110_n2088# 0.122692f
C455 drain_left.n0 a_n3110_n2088# 1.03016f
C456 drain_left.t11 a_n3110_n2088# 0.122692f
C457 drain_left.t13 a_n3110_n2088# 0.122692f
C458 drain_left.n1 a_n3110_n2088# 1.02326f
C459 drain_left.n2 a_n3110_n2088# 0.754715f
C460 drain_left.t9 a_n3110_n2088# 0.122692f
C461 drain_left.t12 a_n3110_n2088# 0.122692f
C462 drain_left.n3 a_n3110_n2088# 1.03016f
C463 drain_left.t3 a_n3110_n2088# 0.122692f
C464 drain_left.t0 a_n3110_n2088# 0.122692f
C465 drain_left.n4 a_n3110_n2088# 1.02326f
C466 drain_left.n5 a_n3110_n2088# 0.754715f
C467 drain_left.n6 a_n3110_n2088# 1.30535f
C468 drain_left.t2 a_n3110_n2088# 0.122692f
C469 drain_left.t10 a_n3110_n2088# 0.122692f
C470 drain_left.n7 a_n3110_n2088# 1.03017f
C471 drain_left.t1 a_n3110_n2088# 0.122692f
C472 drain_left.t7 a_n3110_n2088# 0.122692f
C473 drain_left.n8 a_n3110_n2088# 1.02326f
C474 drain_left.n9 a_n3110_n2088# 0.805963f
C475 drain_left.t4 a_n3110_n2088# 0.122692f
C476 drain_left.t6 a_n3110_n2088# 0.122692f
C477 drain_left.n10 a_n3110_n2088# 1.02326f
C478 drain_left.n11 a_n3110_n2088# 0.401223f
C479 drain_left.t8 a_n3110_n2088# 0.122692f
C480 drain_left.t5 a_n3110_n2088# 0.122692f
C481 drain_left.n12 a_n3110_n2088# 1.02326f
C482 drain_left.n13 a_n3110_n2088# 0.639333f
C483 plus.n0 a_n3110_n2088# 0.049321f
C484 plus.t5 a_n3110_n2088# 0.643263f
C485 plus.t8 a_n3110_n2088# 0.586982f
C486 plus.n1 a_n3110_n2088# 0.033854f
C487 plus.n2 a_n3110_n2088# 0.036962f
C488 plus.t4 a_n3110_n2088# 0.586982f
C489 plus.n3 a_n3110_n2088# 0.04606f
C490 plus.n4 a_n3110_n2088# 0.036962f
C491 plus.t3 a_n3110_n2088# 0.586982f
C492 plus.n5 a_n3110_n2088# 0.032983f
C493 plus.n6 a_n3110_n2088# 0.036962f
C494 plus.t0 a_n3110_n2088# 0.586982f
C495 plus.n7 a_n3110_n2088# 0.045183f
C496 plus.t1 a_n3110_n2088# 0.586982f
C497 plus.n8 a_n3110_n2088# 0.267763f
C498 plus.t15 a_n3110_n2088# 0.664629f
C499 plus.n9 a_n3110_n2088# 0.295416f
C500 plus.n10 a_n3110_n2088# 0.154171f
C501 plus.n11 a_n3110_n2088# 0.036962f
C502 plus.n12 a_n3110_n2088# 0.033854f
C503 plus.n13 a_n3110_n2088# 0.051623f
C504 plus.n14 a_n3110_n2088# 0.241008f
C505 plus.n15 a_n3110_n2088# 0.051618f
C506 plus.n16 a_n3110_n2088# 0.036962f
C507 plus.n17 a_n3110_n2088# 0.036962f
C508 plus.n18 a_n3110_n2088# 0.036962f
C509 plus.n19 a_n3110_n2088# 0.04606f
C510 plus.n20 a_n3110_n2088# 0.241008f
C511 plus.n21 a_n3110_n2088# 0.047978f
C512 plus.t6 a_n3110_n2088# 0.586982f
C513 plus.n22 a_n3110_n2088# 0.241008f
C514 plus.n23 a_n3110_n2088# 0.047978f
C515 plus.n24 a_n3110_n2088# 0.036962f
C516 plus.n25 a_n3110_n2088# 0.036962f
C517 plus.n26 a_n3110_n2088# 0.036962f
C518 plus.n27 a_n3110_n2088# 0.032983f
C519 plus.n28 a_n3110_n2088# 0.051618f
C520 plus.n29 a_n3110_n2088# 0.241008f
C521 plus.n30 a_n3110_n2088# 0.051623f
C522 plus.n31 a_n3110_n2088# 0.036962f
C523 plus.n32 a_n3110_n2088# 0.036962f
C524 plus.n33 a_n3110_n2088# 0.036962f
C525 plus.n34 a_n3110_n2088# 0.045183f
C526 plus.n35 a_n3110_n2088# 0.241008f
C527 plus.n36 a_n3110_n2088# 0.046405f
C528 plus.n37 a_n3110_n2088# 0.29639f
C529 plus.n38 a_n3110_n2088# 0.360731f
C530 plus.n39 a_n3110_n2088# 0.049321f
C531 plus.t14 a_n3110_n2088# 0.643263f
C532 plus.t7 a_n3110_n2088# 0.586982f
C533 plus.n40 a_n3110_n2088# 0.033854f
C534 plus.n41 a_n3110_n2088# 0.036962f
C535 plus.t11 a_n3110_n2088# 0.586982f
C536 plus.n42 a_n3110_n2088# 0.04606f
C537 plus.n43 a_n3110_n2088# 0.036962f
C538 plus.t2 a_n3110_n2088# 0.586982f
C539 plus.n44 a_n3110_n2088# 0.241008f
C540 plus.t9 a_n3110_n2088# 0.586982f
C541 plus.n45 a_n3110_n2088# 0.032983f
C542 plus.n46 a_n3110_n2088# 0.036962f
C543 plus.t13 a_n3110_n2088# 0.586982f
C544 plus.n47 a_n3110_n2088# 0.045183f
C545 plus.t12 a_n3110_n2088# 0.664629f
C546 plus.t10 a_n3110_n2088# 0.586982f
C547 plus.n48 a_n3110_n2088# 0.267763f
C548 plus.n49 a_n3110_n2088# 0.295416f
C549 plus.n50 a_n3110_n2088# 0.154171f
C550 plus.n51 a_n3110_n2088# 0.036962f
C551 plus.n52 a_n3110_n2088# 0.033854f
C552 plus.n53 a_n3110_n2088# 0.051623f
C553 plus.n54 a_n3110_n2088# 0.241008f
C554 plus.n55 a_n3110_n2088# 0.051618f
C555 plus.n56 a_n3110_n2088# 0.036962f
C556 plus.n57 a_n3110_n2088# 0.036962f
C557 plus.n58 a_n3110_n2088# 0.036962f
C558 plus.n59 a_n3110_n2088# 0.04606f
C559 plus.n60 a_n3110_n2088# 0.241008f
C560 plus.n61 a_n3110_n2088# 0.047978f
C561 plus.n62 a_n3110_n2088# 0.047978f
C562 plus.n63 a_n3110_n2088# 0.036962f
C563 plus.n64 a_n3110_n2088# 0.036962f
C564 plus.n65 a_n3110_n2088# 0.036962f
C565 plus.n66 a_n3110_n2088# 0.032983f
C566 plus.n67 a_n3110_n2088# 0.051618f
C567 plus.n68 a_n3110_n2088# 0.241008f
C568 plus.n69 a_n3110_n2088# 0.051623f
C569 plus.n70 a_n3110_n2088# 0.036962f
C570 plus.n71 a_n3110_n2088# 0.036962f
C571 plus.n72 a_n3110_n2088# 0.036962f
C572 plus.n73 a_n3110_n2088# 0.045183f
C573 plus.n74 a_n3110_n2088# 0.241008f
C574 plus.n75 a_n3110_n2088# 0.046405f
C575 plus.n76 a_n3110_n2088# 0.29639f
C576 plus.n77 a_n3110_n2088# 1.23477f
.ends

