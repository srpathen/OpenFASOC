* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t23 minus.t0 source.t30 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X1 source.t18 plus.t0 drain_left.t23 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X2 drain_left.t22 plus.t1 source.t10 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X3 source.t28 minus.t1 drain_right.t22 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X4 a_n2406_n2088# a_n2406_n2088# a_n2406_n2088# a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X5 source.t37 minus.t2 drain_right.t21 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X6 drain_left.t21 plus.t2 source.t7 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X7 drain_left.t20 plus.t3 source.t19 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X8 drain_right.t20 minus.t3 source.t47 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X9 drain_right.t19 minus.t4 source.t39 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X10 drain_right.t18 minus.t5 source.t41 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X11 source.t23 plus.t4 drain_left.t19 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X12 a_n2406_n2088# a_n2406_n2088# a_n2406_n2088# a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X13 source.t35 minus.t6 drain_right.t17 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X14 a_n2406_n2088# a_n2406_n2088# a_n2406_n2088# a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X15 a_n2406_n2088# a_n2406_n2088# a_n2406_n2088# a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X16 source.t24 minus.t7 drain_right.t16 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X17 source.t36 minus.t8 drain_right.t15 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X18 source.t43 minus.t9 drain_right.t14 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X19 drain_right.t13 minus.t10 source.t45 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X20 drain_right.t12 minus.t11 source.t40 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X21 drain_right.t11 minus.t12 source.t42 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X22 source.t13 plus.t5 drain_left.t18 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X23 source.t44 minus.t13 drain_right.t10 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X24 drain_right.t9 minus.t14 source.t25 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X25 drain_right.t8 minus.t15 source.t31 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X26 drain_left.t17 plus.t6 source.t0 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X27 source.t4 plus.t7 drain_left.t16 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X28 drain_right.t7 minus.t16 source.t29 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X29 drain_right.t6 minus.t17 source.t46 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X30 source.t33 minus.t18 drain_right.t5 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X31 source.t5 plus.t8 drain_left.t15 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X32 source.t26 minus.t19 drain_right.t4 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X33 source.t32 minus.t20 drain_right.t3 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X34 source.t14 plus.t9 drain_left.t14 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X35 drain_left.t13 plus.t10 source.t21 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X36 source.t34 minus.t21 drain_right.t2 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X37 drain_left.t12 plus.t11 source.t1 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X38 drain_right.t1 minus.t22 source.t27 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X39 drain_left.t11 plus.t12 source.t9 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X40 source.t12 plus.t13 drain_left.t10 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X41 source.t15 plus.t14 drain_left.t9 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X42 source.t38 minus.t23 drain_right.t0 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X43 drain_left.t8 plus.t15 source.t20 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X44 source.t11 plus.t16 drain_left.t7 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X45 drain_left.t6 plus.t17 source.t16 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X46 drain_left.t5 plus.t18 source.t17 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X47 source.t22 plus.t19 drain_left.t4 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X48 drain_left.t3 plus.t20 source.t3 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X49 drain_left.t2 plus.t21 source.t8 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X50 source.t2 plus.t22 drain_left.t1 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X51 source.t6 plus.t23 drain_left.t0 a_n2406_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
R0 minus.n35 minus.t20 1220.34
R1 minus.n8 minus.t10 1220.34
R2 minus.n72 minus.t0 1220.34
R3 minus.n43 minus.t18 1220.34
R4 minus.n34 minus.t22 1172.87
R5 minus.n32 minus.t23 1172.87
R6 minus.n3 minus.t15 1172.87
R7 minus.n26 minus.t19 1172.87
R8 minus.n24 minus.t17 1172.87
R9 minus.n6 minus.t21 1172.87
R10 minus.n18 minus.t11 1172.87
R11 minus.n16 minus.t13 1172.87
R12 minus.n9 minus.t16 1172.87
R13 minus.n10 minus.t8 1172.87
R14 minus.n71 minus.t9 1172.87
R15 minus.n69 minus.t5 1172.87
R16 minus.n63 minus.t2 1172.87
R17 minus.n62 minus.t14 1172.87
R18 minus.n60 minus.t7 1172.87
R19 minus.n54 minus.t4 1172.87
R20 minus.n53 minus.t1 1172.87
R21 minus.n51 minus.t12 1172.87
R22 minus.n45 minus.t6 1172.87
R23 minus.n44 minus.t3 1172.87
R24 minus.n12 minus.n8 161.489
R25 minus.n47 minus.n43 161.489
R26 minus.n36 minus.n35 161.3
R27 minus.n33 minus.n0 161.3
R28 minus.n31 minus.n30 161.3
R29 minus.n29 minus.n1 161.3
R30 minus.n28 minus.n27 161.3
R31 minus.n25 minus.n2 161.3
R32 minus.n23 minus.n22 161.3
R33 minus.n21 minus.n4 161.3
R34 minus.n20 minus.n19 161.3
R35 minus.n17 minus.n5 161.3
R36 minus.n15 minus.n14 161.3
R37 minus.n13 minus.n7 161.3
R38 minus.n12 minus.n11 161.3
R39 minus.n73 minus.n72 161.3
R40 minus.n70 minus.n37 161.3
R41 minus.n68 minus.n67 161.3
R42 minus.n66 minus.n38 161.3
R43 minus.n65 minus.n64 161.3
R44 minus.n61 minus.n39 161.3
R45 minus.n59 minus.n58 161.3
R46 minus.n57 minus.n40 161.3
R47 minus.n56 minus.n55 161.3
R48 minus.n52 minus.n41 161.3
R49 minus.n50 minus.n49 161.3
R50 minus.n48 minus.n42 161.3
R51 minus.n47 minus.n46 161.3
R52 minus.n31 minus.n1 73.0308
R53 minus.n23 minus.n4 73.0308
R54 minus.n15 minus.n7 73.0308
R55 minus.n50 minus.n42 73.0308
R56 minus.n59 minus.n40 73.0308
R57 minus.n68 minus.n38 73.0308
R58 minus.n33 minus.n32 69.3793
R59 minus.n11 minus.n9 69.3793
R60 minus.n46 minus.n45 69.3793
R61 minus.n70 minus.n69 69.3793
R62 minus.n25 minus.n24 62.0763
R63 minus.n19 minus.n6 62.0763
R64 minus.n55 minus.n54 62.0763
R65 minus.n61 minus.n60 62.0763
R66 minus.n27 minus.n3 54.7732
R67 minus.n17 minus.n16 54.7732
R68 minus.n52 minus.n51 54.7732
R69 minus.n64 minus.n63 54.7732
R70 minus.n35 minus.n34 47.4702
R71 minus.n10 minus.n8 47.4702
R72 minus.n44 minus.n43 47.4702
R73 minus.n72 minus.n71 47.4702
R74 minus.n27 minus.n26 40.1672
R75 minus.n18 minus.n17 40.1672
R76 minus.n53 minus.n52 40.1672
R77 minus.n64 minus.n62 40.1672
R78 minus.n74 minus.n36 33.7126
R79 minus.n26 minus.n25 32.8641
R80 minus.n19 minus.n18 32.8641
R81 minus.n55 minus.n53 32.8641
R82 minus.n62 minus.n61 32.8641
R83 minus.n34 minus.n33 25.5611
R84 minus.n11 minus.n10 25.5611
R85 minus.n46 minus.n44 25.5611
R86 minus.n71 minus.n70 25.5611
R87 minus.n3 minus.n1 18.2581
R88 minus.n16 minus.n15 18.2581
R89 minus.n51 minus.n50 18.2581
R90 minus.n63 minus.n38 18.2581
R91 minus.n24 minus.n23 10.955
R92 minus.n6 minus.n4 10.955
R93 minus.n54 minus.n40 10.955
R94 minus.n60 minus.n59 10.955
R95 minus.n74 minus.n73 6.52323
R96 minus.n32 minus.n31 3.65202
R97 minus.n9 minus.n7 3.65202
R98 minus.n45 minus.n42 3.65202
R99 minus.n69 minus.n68 3.65202
R100 minus.n36 minus.n0 0.189894
R101 minus.n30 minus.n0 0.189894
R102 minus.n30 minus.n29 0.189894
R103 minus.n29 minus.n28 0.189894
R104 minus.n28 minus.n2 0.189894
R105 minus.n22 minus.n2 0.189894
R106 minus.n22 minus.n21 0.189894
R107 minus.n21 minus.n20 0.189894
R108 minus.n20 minus.n5 0.189894
R109 minus.n14 minus.n5 0.189894
R110 minus.n14 minus.n13 0.189894
R111 minus.n13 minus.n12 0.189894
R112 minus.n48 minus.n47 0.189894
R113 minus.n49 minus.n48 0.189894
R114 minus.n49 minus.n41 0.189894
R115 minus.n56 minus.n41 0.189894
R116 minus.n57 minus.n56 0.189894
R117 minus.n58 minus.n57 0.189894
R118 minus.n58 minus.n39 0.189894
R119 minus.n65 minus.n39 0.189894
R120 minus.n66 minus.n65 0.189894
R121 minus.n67 minus.n66 0.189894
R122 minus.n67 minus.n37 0.189894
R123 minus.n73 minus.n37 0.189894
R124 minus minus.n74 0.188
R125 source.n11 source.t4 55.512
R126 source.n12 source.t45 55.512
R127 source.n23 source.t32 55.512
R128 source.n0 source.t8 55.5119
R129 source.n47 source.t30 55.5119
R130 source.n36 source.t33 55.5119
R131 source.n35 source.t7 55.5119
R132 source.n24 source.t6 55.5119
R133 source.n2 source.n1 50.512
R134 source.n4 source.n3 50.512
R135 source.n6 source.n5 50.512
R136 source.n8 source.n7 50.512
R137 source.n10 source.n9 50.512
R138 source.n14 source.n13 50.512
R139 source.n16 source.n15 50.512
R140 source.n18 source.n17 50.512
R141 source.n20 source.n19 50.512
R142 source.n22 source.n21 50.512
R143 source.n46 source.n45 50.5119
R144 source.n44 source.n43 50.5119
R145 source.n42 source.n41 50.5119
R146 source.n40 source.n39 50.5119
R147 source.n38 source.n37 50.5119
R148 source.n34 source.n33 50.5119
R149 source.n32 source.n31 50.5119
R150 source.n30 source.n29 50.5119
R151 source.n28 source.n27 50.5119
R152 source.n26 source.n25 50.5119
R153 source.n24 source.n23 17.3026
R154 source.n48 source.n0 11.7595
R155 source.n48 source.n47 5.5436
R156 source.n45 source.t41 5.0005
R157 source.n45 source.t43 5.0005
R158 source.n43 source.t25 5.0005
R159 source.n43 source.t37 5.0005
R160 source.n41 source.t39 5.0005
R161 source.n41 source.t24 5.0005
R162 source.n39 source.t42 5.0005
R163 source.n39 source.t28 5.0005
R164 source.n37 source.t47 5.0005
R165 source.n37 source.t35 5.0005
R166 source.n33 source.t20 5.0005
R167 source.n33 source.t23 5.0005
R168 source.n31 source.t19 5.0005
R169 source.n31 source.t18 5.0005
R170 source.n29 source.t3 5.0005
R171 source.n29 source.t14 5.0005
R172 source.n27 source.t10 5.0005
R173 source.n27 source.t22 5.0005
R174 source.n25 source.t1 5.0005
R175 source.n25 source.t13 5.0005
R176 source.n1 source.t9 5.0005
R177 source.n1 source.t5 5.0005
R178 source.n3 source.t0 5.0005
R179 source.n3 source.t11 5.0005
R180 source.n5 source.t16 5.0005
R181 source.n5 source.t12 5.0005
R182 source.n7 source.t21 5.0005
R183 source.n7 source.t2 5.0005
R184 source.n9 source.t17 5.0005
R185 source.n9 source.t15 5.0005
R186 source.n13 source.t29 5.0005
R187 source.n13 source.t36 5.0005
R188 source.n15 source.t40 5.0005
R189 source.n15 source.t44 5.0005
R190 source.n17 source.t46 5.0005
R191 source.n17 source.t34 5.0005
R192 source.n19 source.t31 5.0005
R193 source.n19 source.t26 5.0005
R194 source.n21 source.t27 5.0005
R195 source.n21 source.t38 5.0005
R196 source.n23 source.n22 0.560845
R197 source.n22 source.n20 0.560845
R198 source.n20 source.n18 0.560845
R199 source.n18 source.n16 0.560845
R200 source.n16 source.n14 0.560845
R201 source.n14 source.n12 0.560845
R202 source.n11 source.n10 0.560845
R203 source.n10 source.n8 0.560845
R204 source.n8 source.n6 0.560845
R205 source.n6 source.n4 0.560845
R206 source.n4 source.n2 0.560845
R207 source.n2 source.n0 0.560845
R208 source.n26 source.n24 0.560845
R209 source.n28 source.n26 0.560845
R210 source.n30 source.n28 0.560845
R211 source.n32 source.n30 0.560845
R212 source.n34 source.n32 0.560845
R213 source.n35 source.n34 0.560845
R214 source.n38 source.n36 0.560845
R215 source.n40 source.n38 0.560845
R216 source.n42 source.n40 0.560845
R217 source.n44 source.n42 0.560845
R218 source.n46 source.n44 0.560845
R219 source.n47 source.n46 0.560845
R220 source.n12 source.n11 0.470328
R221 source.n36 source.n35 0.470328
R222 source source.n48 0.188
R223 drain_right.n13 drain_right.n11 67.751
R224 drain_right.n7 drain_right.n5 67.751
R225 drain_right.n2 drain_right.n0 67.751
R226 drain_right.n13 drain_right.n12 67.1908
R227 drain_right.n15 drain_right.n14 67.1908
R228 drain_right.n17 drain_right.n16 67.1908
R229 drain_right.n19 drain_right.n18 67.1908
R230 drain_right.n21 drain_right.n20 67.1908
R231 drain_right.n7 drain_right.n6 67.1907
R232 drain_right.n9 drain_right.n8 67.1907
R233 drain_right.n4 drain_right.n3 67.1907
R234 drain_right.n2 drain_right.n1 67.1907
R235 drain_right drain_right.n10 27.5917
R236 drain_right drain_right.n21 6.21356
R237 drain_right.n5 drain_right.t14 5.0005
R238 drain_right.n5 drain_right.t23 5.0005
R239 drain_right.n6 drain_right.t21 5.0005
R240 drain_right.n6 drain_right.t18 5.0005
R241 drain_right.n8 drain_right.t16 5.0005
R242 drain_right.n8 drain_right.t9 5.0005
R243 drain_right.n3 drain_right.t22 5.0005
R244 drain_right.n3 drain_right.t19 5.0005
R245 drain_right.n1 drain_right.t17 5.0005
R246 drain_right.n1 drain_right.t11 5.0005
R247 drain_right.n0 drain_right.t5 5.0005
R248 drain_right.n0 drain_right.t20 5.0005
R249 drain_right.n11 drain_right.t15 5.0005
R250 drain_right.n11 drain_right.t13 5.0005
R251 drain_right.n12 drain_right.t10 5.0005
R252 drain_right.n12 drain_right.t7 5.0005
R253 drain_right.n14 drain_right.t2 5.0005
R254 drain_right.n14 drain_right.t12 5.0005
R255 drain_right.n16 drain_right.t4 5.0005
R256 drain_right.n16 drain_right.t6 5.0005
R257 drain_right.n18 drain_right.t0 5.0005
R258 drain_right.n18 drain_right.t8 5.0005
R259 drain_right.n20 drain_right.t3 5.0005
R260 drain_right.n20 drain_right.t1 5.0005
R261 drain_right.n9 drain_right.n7 0.560845
R262 drain_right.n4 drain_right.n2 0.560845
R263 drain_right.n21 drain_right.n19 0.560845
R264 drain_right.n19 drain_right.n17 0.560845
R265 drain_right.n17 drain_right.n15 0.560845
R266 drain_right.n15 drain_right.n13 0.560845
R267 drain_right.n10 drain_right.n9 0.225326
R268 drain_right.n10 drain_right.n4 0.225326
R269 plus.n6 plus.t7 1220.34
R270 plus.n35 plus.t21 1220.34
R271 plus.n45 plus.t2 1220.34
R272 plus.n72 plus.t23 1220.34
R273 plus.n7 plus.t18 1172.87
R274 plus.n8 plus.t14 1172.87
R275 plus.n14 plus.t10 1172.87
R276 plus.n16 plus.t22 1172.87
R277 plus.n17 plus.t17 1172.87
R278 plus.n23 plus.t13 1172.87
R279 plus.n25 plus.t6 1172.87
R280 plus.n26 plus.t16 1172.87
R281 plus.n32 plus.t12 1172.87
R282 plus.n34 plus.t8 1172.87
R283 plus.n47 plus.t4 1172.87
R284 plus.n46 plus.t15 1172.87
R285 plus.n53 plus.t0 1172.87
R286 plus.n55 plus.t3 1172.87
R287 plus.n43 plus.t9 1172.87
R288 plus.n61 plus.t20 1172.87
R289 plus.n63 plus.t19 1172.87
R290 plus.n40 plus.t1 1172.87
R291 plus.n69 plus.t5 1172.87
R292 plus.n71 plus.t11 1172.87
R293 plus.n10 plus.n6 161.489
R294 plus.n49 plus.n45 161.489
R295 plus.n10 plus.n9 161.3
R296 plus.n11 plus.n5 161.3
R297 plus.n13 plus.n12 161.3
R298 plus.n15 plus.n4 161.3
R299 plus.n19 plus.n18 161.3
R300 plus.n20 plus.n3 161.3
R301 plus.n22 plus.n21 161.3
R302 plus.n24 plus.n2 161.3
R303 plus.n28 plus.n27 161.3
R304 plus.n29 plus.n1 161.3
R305 plus.n31 plus.n30 161.3
R306 plus.n33 plus.n0 161.3
R307 plus.n36 plus.n35 161.3
R308 plus.n49 plus.n48 161.3
R309 plus.n50 plus.n44 161.3
R310 plus.n52 plus.n51 161.3
R311 plus.n54 plus.n42 161.3
R312 plus.n57 plus.n56 161.3
R313 plus.n58 plus.n41 161.3
R314 plus.n60 plus.n59 161.3
R315 plus.n62 plus.n39 161.3
R316 plus.n65 plus.n64 161.3
R317 plus.n66 plus.n38 161.3
R318 plus.n68 plus.n67 161.3
R319 plus.n70 plus.n37 161.3
R320 plus.n73 plus.n72 161.3
R321 plus.n13 plus.n5 73.0308
R322 plus.n22 plus.n3 73.0308
R323 plus.n31 plus.n1 73.0308
R324 plus.n68 plus.n38 73.0308
R325 plus.n60 plus.n41 73.0308
R326 plus.n52 plus.n44 73.0308
R327 plus.n9 plus.n8 69.3793
R328 plus.n33 plus.n32 69.3793
R329 plus.n70 plus.n69 69.3793
R330 plus.n48 plus.n46 69.3793
R331 plus.n18 plus.n17 62.0763
R332 plus.n24 plus.n23 62.0763
R333 plus.n62 plus.n61 62.0763
R334 plus.n56 plus.n43 62.0763
R335 plus.n15 plus.n14 54.7732
R336 plus.n27 plus.n26 54.7732
R337 plus.n64 plus.n40 54.7732
R338 plus.n54 plus.n53 54.7732
R339 plus.n7 plus.n6 47.4702
R340 plus.n35 plus.n34 47.4702
R341 plus.n72 plus.n71 47.4702
R342 plus.n47 plus.n45 47.4702
R343 plus.n16 plus.n15 40.1672
R344 plus.n27 plus.n25 40.1672
R345 plus.n64 plus.n63 40.1672
R346 plus.n55 plus.n54 40.1672
R347 plus.n18 plus.n16 32.8641
R348 plus.n25 plus.n24 32.8641
R349 plus.n63 plus.n62 32.8641
R350 plus.n56 plus.n55 32.8641
R351 plus plus.n73 29.8664
R352 plus.n9 plus.n7 25.5611
R353 plus.n34 plus.n33 25.5611
R354 plus.n71 plus.n70 25.5611
R355 plus.n48 plus.n47 25.5611
R356 plus.n14 plus.n13 18.2581
R357 plus.n26 plus.n1 18.2581
R358 plus.n40 plus.n38 18.2581
R359 plus.n53 plus.n52 18.2581
R360 plus.n17 plus.n3 10.955
R361 plus.n23 plus.n22 10.955
R362 plus.n61 plus.n60 10.955
R363 plus.n43 plus.n41 10.955
R364 plus plus.n36 9.89444
R365 plus.n8 plus.n5 3.65202
R366 plus.n32 plus.n31 3.65202
R367 plus.n69 plus.n68 3.65202
R368 plus.n46 plus.n44 3.65202
R369 plus.n11 plus.n10 0.189894
R370 plus.n12 plus.n11 0.189894
R371 plus.n12 plus.n4 0.189894
R372 plus.n19 plus.n4 0.189894
R373 plus.n20 plus.n19 0.189894
R374 plus.n21 plus.n20 0.189894
R375 plus.n21 plus.n2 0.189894
R376 plus.n28 plus.n2 0.189894
R377 plus.n29 plus.n28 0.189894
R378 plus.n30 plus.n29 0.189894
R379 plus.n30 plus.n0 0.189894
R380 plus.n36 plus.n0 0.189894
R381 plus.n73 plus.n37 0.189894
R382 plus.n67 plus.n37 0.189894
R383 plus.n67 plus.n66 0.189894
R384 plus.n66 plus.n65 0.189894
R385 plus.n65 plus.n39 0.189894
R386 plus.n59 plus.n39 0.189894
R387 plus.n59 plus.n58 0.189894
R388 plus.n58 plus.n57 0.189894
R389 plus.n57 plus.n42 0.189894
R390 plus.n51 plus.n42 0.189894
R391 plus.n51 plus.n50 0.189894
R392 plus.n50 plus.n49 0.189894
R393 drain_left.n13 drain_left.n11 67.7512
R394 drain_left.n7 drain_left.n5 67.751
R395 drain_left.n2 drain_left.n0 67.751
R396 drain_left.n19 drain_left.n18 67.1908
R397 drain_left.n17 drain_left.n16 67.1908
R398 drain_left.n15 drain_left.n14 67.1908
R399 drain_left.n13 drain_left.n12 67.1908
R400 drain_left.n21 drain_left.n20 67.1907
R401 drain_left.n7 drain_left.n6 67.1907
R402 drain_left.n9 drain_left.n8 67.1907
R403 drain_left.n4 drain_left.n3 67.1907
R404 drain_left.n2 drain_left.n1 67.1907
R405 drain_left drain_left.n10 28.1449
R406 drain_left drain_left.n21 6.21356
R407 drain_left.n5 drain_left.t19 5.0005
R408 drain_left.n5 drain_left.t21 5.0005
R409 drain_left.n6 drain_left.t23 5.0005
R410 drain_left.n6 drain_left.t8 5.0005
R411 drain_left.n8 drain_left.t14 5.0005
R412 drain_left.n8 drain_left.t20 5.0005
R413 drain_left.n3 drain_left.t4 5.0005
R414 drain_left.n3 drain_left.t3 5.0005
R415 drain_left.n1 drain_left.t18 5.0005
R416 drain_left.n1 drain_left.t22 5.0005
R417 drain_left.n0 drain_left.t0 5.0005
R418 drain_left.n0 drain_left.t12 5.0005
R419 drain_left.n20 drain_left.t15 5.0005
R420 drain_left.n20 drain_left.t2 5.0005
R421 drain_left.n18 drain_left.t7 5.0005
R422 drain_left.n18 drain_left.t11 5.0005
R423 drain_left.n16 drain_left.t10 5.0005
R424 drain_left.n16 drain_left.t17 5.0005
R425 drain_left.n14 drain_left.t1 5.0005
R426 drain_left.n14 drain_left.t6 5.0005
R427 drain_left.n12 drain_left.t9 5.0005
R428 drain_left.n12 drain_left.t13 5.0005
R429 drain_left.n11 drain_left.t16 5.0005
R430 drain_left.n11 drain_left.t5 5.0005
R431 drain_left.n9 drain_left.n7 0.560845
R432 drain_left.n4 drain_left.n2 0.560845
R433 drain_left.n15 drain_left.n13 0.560845
R434 drain_left.n17 drain_left.n15 0.560845
R435 drain_left.n19 drain_left.n17 0.560845
R436 drain_left.n21 drain_left.n19 0.560845
R437 drain_left.n10 drain_left.n9 0.225326
R438 drain_left.n10 drain_left.n4 0.225326
C0 drain_right source 24.653f
C1 minus source 2.72677f
C2 drain_left plus 3.03881f
C3 plus drain_right 0.392113f
C4 drain_left drain_right 1.29455f
C5 plus minus 5.0304f
C6 drain_left minus 0.171476f
C7 drain_right minus 2.80103f
C8 plus source 2.74079f
C9 drain_left source 24.652302f
C10 drain_right a_n2406_n2088# 5.69685f
C11 drain_left a_n2406_n2088# 6.04656f
C12 source a_n2406_n2088# 5.673229f
C13 minus a_n2406_n2088# 8.420897f
C14 plus a_n2406_n2088# 10.20057f
C15 drain_left.t0 a_n2406_n2088# 0.204046f
C16 drain_left.t12 a_n2406_n2088# 0.204046f
C17 drain_left.n0 a_n2406_n2088# 1.26475f
C18 drain_left.t18 a_n2406_n2088# 0.204046f
C19 drain_left.t22 a_n2406_n2088# 0.204046f
C20 drain_left.n1 a_n2406_n2088# 1.2619f
C21 drain_left.n2 a_n2406_n2088# 0.674786f
C22 drain_left.t4 a_n2406_n2088# 0.204046f
C23 drain_left.t3 a_n2406_n2088# 0.204046f
C24 drain_left.n3 a_n2406_n2088# 1.2619f
C25 drain_left.n4 a_n2406_n2088# 0.305319f
C26 drain_left.t19 a_n2406_n2088# 0.204046f
C27 drain_left.t21 a_n2406_n2088# 0.204046f
C28 drain_left.n5 a_n2406_n2088# 1.26475f
C29 drain_left.t23 a_n2406_n2088# 0.204046f
C30 drain_left.t8 a_n2406_n2088# 0.204046f
C31 drain_left.n6 a_n2406_n2088# 1.2619f
C32 drain_left.n7 a_n2406_n2088# 0.674786f
C33 drain_left.t14 a_n2406_n2088# 0.204046f
C34 drain_left.t20 a_n2406_n2088# 0.204046f
C35 drain_left.n8 a_n2406_n2088# 1.2619f
C36 drain_left.n9 a_n2406_n2088# 0.305319f
C37 drain_left.n10 a_n2406_n2088# 1.18444f
C38 drain_left.t16 a_n2406_n2088# 0.204046f
C39 drain_left.t5 a_n2406_n2088# 0.204046f
C40 drain_left.n11 a_n2406_n2088# 1.26476f
C41 drain_left.t9 a_n2406_n2088# 0.204046f
C42 drain_left.t13 a_n2406_n2088# 0.204046f
C43 drain_left.n12 a_n2406_n2088# 1.26191f
C44 drain_left.n13 a_n2406_n2088# 0.674775f
C45 drain_left.t1 a_n2406_n2088# 0.204046f
C46 drain_left.t6 a_n2406_n2088# 0.204046f
C47 drain_left.n14 a_n2406_n2088# 1.26191f
C48 drain_left.n15 a_n2406_n2088# 0.333092f
C49 drain_left.t10 a_n2406_n2088# 0.204046f
C50 drain_left.t17 a_n2406_n2088# 0.204046f
C51 drain_left.n16 a_n2406_n2088# 1.26191f
C52 drain_left.n17 a_n2406_n2088# 0.333092f
C53 drain_left.t7 a_n2406_n2088# 0.204046f
C54 drain_left.t11 a_n2406_n2088# 0.204046f
C55 drain_left.n18 a_n2406_n2088# 1.26191f
C56 drain_left.n19 a_n2406_n2088# 0.333092f
C57 drain_left.t15 a_n2406_n2088# 0.204046f
C58 drain_left.t2 a_n2406_n2088# 0.204046f
C59 drain_left.n20 a_n2406_n2088# 1.2619f
C60 drain_left.n21 a_n2406_n2088# 0.570295f
C61 plus.n0 a_n2406_n2088# 0.0518f
C62 plus.t8 a_n2406_n2088# 0.132829f
C63 plus.t12 a_n2406_n2088# 0.132829f
C64 plus.n1 a_n2406_n2088# 0.021176f
C65 plus.n2 a_n2406_n2088# 0.0518f
C66 plus.t6 a_n2406_n2088# 0.132829f
C67 plus.t13 a_n2406_n2088# 0.132829f
C68 plus.n3 a_n2406_n2088# 0.019579f
C69 plus.n4 a_n2406_n2088# 0.0518f
C70 plus.t22 a_n2406_n2088# 0.132829f
C71 plus.t10 a_n2406_n2088# 0.132829f
C72 plus.n5 a_n2406_n2088# 0.017982f
C73 plus.t7 a_n2406_n2088# 0.13548f
C74 plus.n6 a_n2406_n2088# 0.087552f
C75 plus.t18 a_n2406_n2088# 0.132829f
C76 plus.n7 a_n2406_n2088# 0.068955f
C77 plus.t14 a_n2406_n2088# 0.132829f
C78 plus.n8 a_n2406_n2088# 0.068955f
C79 plus.n9 a_n2406_n2088# 0.021974f
C80 plus.n10 a_n2406_n2088# 0.11311f
C81 plus.n11 a_n2406_n2088# 0.0518f
C82 plus.n12 a_n2406_n2088# 0.0518f
C83 plus.n13 a_n2406_n2088# 0.021176f
C84 plus.n14 a_n2406_n2088# 0.068955f
C85 plus.n15 a_n2406_n2088# 0.021974f
C86 plus.n16 a_n2406_n2088# 0.068955f
C87 plus.t17 a_n2406_n2088# 0.132829f
C88 plus.n17 a_n2406_n2088# 0.068955f
C89 plus.n18 a_n2406_n2088# 0.021974f
C90 plus.n19 a_n2406_n2088# 0.0518f
C91 plus.n20 a_n2406_n2088# 0.0518f
C92 plus.n21 a_n2406_n2088# 0.0518f
C93 plus.n22 a_n2406_n2088# 0.019579f
C94 plus.n23 a_n2406_n2088# 0.068955f
C95 plus.n24 a_n2406_n2088# 0.021974f
C96 plus.n25 a_n2406_n2088# 0.068955f
C97 plus.t16 a_n2406_n2088# 0.132829f
C98 plus.n26 a_n2406_n2088# 0.068955f
C99 plus.n27 a_n2406_n2088# 0.021974f
C100 plus.n28 a_n2406_n2088# 0.0518f
C101 plus.n29 a_n2406_n2088# 0.0518f
C102 plus.n30 a_n2406_n2088# 0.0518f
C103 plus.n31 a_n2406_n2088# 0.017982f
C104 plus.n32 a_n2406_n2088# 0.068955f
C105 plus.n33 a_n2406_n2088# 0.021974f
C106 plus.n34 a_n2406_n2088# 0.068955f
C107 plus.t21 a_n2406_n2088# 0.13548f
C108 plus.n35 a_n2406_n2088# 0.08748f
C109 plus.n36 a_n2406_n2088# 0.446827f
C110 plus.n37 a_n2406_n2088# 0.0518f
C111 plus.t23 a_n2406_n2088# 0.13548f
C112 plus.t11 a_n2406_n2088# 0.132829f
C113 plus.t5 a_n2406_n2088# 0.132829f
C114 plus.n38 a_n2406_n2088# 0.021176f
C115 plus.n39 a_n2406_n2088# 0.0518f
C116 plus.t1 a_n2406_n2088# 0.132829f
C117 plus.n40 a_n2406_n2088# 0.068955f
C118 plus.t19 a_n2406_n2088# 0.132829f
C119 plus.t20 a_n2406_n2088# 0.132829f
C120 plus.n41 a_n2406_n2088# 0.019579f
C121 plus.n42 a_n2406_n2088# 0.0518f
C122 plus.t9 a_n2406_n2088# 0.132829f
C123 plus.n43 a_n2406_n2088# 0.068955f
C124 plus.t3 a_n2406_n2088# 0.132829f
C125 plus.t0 a_n2406_n2088# 0.132829f
C126 plus.n44 a_n2406_n2088# 0.017982f
C127 plus.t2 a_n2406_n2088# 0.13548f
C128 plus.n45 a_n2406_n2088# 0.087552f
C129 plus.t15 a_n2406_n2088# 0.132829f
C130 plus.n46 a_n2406_n2088# 0.068955f
C131 plus.t4 a_n2406_n2088# 0.132829f
C132 plus.n47 a_n2406_n2088# 0.068955f
C133 plus.n48 a_n2406_n2088# 0.021974f
C134 plus.n49 a_n2406_n2088# 0.11311f
C135 plus.n50 a_n2406_n2088# 0.0518f
C136 plus.n51 a_n2406_n2088# 0.0518f
C137 plus.n52 a_n2406_n2088# 0.021176f
C138 plus.n53 a_n2406_n2088# 0.068955f
C139 plus.n54 a_n2406_n2088# 0.021974f
C140 plus.n55 a_n2406_n2088# 0.068955f
C141 plus.n56 a_n2406_n2088# 0.021974f
C142 plus.n57 a_n2406_n2088# 0.0518f
C143 plus.n58 a_n2406_n2088# 0.0518f
C144 plus.n59 a_n2406_n2088# 0.0518f
C145 plus.n60 a_n2406_n2088# 0.019579f
C146 plus.n61 a_n2406_n2088# 0.068955f
C147 plus.n62 a_n2406_n2088# 0.021974f
C148 plus.n63 a_n2406_n2088# 0.068955f
C149 plus.n64 a_n2406_n2088# 0.021974f
C150 plus.n65 a_n2406_n2088# 0.0518f
C151 plus.n66 a_n2406_n2088# 0.0518f
C152 plus.n67 a_n2406_n2088# 0.0518f
C153 plus.n68 a_n2406_n2088# 0.017982f
C154 plus.n69 a_n2406_n2088# 0.068955f
C155 plus.n70 a_n2406_n2088# 0.021974f
C156 plus.n71 a_n2406_n2088# 0.068955f
C157 plus.n72 a_n2406_n2088# 0.08748f
C158 plus.n73 a_n2406_n2088# 1.47973f
C159 drain_right.t5 a_n2406_n2088# 0.203389f
C160 drain_right.t20 a_n2406_n2088# 0.203389f
C161 drain_right.n0 a_n2406_n2088# 1.26068f
C162 drain_right.t17 a_n2406_n2088# 0.203389f
C163 drain_right.t11 a_n2406_n2088# 0.203389f
C164 drain_right.n1 a_n2406_n2088# 1.25784f
C165 drain_right.n2 a_n2406_n2088# 0.672612f
C166 drain_right.t22 a_n2406_n2088# 0.203389f
C167 drain_right.t19 a_n2406_n2088# 0.203389f
C168 drain_right.n3 a_n2406_n2088# 1.25784f
C169 drain_right.n4 a_n2406_n2088# 0.304336f
C170 drain_right.t14 a_n2406_n2088# 0.203389f
C171 drain_right.t23 a_n2406_n2088# 0.203389f
C172 drain_right.n5 a_n2406_n2088# 1.26068f
C173 drain_right.t21 a_n2406_n2088# 0.203389f
C174 drain_right.t18 a_n2406_n2088# 0.203389f
C175 drain_right.n6 a_n2406_n2088# 1.25784f
C176 drain_right.n7 a_n2406_n2088# 0.672612f
C177 drain_right.t16 a_n2406_n2088# 0.203389f
C178 drain_right.t9 a_n2406_n2088# 0.203389f
C179 drain_right.n8 a_n2406_n2088# 1.25784f
C180 drain_right.n9 a_n2406_n2088# 0.304336f
C181 drain_right.n10 a_n2406_n2088# 1.12367f
C182 drain_right.t15 a_n2406_n2088# 0.203389f
C183 drain_right.t13 a_n2406_n2088# 0.203389f
C184 drain_right.n11 a_n2406_n2088# 1.26068f
C185 drain_right.t10 a_n2406_n2088# 0.203389f
C186 drain_right.t7 a_n2406_n2088# 0.203389f
C187 drain_right.n12 a_n2406_n2088# 1.25784f
C188 drain_right.n13 a_n2406_n2088# 0.672607f
C189 drain_right.t2 a_n2406_n2088# 0.203389f
C190 drain_right.t12 a_n2406_n2088# 0.203389f
C191 drain_right.n14 a_n2406_n2088# 1.25784f
C192 drain_right.n15 a_n2406_n2088# 0.332019f
C193 drain_right.t4 a_n2406_n2088# 0.203389f
C194 drain_right.t6 a_n2406_n2088# 0.203389f
C195 drain_right.n16 a_n2406_n2088# 1.25784f
C196 drain_right.n17 a_n2406_n2088# 0.332019f
C197 drain_right.t0 a_n2406_n2088# 0.203389f
C198 drain_right.t8 a_n2406_n2088# 0.203389f
C199 drain_right.n18 a_n2406_n2088# 1.25784f
C200 drain_right.n19 a_n2406_n2088# 0.332019f
C201 drain_right.t3 a_n2406_n2088# 0.203389f
C202 drain_right.t1 a_n2406_n2088# 0.203389f
C203 drain_right.n20 a_n2406_n2088# 1.25784f
C204 drain_right.n21 a_n2406_n2088# 0.568452f
C205 source.t8 a_n2406_n2088# 1.34405f
C206 source.n0 a_n2406_n2088# 0.988789f
C207 source.t9 a_n2406_n2088# 0.191357f
C208 source.t5 a_n2406_n2088# 0.191357f
C209 source.n1 a_n2406_n2088# 1.11372f
C210 source.n2 a_n2406_n2088# 0.345883f
C211 source.t0 a_n2406_n2088# 0.191357f
C212 source.t11 a_n2406_n2088# 0.191357f
C213 source.n3 a_n2406_n2088# 1.11372f
C214 source.n4 a_n2406_n2088# 0.345883f
C215 source.t16 a_n2406_n2088# 0.191357f
C216 source.t12 a_n2406_n2088# 0.191357f
C217 source.n5 a_n2406_n2088# 1.11372f
C218 source.n6 a_n2406_n2088# 0.345883f
C219 source.t21 a_n2406_n2088# 0.191357f
C220 source.t2 a_n2406_n2088# 0.191357f
C221 source.n7 a_n2406_n2088# 1.11372f
C222 source.n8 a_n2406_n2088# 0.345883f
C223 source.t17 a_n2406_n2088# 0.191357f
C224 source.t15 a_n2406_n2088# 0.191357f
C225 source.n9 a_n2406_n2088# 1.11372f
C226 source.n10 a_n2406_n2088# 0.345883f
C227 source.t4 a_n2406_n2088# 1.34406f
C228 source.n11 a_n2406_n2088# 0.452217f
C229 source.t45 a_n2406_n2088# 1.34406f
C230 source.n12 a_n2406_n2088# 0.452217f
C231 source.t29 a_n2406_n2088# 0.191357f
C232 source.t36 a_n2406_n2088# 0.191357f
C233 source.n13 a_n2406_n2088# 1.11372f
C234 source.n14 a_n2406_n2088# 0.345883f
C235 source.t40 a_n2406_n2088# 0.191357f
C236 source.t44 a_n2406_n2088# 0.191357f
C237 source.n15 a_n2406_n2088# 1.11372f
C238 source.n16 a_n2406_n2088# 0.345883f
C239 source.t46 a_n2406_n2088# 0.191357f
C240 source.t34 a_n2406_n2088# 0.191357f
C241 source.n17 a_n2406_n2088# 1.11372f
C242 source.n18 a_n2406_n2088# 0.345883f
C243 source.t31 a_n2406_n2088# 0.191357f
C244 source.t26 a_n2406_n2088# 0.191357f
C245 source.n19 a_n2406_n2088# 1.11372f
C246 source.n20 a_n2406_n2088# 0.345883f
C247 source.t27 a_n2406_n2088# 0.191357f
C248 source.t38 a_n2406_n2088# 0.191357f
C249 source.n21 a_n2406_n2088# 1.11372f
C250 source.n22 a_n2406_n2088# 0.345883f
C251 source.t32 a_n2406_n2088# 1.34406f
C252 source.n23 a_n2406_n2088# 1.33213f
C253 source.t6 a_n2406_n2088# 1.34405f
C254 source.n24 a_n2406_n2088# 1.33213f
C255 source.t1 a_n2406_n2088# 0.191357f
C256 source.t13 a_n2406_n2088# 0.191357f
C257 source.n25 a_n2406_n2088# 1.11371f
C258 source.n26 a_n2406_n2088# 0.34589f
C259 source.t10 a_n2406_n2088# 0.191357f
C260 source.t22 a_n2406_n2088# 0.191357f
C261 source.n27 a_n2406_n2088# 1.11371f
C262 source.n28 a_n2406_n2088# 0.34589f
C263 source.t3 a_n2406_n2088# 0.191357f
C264 source.t14 a_n2406_n2088# 0.191357f
C265 source.n29 a_n2406_n2088# 1.11371f
C266 source.n30 a_n2406_n2088# 0.34589f
C267 source.t19 a_n2406_n2088# 0.191357f
C268 source.t18 a_n2406_n2088# 0.191357f
C269 source.n31 a_n2406_n2088# 1.11371f
C270 source.n32 a_n2406_n2088# 0.34589f
C271 source.t20 a_n2406_n2088# 0.191357f
C272 source.t23 a_n2406_n2088# 0.191357f
C273 source.n33 a_n2406_n2088# 1.11371f
C274 source.n34 a_n2406_n2088# 0.34589f
C275 source.t7 a_n2406_n2088# 1.34405f
C276 source.n35 a_n2406_n2088# 0.452224f
C277 source.t33 a_n2406_n2088# 1.34405f
C278 source.n36 a_n2406_n2088# 0.452224f
C279 source.t47 a_n2406_n2088# 0.191357f
C280 source.t35 a_n2406_n2088# 0.191357f
C281 source.n37 a_n2406_n2088# 1.11371f
C282 source.n38 a_n2406_n2088# 0.34589f
C283 source.t42 a_n2406_n2088# 0.191357f
C284 source.t28 a_n2406_n2088# 0.191357f
C285 source.n39 a_n2406_n2088# 1.11371f
C286 source.n40 a_n2406_n2088# 0.34589f
C287 source.t39 a_n2406_n2088# 0.191357f
C288 source.t24 a_n2406_n2088# 0.191357f
C289 source.n41 a_n2406_n2088# 1.11371f
C290 source.n42 a_n2406_n2088# 0.34589f
C291 source.t25 a_n2406_n2088# 0.191357f
C292 source.t37 a_n2406_n2088# 0.191357f
C293 source.n43 a_n2406_n2088# 1.11371f
C294 source.n44 a_n2406_n2088# 0.34589f
C295 source.t41 a_n2406_n2088# 0.191357f
C296 source.t43 a_n2406_n2088# 0.191357f
C297 source.n45 a_n2406_n2088# 1.11371f
C298 source.n46 a_n2406_n2088# 0.34589f
C299 source.t30 a_n2406_n2088# 1.34405f
C300 source.n47 a_n2406_n2088# 0.603771f
C301 source.n48 a_n2406_n2088# 1.09065f
C302 minus.n0 a_n2406_n2088# 0.050339f
C303 minus.t20 a_n2406_n2088# 0.131659f
C304 minus.t22 a_n2406_n2088# 0.129083f
C305 minus.t23 a_n2406_n2088# 0.129083f
C306 minus.n1 a_n2406_n2088# 0.020579f
C307 minus.n2 a_n2406_n2088# 0.050339f
C308 minus.t15 a_n2406_n2088# 0.129083f
C309 minus.n3 a_n2406_n2088# 0.06701f
C310 minus.t19 a_n2406_n2088# 0.129083f
C311 minus.t17 a_n2406_n2088# 0.129083f
C312 minus.n4 a_n2406_n2088# 0.019027f
C313 minus.n5 a_n2406_n2088# 0.050339f
C314 minus.t21 a_n2406_n2088# 0.129083f
C315 minus.n6 a_n2406_n2088# 0.06701f
C316 minus.t11 a_n2406_n2088# 0.129083f
C317 minus.t13 a_n2406_n2088# 0.129083f
C318 minus.n7 a_n2406_n2088# 0.017475f
C319 minus.t10 a_n2406_n2088# 0.131659f
C320 minus.n8 a_n2406_n2088# 0.085082f
C321 minus.t16 a_n2406_n2088# 0.129083f
C322 minus.n9 a_n2406_n2088# 0.06701f
C323 minus.t8 a_n2406_n2088# 0.129083f
C324 minus.n10 a_n2406_n2088# 0.06701f
C325 minus.n11 a_n2406_n2088# 0.021355f
C326 minus.n12 a_n2406_n2088# 0.109919f
C327 minus.n13 a_n2406_n2088# 0.050339f
C328 minus.n14 a_n2406_n2088# 0.050339f
C329 minus.n15 a_n2406_n2088# 0.020579f
C330 minus.n16 a_n2406_n2088# 0.06701f
C331 minus.n17 a_n2406_n2088# 0.021355f
C332 minus.n18 a_n2406_n2088# 0.06701f
C333 minus.n19 a_n2406_n2088# 0.021355f
C334 minus.n20 a_n2406_n2088# 0.050339f
C335 minus.n21 a_n2406_n2088# 0.050339f
C336 minus.n22 a_n2406_n2088# 0.050339f
C337 minus.n23 a_n2406_n2088# 0.019027f
C338 minus.n24 a_n2406_n2088# 0.06701f
C339 minus.n25 a_n2406_n2088# 0.021355f
C340 minus.n26 a_n2406_n2088# 0.06701f
C341 minus.n27 a_n2406_n2088# 0.021355f
C342 minus.n28 a_n2406_n2088# 0.050339f
C343 minus.n29 a_n2406_n2088# 0.050339f
C344 minus.n30 a_n2406_n2088# 0.050339f
C345 minus.n31 a_n2406_n2088# 0.017475f
C346 minus.n32 a_n2406_n2088# 0.06701f
C347 minus.n33 a_n2406_n2088# 0.021355f
C348 minus.n34 a_n2406_n2088# 0.06701f
C349 minus.n35 a_n2406_n2088# 0.085012f
C350 minus.n36 a_n2406_n2088# 1.59025f
C351 minus.n37 a_n2406_n2088# 0.050339f
C352 minus.t9 a_n2406_n2088# 0.129083f
C353 minus.t5 a_n2406_n2088# 0.129083f
C354 minus.n38 a_n2406_n2088# 0.020579f
C355 minus.n39 a_n2406_n2088# 0.050339f
C356 minus.t14 a_n2406_n2088# 0.129083f
C357 minus.t7 a_n2406_n2088# 0.129083f
C358 minus.n40 a_n2406_n2088# 0.019027f
C359 minus.n41 a_n2406_n2088# 0.050339f
C360 minus.t1 a_n2406_n2088# 0.129083f
C361 minus.t12 a_n2406_n2088# 0.129083f
C362 minus.n42 a_n2406_n2088# 0.017475f
C363 minus.t18 a_n2406_n2088# 0.131659f
C364 minus.n43 a_n2406_n2088# 0.085082f
C365 minus.t3 a_n2406_n2088# 0.129083f
C366 minus.n44 a_n2406_n2088# 0.06701f
C367 minus.t6 a_n2406_n2088# 0.129083f
C368 minus.n45 a_n2406_n2088# 0.06701f
C369 minus.n46 a_n2406_n2088# 0.021355f
C370 minus.n47 a_n2406_n2088# 0.109919f
C371 minus.n48 a_n2406_n2088# 0.050339f
C372 minus.n49 a_n2406_n2088# 0.050339f
C373 minus.n50 a_n2406_n2088# 0.020579f
C374 minus.n51 a_n2406_n2088# 0.06701f
C375 minus.n52 a_n2406_n2088# 0.021355f
C376 minus.n53 a_n2406_n2088# 0.06701f
C377 minus.t4 a_n2406_n2088# 0.129083f
C378 minus.n54 a_n2406_n2088# 0.06701f
C379 minus.n55 a_n2406_n2088# 0.021355f
C380 minus.n56 a_n2406_n2088# 0.050339f
C381 minus.n57 a_n2406_n2088# 0.050339f
C382 minus.n58 a_n2406_n2088# 0.050339f
C383 minus.n59 a_n2406_n2088# 0.019027f
C384 minus.n60 a_n2406_n2088# 0.06701f
C385 minus.n61 a_n2406_n2088# 0.021355f
C386 minus.n62 a_n2406_n2088# 0.06701f
C387 minus.t2 a_n2406_n2088# 0.129083f
C388 minus.n63 a_n2406_n2088# 0.06701f
C389 minus.n64 a_n2406_n2088# 0.021355f
C390 minus.n65 a_n2406_n2088# 0.050339f
C391 minus.n66 a_n2406_n2088# 0.050339f
C392 minus.n67 a_n2406_n2088# 0.050339f
C393 minus.n68 a_n2406_n2088# 0.017475f
C394 minus.n69 a_n2406_n2088# 0.06701f
C395 minus.n70 a_n2406_n2088# 0.021355f
C396 minus.n71 a_n2406_n2088# 0.06701f
C397 minus.t0 a_n2406_n2088# 0.131659f
C398 minus.n72 a_n2406_n2088# 0.085012f
C399 minus.n73 a_n2406_n2088# 0.331856f
C400 minus.n74 a_n2406_n2088# 1.94427f
.ends

