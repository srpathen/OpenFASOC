* NGSPICE file created from opamp197.ext - technology: sky130A

.subckt opamp197 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X2 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X4 a_n2472_13878# a_n2650_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 outputibias outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X7 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=337.44 ps=1.95024k w=7 l=1
X8 a_n8964_8799# plus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X9 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X10 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X11 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 CSoutput a_n2650_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X13 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 minus gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X16 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X17 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X22 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 outputibias outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X25 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X27 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 a_n2650_13878# minus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X29 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 a_n8964_8799# plus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X31 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X32 a_n2650_13878# minus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X33 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X36 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X40 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X41 a_n2903_n3924# plus a_n8964_8799# gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X42 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 a_n2903_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X45 a_n2903_n3924# minus a_n2650_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X46 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X51 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=348.84 ps=2.0286k w=9 l=0.5
X52 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 outputibias outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X54 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X55 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X56 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X59 CSoutput a_n2650_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X60 gnd gnd plus gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X61 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X63 a_n2903_n3924# plus a_n8964_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X64 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X67 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X68 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X70 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X71 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X74 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X77 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X79 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X82 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X85 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 a_n2903_n3924# minus a_n2650_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X89 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X90 a_n2903_n3924# plus a_n8964_8799# gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X91 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X95 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 a_n2903_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X97 CSoutput a_n2650_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X98 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X101 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X102 a_n2903_n3924# plus a_n8964_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X103 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X105 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X106 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X107 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X112 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X114 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X115 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X117 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X119 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X121 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 vdd a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 gnd gnd minus gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X127 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X128 a_n2650_8322# a_n2650_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 a_n2903_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X130 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X134 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 vdd a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X137 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X138 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X140 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X142 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 outputibias outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X144 a_n8964_8799# plus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X145 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X146 a_n2650_8322# a_n2650_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X147 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X148 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X152 a_n8964_8799# plus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X153 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X155 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X159 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X160 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X162 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X164 output outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X165 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X166 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X170 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X171 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 vdd a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X174 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X175 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X177 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X178 a_n2650_13878# minus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X179 a_n2903_n3924# plus a_n8964_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X180 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X181 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X182 plus gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X183 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 a_n2903_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 gnd gnd minus gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X187 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X188 a_n2903_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X189 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X190 a_n8964_8799# plus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X191 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X192 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X195 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X196 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X197 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X199 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X202 a_n8964_8799# plus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X203 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X204 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X205 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X206 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X211 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X212 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X214 a_n2472_13878# a_n2650_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X215 a_n2650_13878# minus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X216 vdd a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X217 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 a_n2903_n3924# plus a_n8964_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X219 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X220 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X222 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X224 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X226 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X229 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 a_n2903_n3924# minus a_n2650_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X231 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X232 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X233 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X234 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X236 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X239 vdd a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X240 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X243 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 plus gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X245 gnd gnd minus gnd sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X246 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X249 a_n2472_13878# a_n2650_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X250 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X251 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X253 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X257 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X258 a_n2903_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X259 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X261 vdd a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X262 CSoutput a_n2650_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X263 a_n8964_8799# plus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X264 a_n2650_13878# minus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X265 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X268 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 a_n2903_n3924# minus a_n2650_13878# gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X270 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X271 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X276 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X277 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X279 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X282 a_n2903_n3924# minus a_n2650_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X283 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X284 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X286 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 a_n2903_n3924# minus a_n2650_13878# gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X288 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X289 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X292 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X294 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X295 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X296 CSoutput a_n2650_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X297 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X304 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X305 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X306 a_n2650_8322# a_n2650_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X307 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X310 a_n2903_n3924# minus a_n2650_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X311 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X313 output outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X314 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 vdd a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X317 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X320 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X322 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X323 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 output outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X331 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X332 gnd gnd plus gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X333 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X334 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X335 a_n2472_13878# a_n2650_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X336 output outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X337 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X338 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X339 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X341 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X344 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X345 a_n2903_n3924# plus a_n8964_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X346 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X347 a_n2650_13878# minus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X348 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X350 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X351 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X356 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X357 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X360 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X361 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 a_n2903_n3924# minus a_n2650_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X364 a_n2903_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X365 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X366 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X367 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X369 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X372 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 a_n8964_8799# a_n2650_13878# a_n2650_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X374 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X375 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X377 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X379 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X380 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 gnd gnd plus gnd sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X382 minus gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X383 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X385 a_n2650_13878# minus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X386 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X390 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X391 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X392 CSoutput a_n2650_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X393 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X394 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X395 vdd a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X396 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X397 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X398 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X399 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X400 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X401 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X403 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X404 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X407 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X408 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X409 a_n8964_8799# plus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X410 a_n2650_13878# minus a_n2903_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X411 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X412 a_n2650_8322# a_n2650_13878# a_n8964_8799# vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X413 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X414 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 vdd a_n8964_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X416 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X417 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X418 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X419 a_n2650_8322# a_n2650_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X420 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X421 a_n2472_13878# a_n2650_13878# a_n2650_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X422 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X423 a_n2903_n3924# plus a_n8964_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X424 a_n2903_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X425 CSoutput a_n8964_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X426 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X427 a_n2650_13878# a_n2650_13878# a_n2472_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
.ends

