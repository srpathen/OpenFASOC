* NGSPICE file created from opamp683.ext - technology: sky130A

.subckt opamp683 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n9628_8799.t34 plus.t5 a_n2903_n3924.t31 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 CSoutput.t71 commonsourceibias.t48 gnd.t160 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n2804_13878.t7 a_n2982_13878.t64 vdd.t291 vdd.t290 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2804_13878.t31 a_n2982_13878.t17 a_n2982_13878.t18 vdd.t278 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 vdd.t159 a_n9628_8799.t40 CSoutput.t181 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 gnd.t72 commonsourceibias.t49 CSoutput.t70 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 CSoutput.t69 commonsourceibias.t50 gnd.t104 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t68 commonsourceibias.t51 gnd.t159 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 CSoutput.t180 a_n9628_8799.t41 vdd.t158 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 a_n2903_n3924.t32 plus.t6 a_n9628_8799.t33 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X10 plus.t0 gnd.t288 gnd.t290 gnd.t289 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X11 vdd.t157 a_n9628_8799.t42 CSoutput.t140 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 a_n2982_8322.t23 a_n2982_13878.t65 a_n9628_8799.t38 vdd.t288 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 CSoutput.t139 a_n9628_8799.t43 vdd.t156 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X14 vdd.t155 a_n9628_8799.t44 CSoutput.t138 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 output.t18 CSoutput.t192 vdd.t304 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X16 CSoutput.t137 a_n9628_8799.t45 vdd.t154 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X17 gnd.t161 commonsourceibias.t52 CSoutput.t67 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X18 vdd.t298 CSoutput.t193 output.t17 gnd.t67 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X19 CSoutput.t66 commonsourceibias.t53 gnd.t59 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 gnd.t82 commonsourceibias.t54 CSoutput.t65 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X21 vdd.t153 a_n9628_8799.t46 CSoutput.t150 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 vdd.t152 a_n9628_8799.t47 CSoutput.t149 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X23 CSoutput.t64 commonsourceibias.t55 gnd.t60 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 CSoutput.t63 commonsourceibias.t56 gnd.t83 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 CSoutput.t148 a_n9628_8799.t48 vdd.t151 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X26 CSoutput.t62 commonsourceibias.t57 gnd.t139 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 a_n9628_8799.t10 a_n2982_13878.t66 a_n2982_8322.t22 vdd.t274 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X28 vdd.t150 a_n9628_8799.t49 CSoutput.t147 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 a_n2982_13878.t6 minus.t5 a_n2903_n3924.t6 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X30 vdd.t149 a_n9628_8799.t50 CSoutput.t75 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 CSoutput.t74 a_n9628_8799.t51 vdd.t148 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 a_n9628_8799.t12 a_n2982_13878.t67 a_n2982_8322.t21 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 CSoutput.t61 commonsourceibias.t58 gnd.t110 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 gnd.t71 commonsourceibias.t59 CSoutput.t60 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t287 gnd.t285 gnd.t286 gnd.t211 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X36 CSoutput.t59 commonsourceibias.t60 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 a_n2903_n3924.t2 minus.t6 a_n2982_13878.t2 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X38 gnd.t284 gnd.t282 minus.t4 gnd.t283 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X39 CSoutput.t58 commonsourceibias.t61 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 vdd.t297 CSoutput.t194 output.t16 gnd.t68 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X41 CSoutput.t73 a_n9628_8799.t52 vdd.t147 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X42 a_n2903_n3924.t9 diffpairibias.t16 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 CSoutput.t72 a_n9628_8799.t53 vdd.t146 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 vdd.t145 a_n9628_8799.t54 CSoutput.t83 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 gnd.t96 commonsourceibias.t62 CSoutput.t57 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 gnd.t281 gnd.t279 gnd.t280 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X47 vdd.t144 a_n9628_8799.t55 CSoutput.t82 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 CSoutput.t56 commonsourceibias.t63 gnd.t129 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X49 output.t2 outputibias.t8 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X50 gnd.t50 commonsourceibias.t46 commonsourceibias.t47 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 CSoutput.t55 commonsourceibias.t64 gnd.t295 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 CSoutput.t195 a_n2982_8322.t37 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X53 vdd.t235 vdd.t233 vdd.t234 vdd.t224 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X54 a_n2903_n3924.t33 plus.t7 a_n9628_8799.t32 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X55 vdd.t143 a_n9628_8799.t56 CSoutput.t81 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X56 vdd.t306 CSoutput.t196 output.t15 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X57 a_n2804_13878.t30 a_n2982_13878.t45 a_n2982_13878.t46 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 CSoutput.t54 commonsourceibias.t65 gnd.t306 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 output.t14 CSoutput.t197 vdd.t299 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X60 a_n2982_13878.t36 a_n2982_13878.t35 a_n2804_13878.t29 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X61 vdd.t232 vdd.t230 vdd.t231 vdd.t224 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X62 gnd.t130 commonsourceibias.t66 CSoutput.t53 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 a_n9628_8799.t31 plus.t8 a_n2903_n3924.t21 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X64 CSoutput.t80 a_n9628_8799.t57 vdd.t142 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 gnd.t140 commonsourceibias.t44 commonsourceibias.t45 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 vdd.t229 vdd.t227 vdd.t228 vdd.t206 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X67 CSoutput.t52 commonsourceibias.t67 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 vdd.t141 a_n9628_8799.t58 CSoutput.t153 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X69 vdd.t140 a_n9628_8799.t59 CSoutput.t152 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 gnd.t278 gnd.t276 gnd.t277 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X71 gnd.t275 gnd.t272 gnd.t274 gnd.t273 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X72 gnd.t271 gnd.t269 gnd.t270 gnd.t211 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X73 CSoutput.t51 commonsourceibias.t68 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 diffpairibias.t15 diffpairibias.t14 gnd.t135 gnd.t134 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X75 CSoutput.t151 a_n9628_8799.t60 vdd.t138 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 a_n2982_13878.t61 minus.t7 a_n2903_n3924.t17 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X77 a_n2982_13878.t44 a_n2982_13878.t43 a_n2804_13878.t28 vdd.t273 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X78 CSoutput.t50 commonsourceibias.t69 gnd.t307 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X79 CSoutput.t79 a_n9628_8799.t61 vdd.t137 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 CSoutput.t49 commonsourceibias.t70 gnd.t133 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X81 gnd.t150 commonsourceibias.t71 CSoutput.t48 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 vdd.t136 a_n9628_8799.t62 CSoutput.t78 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 a_n9628_8799.t14 a_n2982_13878.t68 a_n2982_8322.t20 vdd.t268 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X84 CSoutput.t77 a_n9628_8799.t63 vdd.t135 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X85 gnd.t163 commonsourceibias.t72 CSoutput.t47 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 CSoutput.t198 a_n2982_8322.t36 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X87 a_n2982_13878.t50 a_n2982_13878.t49 a_n2804_13878.t27 vdd.t289 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X88 vdd.t134 a_n9628_8799.t64 CSoutput.t76 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 vdd.t133 a_n9628_8799.t65 CSoutput.t108 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 a_n9628_8799.t37 a_n2982_13878.t69 a_n2982_8322.t19 vdd.t266 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X91 CSoutput.t107 a_n9628_8799.t66 vdd.t132 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 CSoutput.t46 commonsourceibias.t73 gnd.t301 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X93 diffpairibias.t13 diffpairibias.t12 gnd.t90 gnd.t89 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X94 CSoutput.t106 a_n9628_8799.t67 vdd.t131 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 gnd.t42 commonsourceibias.t42 commonsourceibias.t43 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 a_n9628_8799.t9 a_n2982_13878.t70 a_n2982_8322.t18 vdd.t283 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X97 CSoutput.t45 commonsourceibias.t74 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 gnd.t297 commonsourceibias.t75 CSoutput.t44 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 CSoutput.t43 commonsourceibias.t76 gnd.t86 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 a_n2982_8322.t17 a_n2982_13878.t71 a_n9628_8799.t8 vdd.t289 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X101 gnd.t34 commonsourceibias.t77 CSoutput.t42 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 CSoutput.t105 a_n9628_8799.t68 vdd.t130 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 output.t13 CSoutput.t199 vdd.t293 gnd.t47 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X104 vdd.t294 CSoutput.t200 output.t12 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X105 vdd.t226 vdd.t223 vdd.t225 vdd.t224 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X106 a_n2903_n3924.t22 plus.t9 a_n9628_8799.t30 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X107 gnd.t268 gnd.t266 minus.t3 gnd.t267 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X108 gnd.t100 commonsourceibias.t78 CSoutput.t41 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 a_n2903_n3924.t8 diffpairibias.t17 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X110 CSoutput.t93 a_n9628_8799.t69 vdd.t129 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 vdd.t127 a_n9628_8799.t70 CSoutput.t92 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X112 gnd.t265 gnd.t263 gnd.t264 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X113 vdd.t126 a_n9628_8799.t71 CSoutput.t91 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 a_n2982_13878.t56 a_n2982_13878.t55 a_n2804_13878.t26 vdd.t288 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X115 vdd.t125 a_n9628_8799.t72 CSoutput.t87 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 gnd.t158 commonsourceibias.t79 CSoutput.t40 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 a_n9628_8799.t4 a_n2982_13878.t72 a_n2982_8322.t16 vdd.t277 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X118 a_n2982_13878.t42 a_n2982_13878.t41 a_n2804_13878.t25 vdd.t240 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X119 gnd.t262 gnd.t260 gnd.t261 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X120 vdd.t295 CSoutput.t201 output.t11 gnd.t298 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X121 vdd.t124 a_n9628_8799.t73 CSoutput.t86 vdd.t87 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X122 CSoutput.t85 a_n9628_8799.t74 vdd.t123 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 gnd.t164 commonsourceibias.t80 CSoutput.t39 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 CSoutput.t84 a_n9628_8799.t75 vdd.t122 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X125 a_n2982_13878.t4 minus.t8 a_n2903_n3924.t4 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X126 vdd.t222 vdd.t220 vdd.t221 vdd.t213 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X127 gnd.t319 commonsourceibias.t40 commonsourceibias.t41 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X128 output.t10 CSoutput.t202 vdd.t300 gnd.t299 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X129 gnd.t114 commonsourceibias.t81 CSoutput.t38 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 CSoutput.t171 a_n9628_8799.t76 vdd.t121 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 vdd.t219 vdd.t216 vdd.t218 vdd.t217 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X132 gnd.t259 gnd.t257 gnd.t258 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X133 a_n2804_13878.t24 a_n2982_13878.t57 a_n2982_13878.t58 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X134 a_n2903_n3924.t11 minus.t9 a_n2982_13878.t9 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X135 CSoutput.t170 a_n9628_8799.t77 vdd.t120 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X136 vdd.t119 a_n9628_8799.t78 CSoutput.t169 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X137 vdd.t282 a_n2982_13878.t73 a_n2982_8322.t31 vdd.t281 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X138 a_n2982_13878.t54 a_n2982_13878.t53 a_n2804_13878.t23 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X139 a_n2982_8322.t30 a_n2982_13878.t74 vdd.t287 vdd.t286 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X140 a_n2903_n3924.t39 diffpairibias.t18 gnd.t317 gnd.t316 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X141 CSoutput.t168 a_n9628_8799.t79 vdd.t118 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 output.t9 CSoutput.t203 vdd.t303 gnd.t300 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X143 CSoutput.t37 commonsourceibias.t82 gnd.t101 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X144 CSoutput.t36 commonsourceibias.t83 gnd.t136 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 gnd.t256 gnd.t254 gnd.t255 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X146 a_n2903_n3924.t10 minus.t10 a_n2982_13878.t8 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X147 gnd.t253 gnd.t251 plus.t3 gnd.t252 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X148 vdd.t285 a_n2982_13878.t75 a_n2804_13878.t6 vdd.t284 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X149 a_n2903_n3924.t19 plus.t10 a_n9628_8799.t29 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X150 vdd.t215 vdd.t212 vdd.t214 vdd.t213 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X151 gnd.t250 gnd.t248 gnd.t249 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X152 a_n2804_13878.t22 a_n2982_13878.t47 a_n2982_13878.t48 vdd.t283 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 vdd.t117 a_n9628_8799.t80 CSoutput.t131 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 vdd.t115 a_n9628_8799.t81 CSoutput.t130 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 a_n2982_8322.t15 a_n2982_13878.t76 a_n9628_8799.t7 vdd.t267 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 a_n9628_8799.t28 plus.t11 a_n2903_n3924.t23 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X157 a_n9628_8799.t27 plus.t12 a_n2903_n3924.t25 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X158 vdd.t211 vdd.t209 vdd.t210 vdd.t186 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X159 vdd.t208 vdd.t205 vdd.t207 vdd.t206 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X160 a_n2982_8322.t29 a_n2982_13878.t77 vdd.t280 vdd.t279 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X161 a_n9628_8799.t18 a_n2982_13878.t78 a_n2982_8322.t14 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 CSoutput.t129 a_n9628_8799.t82 vdd.t114 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X163 diffpairibias.t11 diffpairibias.t10 gnd.t116 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X164 vdd.t113 a_n9628_8799.t83 CSoutput.t183 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X165 a_n2982_13878.t63 minus.t11 a_n2903_n3924.t36 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X166 a_n2982_13878.t32 a_n2982_13878.t31 a_n2804_13878.t21 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X167 CSoutput.t35 commonsourceibias.t84 gnd.t91 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 a_n9628_8799.t39 a_n2982_13878.t79 a_n2982_8322.t13 vdd.t278 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X169 CSoutput.t182 a_n9628_8799.t84 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 CSoutput.t144 a_n9628_8799.t85 vdd.t109 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 commonsourceibias.t39 commonsourceibias.t38 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 gnd.t79 commonsourceibias.t85 CSoutput.t34 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 a_n2804_13878.t20 a_n2982_13878.t11 a_n2982_13878.t12 vdd.t277 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X174 gnd.t247 gnd.t244 gnd.t246 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X175 a_n2903_n3924.t5 minus.t12 a_n2982_13878.t5 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X176 minus.t2 gnd.t241 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X177 vdd.t204 vdd.t202 vdd.t203 vdd.t165 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X178 outputibias.t7 outputibias.t6 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X179 vdd.t302 CSoutput.t204 output.t8 gnd.t296 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X180 CSoutput.t143 a_n9628_8799.t86 vdd.t108 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X181 CSoutput.t33 commonsourceibias.t86 gnd.t128 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 vdd.t276 a_n2982_13878.t80 a_n2982_8322.t28 vdd.t275 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X183 a_n2804_13878.t19 a_n2982_13878.t51 a_n2982_13878.t52 vdd.t274 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X184 vdd.t107 a_n9628_8799.t87 CSoutput.t142 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 vdd.t106 a_n9628_8799.t88 CSoutput.t141 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X186 a_n2982_13878.t16 a_n2982_13878.t15 a_n2804_13878.t18 vdd.t244 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X187 gnd.t119 commonsourceibias.t87 CSoutput.t32 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 gnd.t113 commonsourceibias.t88 CSoutput.t31 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 commonsourceibias.t37 commonsourceibias.t36 gnd.t65 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 outputibias.t5 outputibias.t4 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X191 gnd.t122 commonsourceibias.t89 CSoutput.t30 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X192 vdd.t105 a_n9628_8799.t89 CSoutput.t162 vdd.t87 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X193 vdd.t104 a_n9628_8799.t90 CSoutput.t161 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X194 CSoutput.t29 commonsourceibias.t90 gnd.t131 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 CSoutput.t160 a_n9628_8799.t91 vdd.t103 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 a_n2903_n3924.t13 diffpairibias.t19 gnd.t106 gnd.t105 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X197 gnd.t240 gnd.t237 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X198 vdd.t201 vdd.t199 vdd.t200 vdd.t173 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X199 a_n2903_n3924.t12 diffpairibias.t20 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X200 commonsourceibias.t35 commonsourceibias.t34 gnd.t303 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 vdd.t102 a_n9628_8799.t92 CSoutput.t159 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 vdd.t101 a_n9628_8799.t93 CSoutput.t115 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 CSoutput.t114 a_n9628_8799.t94 vdd.t100 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X204 gnd.t236 gnd.t234 gnd.t235 gnd.t211 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X205 vdd.t198 vdd.t196 vdd.t197 vdd.t186 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X206 CSoutput.t28 commonsourceibias.t91 gnd.t97 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 CSoutput.t27 commonsourceibias.t92 gnd.t293 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 a_n2804_13878.t17 a_n2982_13878.t25 a_n2982_13878.t26 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 gnd.t233 gnd.t231 gnd.t232 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X210 a_n2982_8322.t12 a_n2982_13878.t81 a_n9628_8799.t6 vdd.t273 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X211 CSoutput.t113 a_n9628_8799.t95 vdd.t99 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X212 CSoutput.t112 a_n9628_8799.t96 vdd.t98 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 commonsourceibias.t33 commonsourceibias.t32 gnd.t147 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 CSoutput.t205 a_n2982_8322.t35 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X215 diffpairibias.t9 diffpairibias.t8 gnd.t311 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X216 a_n2804_13878.t5 a_n2982_13878.t82 vdd.t272 vdd.t271 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X217 vdd.t270 a_n2982_13878.t83 a_n2804_13878.t4 vdd.t269 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X218 CSoutput.t26 commonsourceibias.t93 gnd.t170 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 CSoutput.t25 commonsourceibias.t94 gnd.t292 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 CSoutput.t117 a_n9628_8799.t97 vdd.t97 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 CSoutput.t206 a_n2982_8322.t34 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X222 gnd.t18 commonsourceibias.t30 commonsourceibias.t31 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 vdd.t95 a_n9628_8799.t98 CSoutput.t116 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 vdd.t93 a_n9628_8799.t99 CSoutput.t173 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 gnd.t230 gnd.t227 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X226 gnd.t226 gnd.t224 plus.t2 gnd.t225 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X227 vdd.t91 a_n9628_8799.t100 CSoutput.t172 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 commonsourceibias.t29 commonsourceibias.t28 gnd.t53 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 CSoutput.t134 a_n9628_8799.t101 vdd.t89 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 a_n2804_13878.t16 a_n2982_13878.t13 a_n2982_13878.t14 vdd.t268 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X231 a_n2903_n3924.t14 minus.t13 a_n2982_13878.t10 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X232 gnd.t302 commonsourceibias.t95 CSoutput.t24 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X233 commonsourceibias.t27 commonsourceibias.t26 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X234 vdd.t88 a_n9628_8799.t102 CSoutput.t133 vdd.t87 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X235 vdd.t86 a_n9628_8799.t103 CSoutput.t132 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X236 output.t0 outputibias.t9 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X237 CSoutput.t125 a_n9628_8799.t104 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 gnd.t162 commonsourceibias.t24 commonsourceibias.t25 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 a_n2982_8322.t11 a_n2982_13878.t84 a_n9628_8799.t5 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X240 a_n2982_13878.t38 a_n2982_13878.t37 a_n2804_13878.t15 vdd.t267 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X241 CSoutput.t124 a_n9628_8799.t105 vdd.t83 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X242 diffpairibias.t7 diffpairibias.t6 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X243 gnd.t223 gnd.t221 gnd.t222 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X244 vdd.t82 a_n9628_8799.t106 CSoutput.t123 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X245 a_n2804_13878.t14 a_n2982_13878.t23 a_n2982_13878.t24 vdd.t266 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X246 commonsourceibias.t23 commonsourceibias.t22 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X247 a_n2982_13878.t0 minus.t14 a_n2903_n3924.t0 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X248 a_n2982_13878.t59 minus.t15 a_n2903_n3924.t15 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X249 vdd.t265 a_n2982_13878.t85 a_n2982_8322.t27 vdd.t264 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X250 vdd.t292 CSoutput.t207 output.t7 gnd.t152 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X251 vdd.t80 a_n9628_8799.t107 CSoutput.t119 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 a_n9628_8799.t26 plus.t13 a_n2903_n3924.t30 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X253 gnd.t14 commonsourceibias.t96 CSoutput.t23 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 a_n2903_n3924.t16 minus.t16 a_n2982_13878.t60 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X255 CSoutput.t118 a_n9628_8799.t108 vdd.t78 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 gnd.t98 commonsourceibias.t20 commonsourceibias.t21 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 a_n2804_13878.t3 a_n2982_13878.t86 vdd.t263 vdd.t262 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X258 vdd.t77 a_n9628_8799.t109 CSoutput.t185 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X259 CSoutput.t184 a_n9628_8799.t110 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X260 CSoutput.t157 a_n9628_8799.t111 vdd.t73 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 gnd.t220 gnd.t217 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X262 vdd.t195 vdd.t193 vdd.t194 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X263 vdd.t72 a_n9628_8799.t112 CSoutput.t156 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X264 a_n2903_n3924.t35 diffpairibias.t21 gnd.t305 gnd.t304 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X265 vdd.t261 a_n2982_13878.t87 a_n2982_8322.t26 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X266 a_n2982_8322.t10 a_n2982_13878.t88 a_n9628_8799.t13 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X267 gnd.t99 commonsourceibias.t18 commonsourceibias.t19 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 vdd.t71 a_n9628_8799.t113 CSoutput.t155 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 a_n9628_8799.t25 plus.t14 a_n2903_n3924.t34 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X270 gnd.t216 gnd.t214 plus.t4 gnd.t215 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X271 gnd.t294 commonsourceibias.t16 commonsourceibias.t17 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 vdd.t192 vdd.t189 vdd.t191 vdd.t190 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X273 vdd.t70 a_n9628_8799.t114 CSoutput.t154 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 a_n2903_n3924.t29 plus.t15 a_n9628_8799.t24 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X275 vdd.t69 a_n9628_8799.t115 CSoutput.t111 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 output.t6 CSoutput.t208 vdd.t301 gnd.t153 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X277 vdd.t68 a_n9628_8799.t116 CSoutput.t110 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X278 CSoutput.t109 a_n9628_8799.t117 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 CSoutput.t96 a_n9628_8799.t118 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X280 CSoutput.t22 commonsourceibias.t97 gnd.t107 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 a_n2804_13878.t13 a_n2982_13878.t27 a_n2982_13878.t28 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X282 CSoutput.t95 a_n9628_8799.t119 vdd.t63 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 CSoutput.t94 a_n9628_8799.t120 vdd.t62 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X284 a_n2982_8322.t9 a_n2982_13878.t89 a_n9628_8799.t2 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X285 diffpairibias.t5 diffpairibias.t4 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X286 gnd.t213 gnd.t210 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X287 CSoutput.t90 a_n9628_8799.t121 vdd.t61 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 CSoutput.t89 a_n9628_8799.t122 vdd.t59 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 vdd.t188 vdd.t185 vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X290 CSoutput.t21 commonsourceibias.t98 gnd.t22 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X291 vdd.t58 a_n9628_8799.t123 CSoutput.t88 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 CSoutput.t209 a_n2982_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X293 a_n2982_8322.t25 a_n2982_13878.t90 vdd.t257 vdd.t256 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X294 CSoutput.t176 a_n9628_8799.t124 vdd.t57 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 outputibias.t3 outputibias.t2 gnd.t121 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X296 gnd.t209 gnd.t206 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X297 vdd.t55 a_n9628_8799.t125 CSoutput.t175 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 gnd.t205 gnd.t203 gnd.t204 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X299 gnd.t24 commonsourceibias.t99 CSoutput.t20 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 CSoutput.t174 a_n9628_8799.t126 vdd.t54 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 output.t1 outputibias.t10 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X302 vdd.t255 a_n2982_13878.t91 a_n2804_13878.t2 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X303 vdd.t53 a_n9628_8799.t127 CSoutput.t136 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 CSoutput.t135 a_n9628_8799.t128 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 vdd.t49 a_n9628_8799.t129 CSoutput.t128 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 gnd.t80 commonsourceibias.t100 CSoutput.t19 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 output.t19 outputibias.t11 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X308 gnd.t52 commonsourceibias.t101 CSoutput.t18 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 gnd.t177 gnd.t174 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X310 a_n2982_8322.t8 a_n2982_13878.t92 a_n9628_8799.t0 vdd.t246 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X311 commonsourceibias.t15 commonsourceibias.t14 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 gnd.t202 gnd.t200 minus.t1 gnd.t201 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X313 a_n9628_8799.t15 a_n2982_13878.t93 a_n2982_8322.t7 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X314 a_n2804_13878.t1 a_n2982_13878.t94 vdd.t252 vdd.t251 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X315 gnd.t26 commonsourceibias.t102 CSoutput.t17 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 vdd.t47 a_n9628_8799.t130 CSoutput.t127 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 vdd.t184 vdd.t182 vdd.t183 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X318 vdd.t181 vdd.t179 vdd.t180 vdd.t173 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X319 vdd.t46 a_n9628_8799.t131 CSoutput.t126 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 a_n2982_13878.t1 minus.t17 a_n2903_n3924.t1 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X321 CSoutput.t104 a_n9628_8799.t132 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 CSoutput.t103 a_n9628_8799.t133 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X323 CSoutput.t187 a_n9628_8799.t134 vdd.t41 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 a_n2982_13878.t30 a_n2982_13878.t29 a_n2804_13878.t12 vdd.t241 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X325 a_n9628_8799.t1 a_n2982_13878.t95 a_n2982_8322.t6 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X326 minus.t0 gnd.t197 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X327 a_n9628_8799.t36 a_n2982_13878.t96 a_n2982_8322.t5 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X328 gnd.t108 commonsourceibias.t103 CSoutput.t16 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 commonsourceibias.t13 commonsourceibias.t12 gnd.t84 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 a_n9628_8799.t23 plus.t16 a_n2903_n3924.t28 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X331 a_n2982_8322.t4 a_n2982_13878.t97 a_n9628_8799.t11 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X332 gnd.t123 commonsourceibias.t104 CSoutput.t15 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 a_n2903_n3924.t7 minus.t18 a_n2982_13878.t7 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X334 vdd.t40 a_n9628_8799.t135 CSoutput.t186 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 gnd.t3 commonsourceibias.t10 commonsourceibias.t11 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 CSoutput.t178 a_n9628_8799.t136 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 CSoutput.t177 a_n9628_8799.t137 vdd.t36 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X338 CSoutput.t164 a_n9628_8799.t138 vdd.t35 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 CSoutput.t163 a_n9628_8799.t139 vdd.t34 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 a_n2804_13878.t11 a_n2982_13878.t21 a_n2982_13878.t22 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X341 vdd.t33 a_n9628_8799.t140 CSoutput.t100 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 vdd.t31 a_n9628_8799.t141 CSoutput.t121 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 a_n2903_n3924.t20 plus.t17 a_n9628_8799.t22 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X344 vdd.t30 a_n9628_8799.t142 CSoutput.t97 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X345 gnd.t157 commonsourceibias.t8 commonsourceibias.t9 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X346 commonsourceibias.t7 commonsourceibias.t6 gnd.t49 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 gnd.t166 commonsourceibias.t105 CSoutput.t14 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X348 a_n2903_n3924.t37 diffpairibias.t22 gnd.t309 gnd.t308 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X349 CSoutput.t13 commonsourceibias.t106 gnd.t27 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 output.t5 CSoutput.t210 vdd.t307 gnd.t154 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X351 vdd.t29 a_n9628_8799.t143 CSoutput.t120 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 gnd.t168 commonsourceibias.t107 CSoutput.t12 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 CSoutput.t165 a_n9628_8799.t144 vdd.t28 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 a_n2982_13878.t20 a_n2982_13878.t19 a_n2804_13878.t10 vdd.t246 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X355 gnd.t196 gnd.t193 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X356 a_n9628_8799.t16 a_n2982_13878.t98 a_n2982_8322.t3 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X357 gnd.t192 gnd.t190 gnd.t191 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X358 vdd.t27 a_n9628_8799.t145 CSoutput.t102 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 CSoutput.t211 a_n2982_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X360 CSoutput.t189 a_n9628_8799.t146 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 a_n9628_8799.t21 plus.t18 a_n2903_n3924.t26 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X362 vdd.t178 vdd.t176 vdd.t177 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X363 CSoutput.t11 commonsourceibias.t108 gnd.t167 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 gnd.t124 commonsourceibias.t109 CSoutput.t10 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X365 commonsourceibias.t5 commonsourceibias.t4 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 diffpairibias.t3 diffpairibias.t2 gnd.t118 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X367 gnd.t189 gnd.t186 gnd.t188 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X368 CSoutput.t101 a_n9628_8799.t147 vdd.t24 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X369 outputibias.t1 outputibias.t0 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X370 a_n2982_8322.t2 a_n2982_13878.t99 a_n9628_8799.t35 vdd.t244 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X371 gnd.t165 commonsourceibias.t110 CSoutput.t9 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X372 a_n2903_n3924.t24 plus.t19 a_n9628_8799.t20 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X373 vdd.t23 a_n9628_8799.t148 CSoutput.t179 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 vdd.t175 vdd.t172 vdd.t174 vdd.t173 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X375 gnd.t185 gnd.t182 gnd.t184 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X376 CSoutput.t190 a_n9628_8799.t149 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X377 CSoutput.t188 a_n9628_8799.t150 vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 diffpairibias.t1 diffpairibias.t0 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X379 commonsourceibias.t3 commonsourceibias.t2 gnd.t85 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 gnd.t127 commonsourceibias.t111 CSoutput.t8 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X381 a_n2903_n3924.t27 plus.t20 a_n9628_8799.t19 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X382 CSoutput.t7 commonsourceibias.t112 gnd.t146 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X383 vdd.t243 a_n2982_13878.t100 a_n2804_13878.t0 vdd.t242 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X384 CSoutput.t166 a_n9628_8799.t151 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X385 CSoutput.t122 a_n9628_8799.t152 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X386 a_n2903_n3924.t18 minus.t19 a_n2982_13878.t62 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X387 vdd.t13 a_n9628_8799.t153 CSoutput.t158 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 vdd.t11 a_n9628_8799.t154 CSoutput.t145 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X389 gnd.t94 commonsourceibias.t0 commonsourceibias.t1 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 vdd.t305 CSoutput.t212 output.t4 gnd.t155 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X391 a_n2982_8322.t1 a_n2982_13878.t101 a_n9628_8799.t3 vdd.t241 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X392 a_n2982_13878.t3 minus.t20 a_n2903_n3924.t3 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X393 output.t3 CSoutput.t213 vdd.t296 gnd.t156 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X394 gnd.t148 commonsourceibias.t113 CSoutput.t6 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X395 gnd.t57 commonsourceibias.t114 CSoutput.t5 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 gnd.t181 gnd.t178 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X397 a_n2982_8322.t0 a_n2982_13878.t102 a_n9628_8799.t17 vdd.t240 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X398 vdd.t9 a_n9628_8799.t155 CSoutput.t167 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X399 vdd.t7 a_n9628_8799.t156 CSoutput.t146 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X400 CSoutput.t191 a_n9628_8799.t157 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X401 gnd.t132 commonsourceibias.t115 CSoutput.t4 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 plus.t1 gnd.t171 gnd.t173 gnd.t172 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X403 vdd.t171 vdd.t168 vdd.t170 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X404 a_n2982_8322.t24 a_n2982_13878.t103 vdd.t239 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X405 gnd.t145 commonsourceibias.t116 CSoutput.t3 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 a_n2804_13878.t9 a_n2982_13878.t33 a_n2982_13878.t34 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X407 gnd.t318 commonsourceibias.t117 CSoutput.t2 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X408 CSoutput.t1 commonsourceibias.t118 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 CSoutput.t0 commonsourceibias.t119 gnd.t169 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X410 vdd.t167 vdd.t164 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X411 a_n2903_n3924.t38 diffpairibias.t23 gnd.t315 gnd.t314 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X412 vdd.t163 vdd.t160 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X413 vdd.t3 a_n9628_8799.t158 CSoutput.t99 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X414 CSoutput.t98 a_n9628_8799.t159 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 a_n2982_13878.t40 a_n2982_13878.t39 a_n2804_13878.t8 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 plus.n33 plus.t15 321.495
R1 plus.n7 plus.t12 321.495
R2 plus.n32 plus.t14 297.12
R3 plus.n36 plus.t19 297.12
R4 plus.n38 plus.t18 297.12
R5 plus.n42 plus.t20 297.12
R6 plus.n44 plus.t8 297.12
R7 plus.n48 plus.t7 297.12
R8 plus.n50 plus.t11 297.12
R9 plus.n24 plus.t9 297.12
R10 plus.n22 plus.t5 297.12
R11 plus.n2 plus.t6 297.12
R12 plus.n16 plus.t16 297.12
R13 plus.n4 plus.t17 297.12
R14 plus.n10 plus.t13 297.12
R15 plus.n6 plus.t10 297.12
R16 plus.n54 plus.t3 243.97
R17 plus.n54 plus.n53 223.454
R18 plus.n56 plus.n55 223.454
R19 plus.n51 plus.n50 161.3
R20 plus.n49 plus.n26 161.3
R21 plus.n48 plus.n47 161.3
R22 plus.n46 plus.n27 161.3
R23 plus.n45 plus.n44 161.3
R24 plus.n43 plus.n28 161.3
R25 plus.n42 plus.n41 161.3
R26 plus.n40 plus.n29 161.3
R27 plus.n39 plus.n38 161.3
R28 plus.n37 plus.n30 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n34 plus.n31 161.3
R31 plus.n9 plus.n8 161.3
R32 plus.n10 plus.n5 161.3
R33 plus.n12 plus.n11 161.3
R34 plus.n13 plus.n4 161.3
R35 plus.n15 plus.n14 161.3
R36 plus.n16 plus.n3 161.3
R37 plus.n18 plus.n17 161.3
R38 plus.n19 plus.n2 161.3
R39 plus.n21 plus.n20 161.3
R40 plus.n22 plus.n1 161.3
R41 plus.n23 plus.n0 161.3
R42 plus.n25 plus.n24 161.3
R43 plus.n34 plus.n33 44.9377
R44 plus.n8 plus.n7 44.9377
R45 plus.n50 plus.n49 37.246
R46 plus.n24 plus.n23 37.246
R47 plus.n32 plus.n31 32.8641
R48 plus.n48 plus.n27 32.8641
R49 plus.n22 plus.n21 32.8641
R50 plus.n9 plus.n6 32.8641
R51 plus.n52 plus.n51 30.0327
R52 plus.n37 plus.n36 28.4823
R53 plus.n44 plus.n43 28.4823
R54 plus.n17 plus.n2 28.4823
R55 plus.n11 plus.n10 28.4823
R56 plus.n38 plus.n29 24.1005
R57 plus.n42 plus.n29 24.1005
R58 plus.n16 plus.n15 24.1005
R59 plus.n15 plus.n4 24.1005
R60 plus.n53 plus.t2 19.8005
R61 plus.n53 plus.t0 19.8005
R62 plus.n55 plus.t4 19.8005
R63 plus.n55 plus.t1 19.8005
R64 plus.n38 plus.n37 19.7187
R65 plus.n43 plus.n42 19.7187
R66 plus.n17 plus.n16 19.7187
R67 plus.n11 plus.n4 19.7187
R68 plus.n33 plus.n32 17.0522
R69 plus.n7 plus.n6 17.0522
R70 plus.n36 plus.n31 15.3369
R71 plus.n44 plus.n27 15.3369
R72 plus.n21 plus.n2 15.3369
R73 plus.n10 plus.n9 15.3369
R74 plus plus.n57 14.3956
R75 plus.n52 plus.n25 11.8547
R76 plus.n49 plus.n48 10.955
R77 plus.n23 plus.n22 10.955
R78 plus.n57 plus.n56 5.40567
R79 plus.n57 plus.n52 1.188
R80 plus.n56 plus.n54 0.716017
R81 plus.n35 plus.n34 0.189894
R82 plus.n35 plus.n30 0.189894
R83 plus.n39 plus.n30 0.189894
R84 plus.n40 plus.n39 0.189894
R85 plus.n41 plus.n40 0.189894
R86 plus.n41 plus.n28 0.189894
R87 plus.n45 plus.n28 0.189894
R88 plus.n46 plus.n45 0.189894
R89 plus.n47 plus.n46 0.189894
R90 plus.n47 plus.n26 0.189894
R91 plus.n51 plus.n26 0.189894
R92 plus.n25 plus.n0 0.189894
R93 plus.n1 plus.n0 0.189894
R94 plus.n20 plus.n1 0.189894
R95 plus.n20 plus.n19 0.189894
R96 plus.n19 plus.n18 0.189894
R97 plus.n18 plus.n3 0.189894
R98 plus.n14 plus.n3 0.189894
R99 plus.n14 plus.n13 0.189894
R100 plus.n13 plus.n12 0.189894
R101 plus.n12 plus.n5 0.189894
R102 plus.n8 plus.n5 0.189894
R103 a_n2903_n3924.n6 a_n2903_n3924.t35 214.994
R104 a_n2903_n3924.n9 a_n2903_n3924.t39 214.714
R105 a_n2903_n3924.n9 a_n2903_n3924.t37 214.321
R106 a_n2903_n3924.n5 a_n2903_n3924.t12 214.321
R107 a_n2903_n3924.n5 a_n2903_n3924.t38 214.321
R108 a_n2903_n3924.n4 a_n2903_n3924.t13 214.321
R109 a_n2903_n3924.n6 a_n2903_n3924.t9 214.321
R110 a_n2903_n3924.n6 a_n2903_n3924.t8 214.321
R111 a_n2903_n3924.n3 a_n2903_n3924.t29 55.8337
R112 a_n2903_n3924.n3 a_n2903_n3924.t3 55.8337
R113 a_n2903_n3924.n7 a_n2903_n3924.t7 55.8337
R114 a_n2903_n3924.n1 a_n2903_n3924.t23 55.8335
R115 a_n2903_n3924.n0 a_n2903_n3924.t1 55.8335
R116 a_n2903_n3924.n2 a_n2903_n3924.t2 55.8335
R117 a_n2903_n3924.n2 a_n2903_n3924.t25 55.8335
R118 a_n2903_n3924.n8 a_n2903_n3924.t22 55.8335
R119 a_n2903_n3924.n23 a_n2903_n3924.n0 53.0054
R120 a_n2903_n3924.n1 a_n2903_n3924.n11 53.0052
R121 a_n2903_n3924.n1 a_n2903_n3924.n12 53.0052
R122 a_n2903_n3924.n1 a_n2903_n3924.n13 53.0052
R123 a_n2903_n3924.n3 a_n2903_n3924.n14 53.0052
R124 a_n2903_n3924.n3 a_n2903_n3924.n15 53.0052
R125 a_n2903_n3924.n7 a_n2903_n3924.n16 53.0052
R126 a_n2903_n3924.n0 a_n2903_n3924.n10 53.0051
R127 a_n2903_n3924.n0 a_n2903_n3924.n17 53.0051
R128 a_n2903_n3924.n2 a_n2903_n3924.n18 53.0051
R129 a_n2903_n3924.n2 a_n2903_n3924.n19 53.0051
R130 a_n2903_n3924.n8 a_n2903_n3924.n20 53.0051
R131 a_n2903_n3924.n21 a_n2903_n3924.n7 12.1986
R132 a_n2903_n3924.n22 a_n2903_n3924.n1 12.1986
R133 a_n2903_n3924.n21 a_n2903_n3924.n8 5.11903
R134 a_n2903_n3924.n0 a_n2903_n3924.n22 5.11903
R135 a_n2903_n3924.n10 a_n2903_n3924.t4 2.82907
R136 a_n2903_n3924.n10 a_n2903_n3924.t10 2.82907
R137 a_n2903_n3924.n17 a_n2903_n3924.t6 2.82907
R138 a_n2903_n3924.n17 a_n2903_n3924.t11 2.82907
R139 a_n2903_n3924.n18 a_n2903_n3924.t30 2.82907
R140 a_n2903_n3924.n18 a_n2903_n3924.t19 2.82907
R141 a_n2903_n3924.n19 a_n2903_n3924.t28 2.82907
R142 a_n2903_n3924.n19 a_n2903_n3924.t20 2.82907
R143 a_n2903_n3924.n20 a_n2903_n3924.t31 2.82907
R144 a_n2903_n3924.n20 a_n2903_n3924.t32 2.82907
R145 a_n2903_n3924.n11 a_n2903_n3924.t21 2.82907
R146 a_n2903_n3924.n11 a_n2903_n3924.t33 2.82907
R147 a_n2903_n3924.n12 a_n2903_n3924.t26 2.82907
R148 a_n2903_n3924.n12 a_n2903_n3924.t27 2.82907
R149 a_n2903_n3924.n13 a_n2903_n3924.t34 2.82907
R150 a_n2903_n3924.n13 a_n2903_n3924.t24 2.82907
R151 a_n2903_n3924.n14 a_n2903_n3924.t17 2.82907
R152 a_n2903_n3924.n14 a_n2903_n3924.t18 2.82907
R153 a_n2903_n3924.n15 a_n2903_n3924.t36 2.82907
R154 a_n2903_n3924.n15 a_n2903_n3924.t5 2.82907
R155 a_n2903_n3924.n16 a_n2903_n3924.t15 2.82907
R156 a_n2903_n3924.n16 a_n2903_n3924.t16 2.82907
R157 a_n2903_n3924.t0 a_n2903_n3924.n23 2.82907
R158 a_n2903_n3924.n23 a_n2903_n3924.t14 2.82907
R159 a_n2903_n3924.n3 a_n2903_n3924.n1 2.45524
R160 a_n2903_n3924.n2 a_n2903_n3924.n0 2.45524
R161 a_n2903_n3924.n6 a_n2903_n3924.n21 1.95694
R162 a_n2903_n3924.n22 a_n2903_n3924.n9 1.95694
R163 a_n2903_n3924.n5 a_n2903_n3924.n4 1.34352
R164 a_n2903_n3924.n4 a_n2903_n3924.n6 1.34352
R165 a_n2903_n3924.n8 a_n2903_n3924.n2 1.3324
R166 a_n2903_n3924.n7 a_n2903_n3924.n3 1.3324
R167 a_n2903_n3924.n9 a_n2903_n3924.n5 0.951808
R168 a_n9628_8799.n228 a_n9628_8799.t137 485.149
R169 a_n9628_8799.n290 a_n9628_8799.t152 485.149
R170 a_n9628_8799.n353 a_n9628_8799.t75 485.149
R171 a_n9628_8799.n38 a_n9628_8799.t89 485.149
R172 a_n9628_8799.n100 a_n9628_8799.t102 485.149
R173 a_n9628_8799.n163 a_n9628_8799.t73 485.149
R174 a_n9628_8799.n271 a_n9628_8799.t47 464.166
R175 a_n9628_8799.n270 a_n9628_8799.t45 464.166
R176 a_n9628_8799.n212 a_n9628_8799.t131 464.166
R177 a_n9628_8799.n264 a_n9628_8799.t67 464.166
R178 a_n9628_8799.n263 a_n9628_8799.t50 464.166
R179 a_n9628_8799.n215 a_n9628_8799.t138 464.166
R180 a_n9628_8799.n257 a_n9628_8799.t93 464.166
R181 a_n9628_8799.n256 a_n9628_8799.t68 464.166
R182 a_n9628_8799.n218 a_n9628_8799.t156 464.166
R183 a_n9628_8799.n250 a_n9628_8799.t111 464.166
R184 a_n9628_8799.n249 a_n9628_8799.t71 464.166
R185 a_n9628_8799.n221 a_n9628_8799.t150 464.166
R186 a_n9628_8799.n243 a_n9628_8799.t113 464.166
R187 a_n9628_8799.n242 a_n9628_8799.t85 464.166
R188 a_n9628_8799.n224 a_n9628_8799.t46 464.166
R189 a_n9628_8799.n236 a_n9628_8799.t134 464.166
R190 a_n9628_8799.n235 a_n9628_8799.t115 464.166
R191 a_n9628_8799.n227 a_n9628_8799.t51 464.166
R192 a_n9628_8799.n229 a_n9628_8799.t141 464.166
R193 a_n9628_8799.n333 a_n9628_8799.t58 464.166
R194 a_n9628_8799.n332 a_n9628_8799.t57 464.166
R195 a_n9628_8799.n274 a_n9628_8799.t148 464.166
R196 a_n9628_8799.n326 a_n9628_8799.t76 464.166
R197 a_n9628_8799.n325 a_n9628_8799.t65 464.166
R198 a_n9628_8799.n277 a_n9628_8799.t151 464.166
R199 a_n9628_8799.n319 a_n9628_8799.t107 464.166
R200 a_n9628_8799.n318 a_n9628_8799.t79 464.166
R201 a_n9628_8799.n280 a_n9628_8799.t49 464.166
R202 a_n9628_8799.n312 a_n9628_8799.t124 464.166
R203 a_n9628_8799.n311 a_n9628_8799.t80 464.166
R204 a_n9628_8799.n283 a_n9628_8799.t41 464.166
R205 a_n9628_8799.n305 a_n9628_8799.t129 464.166
R206 a_n9628_8799.n304 a_n9628_8799.t95 464.166
R207 a_n9628_8799.n286 a_n9628_8799.t59 464.166
R208 a_n9628_8799.n298 a_n9628_8799.t149 464.166
R209 a_n9628_8799.n297 a_n9628_8799.t130 464.166
R210 a_n9628_8799.n289 a_n9628_8799.t66 464.166
R211 a_n9628_8799.n291 a_n9628_8799.t153 464.166
R212 a_n9628_8799.n396 a_n9628_8799.t106 464.166
R213 a_n9628_8799.n395 a_n9628_8799.t128 464.166
R214 a_n9628_8799.n337 a_n9628_8799.t64 464.166
R215 a_n9628_8799.n389 a_n9628_8799.t146 464.166
R216 a_n9628_8799.n388 a_n9628_8799.t83 464.166
R217 a_n9628_8799.n340 a_n9628_8799.t139 464.166
R218 a_n9628_8799.n382 a_n9628_8799.t70 464.166
R219 a_n9628_8799.n381 a_n9628_8799.t118 464.166
R220 a_n9628_8799.n343 a_n9628_8799.t55 464.166
R221 a_n9628_8799.n375 a_n9628_8799.t101 464.166
R222 a_n9628_8799.n374 a_n9628_8799.t78 464.166
R223 a_n9628_8799.n346 a_n9628_8799.t126 464.166
R224 a_n9628_8799.n368 a_n9628_8799.t62 464.166
R225 a_n9628_8799.n367 a_n9628_8799.t110 464.166
R226 a_n9628_8799.n349 a_n9628_8799.t44 464.166
R227 a_n9628_8799.n361 a_n9628_8799.t94 464.166
R228 a_n9628_8799.n360 a_n9628_8799.t158 464.166
R229 a_n9628_8799.n352 a_n9628_8799.t117 464.166
R230 a_n9628_8799.n354 a_n9628_8799.t54 464.166
R231 a_n9628_8799.n39 a_n9628_8799.t91 464.166
R232 a_n9628_8799.n41 a_n9628_8799.t123 464.166
R233 a_n9628_8799.n45 a_n9628_8799.t48 464.166
R234 a_n9628_8799.n46 a_n9628_8799.t87 464.166
R235 a_n9628_8799.n34 a_n9628_8799.t119 464.166
R236 a_n9628_8799.n52 a_n9628_8799.t42 464.166
R237 a_n9628_8799.n53 a_n9628_8799.t74 464.166
R238 a_n9628_8799.n57 a_n9628_8799.t112 464.166
R239 a_n9628_8799.n59 a_n9628_8799.t147 464.166
R240 a_n9628_8799.n30 a_n9628_8799.t72 464.166
R241 a_n9628_8799.n64 a_n9628_8799.t108 464.166
R242 a_n9628_8799.n28 a_n9628_8799.t143 464.166
R243 a_n9628_8799.n69 a_n9628_8799.t144 464.166
R244 a_n9628_8799.n71 a_n9628_8799.t90 464.166
R245 a_n9628_8799.n75 a_n9628_8799.t122 464.166
R246 a_n9628_8799.n76 a_n9628_8799.t142 464.166
R247 a_n9628_8799.n24 a_n9628_8799.t86 464.166
R248 a_n9628_8799.n82 a_n9628_8799.t88 464.166
R249 a_n9628_8799.n83 a_n9628_8799.t120 464.166
R250 a_n9628_8799.n101 a_n9628_8799.t104 464.166
R251 a_n9628_8799.n103 a_n9628_8799.t140 464.166
R252 a_n9628_8799.n107 a_n9628_8799.t60 464.166
R253 a_n9628_8799.n108 a_n9628_8799.t98 464.166
R254 a_n9628_8799.n96 a_n9628_8799.t132 464.166
R255 a_n9628_8799.n114 a_n9628_8799.t56 464.166
R256 a_n9628_8799.n115 a_n9628_8799.t84 464.166
R257 a_n9628_8799.n119 a_n9628_8799.t125 464.166
R258 a_n9628_8799.n121 a_n9628_8799.t159 464.166
R259 a_n9628_8799.n92 a_n9628_8799.t81 464.166
R260 a_n9628_8799.n126 a_n9628_8799.t121 464.166
R261 a_n9628_8799.n90 a_n9628_8799.t155 464.166
R262 a_n9628_8799.n131 a_n9628_8799.t157 464.166
R263 a_n9628_8799.n133 a_n9628_8799.t103 464.166
R264 a_n9628_8799.n137 a_n9628_8799.t136 464.166
R265 a_n9628_8799.n138 a_n9628_8799.t154 464.166
R266 a_n9628_8799.n86 a_n9628_8799.t97 464.166
R267 a_n9628_8799.n144 a_n9628_8799.t99 464.166
R268 a_n9628_8799.n145 a_n9628_8799.t133 464.166
R269 a_n9628_8799.n164 a_n9628_8799.t52 464.166
R270 a_n9628_8799.n166 a_n9628_8799.t114 464.166
R271 a_n9628_8799.n170 a_n9628_8799.t69 464.166
R272 a_n9628_8799.n171 a_n9628_8799.t92 464.166
R273 a_n9628_8799.n159 a_n9628_8799.t43 464.166
R274 a_n9628_8799.n177 a_n9628_8799.t109 464.166
R275 a_n9628_8799.n178 a_n9628_8799.t61 464.166
R276 a_n9628_8799.n182 a_n9628_8799.t127 464.166
R277 a_n9628_8799.n184 a_n9628_8799.t77 464.166
R278 a_n9628_8799.n155 a_n9628_8799.t100 464.166
R279 a_n9628_8799.n189 a_n9628_8799.t53 464.166
R280 a_n9628_8799.n153 a_n9628_8799.t116 464.166
R281 a_n9628_8799.n194 a_n9628_8799.t96 464.166
R282 a_n9628_8799.n196 a_n9628_8799.t135 464.166
R283 a_n9628_8799.n200 a_n9628_8799.t82 464.166
R284 a_n9628_8799.n201 a_n9628_8799.t145 464.166
R285 a_n9628_8799.n149 a_n9628_8799.t63 464.166
R286 a_n9628_8799.n207 a_n9628_8799.t40 464.166
R287 a_n9628_8799.n208 a_n9628_8799.t105 464.166
R288 a_n9628_8799.n231 a_n9628_8799.n230 161.3
R289 a_n9628_8799.n232 a_n9628_8799.n227 161.3
R290 a_n9628_8799.n234 a_n9628_8799.n233 161.3
R291 a_n9628_8799.n235 a_n9628_8799.n226 161.3
R292 a_n9628_8799.n236 a_n9628_8799.n225 161.3
R293 a_n9628_8799.n238 a_n9628_8799.n237 161.3
R294 a_n9628_8799.n239 a_n9628_8799.n224 161.3
R295 a_n9628_8799.n241 a_n9628_8799.n240 161.3
R296 a_n9628_8799.n242 a_n9628_8799.n223 161.3
R297 a_n9628_8799.n243 a_n9628_8799.n222 161.3
R298 a_n9628_8799.n245 a_n9628_8799.n244 161.3
R299 a_n9628_8799.n246 a_n9628_8799.n221 161.3
R300 a_n9628_8799.n248 a_n9628_8799.n247 161.3
R301 a_n9628_8799.n249 a_n9628_8799.n220 161.3
R302 a_n9628_8799.n250 a_n9628_8799.n219 161.3
R303 a_n9628_8799.n252 a_n9628_8799.n251 161.3
R304 a_n9628_8799.n253 a_n9628_8799.n218 161.3
R305 a_n9628_8799.n255 a_n9628_8799.n254 161.3
R306 a_n9628_8799.n256 a_n9628_8799.n217 161.3
R307 a_n9628_8799.n257 a_n9628_8799.n216 161.3
R308 a_n9628_8799.n259 a_n9628_8799.n258 161.3
R309 a_n9628_8799.n260 a_n9628_8799.n215 161.3
R310 a_n9628_8799.n262 a_n9628_8799.n261 161.3
R311 a_n9628_8799.n263 a_n9628_8799.n214 161.3
R312 a_n9628_8799.n264 a_n9628_8799.n213 161.3
R313 a_n9628_8799.n266 a_n9628_8799.n265 161.3
R314 a_n9628_8799.n267 a_n9628_8799.n212 161.3
R315 a_n9628_8799.n269 a_n9628_8799.n268 161.3
R316 a_n9628_8799.n270 a_n9628_8799.n211 161.3
R317 a_n9628_8799.n272 a_n9628_8799.n271 161.3
R318 a_n9628_8799.n293 a_n9628_8799.n292 161.3
R319 a_n9628_8799.n294 a_n9628_8799.n289 161.3
R320 a_n9628_8799.n296 a_n9628_8799.n295 161.3
R321 a_n9628_8799.n297 a_n9628_8799.n288 161.3
R322 a_n9628_8799.n298 a_n9628_8799.n287 161.3
R323 a_n9628_8799.n300 a_n9628_8799.n299 161.3
R324 a_n9628_8799.n301 a_n9628_8799.n286 161.3
R325 a_n9628_8799.n303 a_n9628_8799.n302 161.3
R326 a_n9628_8799.n304 a_n9628_8799.n285 161.3
R327 a_n9628_8799.n305 a_n9628_8799.n284 161.3
R328 a_n9628_8799.n307 a_n9628_8799.n306 161.3
R329 a_n9628_8799.n308 a_n9628_8799.n283 161.3
R330 a_n9628_8799.n310 a_n9628_8799.n309 161.3
R331 a_n9628_8799.n311 a_n9628_8799.n282 161.3
R332 a_n9628_8799.n312 a_n9628_8799.n281 161.3
R333 a_n9628_8799.n314 a_n9628_8799.n313 161.3
R334 a_n9628_8799.n315 a_n9628_8799.n280 161.3
R335 a_n9628_8799.n317 a_n9628_8799.n316 161.3
R336 a_n9628_8799.n318 a_n9628_8799.n279 161.3
R337 a_n9628_8799.n319 a_n9628_8799.n278 161.3
R338 a_n9628_8799.n321 a_n9628_8799.n320 161.3
R339 a_n9628_8799.n322 a_n9628_8799.n277 161.3
R340 a_n9628_8799.n324 a_n9628_8799.n323 161.3
R341 a_n9628_8799.n325 a_n9628_8799.n276 161.3
R342 a_n9628_8799.n326 a_n9628_8799.n275 161.3
R343 a_n9628_8799.n328 a_n9628_8799.n327 161.3
R344 a_n9628_8799.n329 a_n9628_8799.n274 161.3
R345 a_n9628_8799.n331 a_n9628_8799.n330 161.3
R346 a_n9628_8799.n332 a_n9628_8799.n273 161.3
R347 a_n9628_8799.n334 a_n9628_8799.n333 161.3
R348 a_n9628_8799.n356 a_n9628_8799.n355 161.3
R349 a_n9628_8799.n357 a_n9628_8799.n352 161.3
R350 a_n9628_8799.n359 a_n9628_8799.n358 161.3
R351 a_n9628_8799.n360 a_n9628_8799.n351 161.3
R352 a_n9628_8799.n361 a_n9628_8799.n350 161.3
R353 a_n9628_8799.n363 a_n9628_8799.n362 161.3
R354 a_n9628_8799.n364 a_n9628_8799.n349 161.3
R355 a_n9628_8799.n366 a_n9628_8799.n365 161.3
R356 a_n9628_8799.n367 a_n9628_8799.n348 161.3
R357 a_n9628_8799.n368 a_n9628_8799.n347 161.3
R358 a_n9628_8799.n370 a_n9628_8799.n369 161.3
R359 a_n9628_8799.n371 a_n9628_8799.n346 161.3
R360 a_n9628_8799.n373 a_n9628_8799.n372 161.3
R361 a_n9628_8799.n374 a_n9628_8799.n345 161.3
R362 a_n9628_8799.n375 a_n9628_8799.n344 161.3
R363 a_n9628_8799.n377 a_n9628_8799.n376 161.3
R364 a_n9628_8799.n378 a_n9628_8799.n343 161.3
R365 a_n9628_8799.n380 a_n9628_8799.n379 161.3
R366 a_n9628_8799.n381 a_n9628_8799.n342 161.3
R367 a_n9628_8799.n382 a_n9628_8799.n341 161.3
R368 a_n9628_8799.n384 a_n9628_8799.n383 161.3
R369 a_n9628_8799.n385 a_n9628_8799.n340 161.3
R370 a_n9628_8799.n387 a_n9628_8799.n386 161.3
R371 a_n9628_8799.n388 a_n9628_8799.n339 161.3
R372 a_n9628_8799.n389 a_n9628_8799.n338 161.3
R373 a_n9628_8799.n391 a_n9628_8799.n390 161.3
R374 a_n9628_8799.n392 a_n9628_8799.n337 161.3
R375 a_n9628_8799.n394 a_n9628_8799.n393 161.3
R376 a_n9628_8799.n395 a_n9628_8799.n336 161.3
R377 a_n9628_8799.n397 a_n9628_8799.n396 161.3
R378 a_n9628_8799.n84 a_n9628_8799.n83 161.3
R379 a_n9628_8799.n82 a_n9628_8799.n23 161.3
R380 a_n9628_8799.n81 a_n9628_8799.n80 161.3
R381 a_n9628_8799.n79 a_n9628_8799.n24 161.3
R382 a_n9628_8799.n78 a_n9628_8799.n77 161.3
R383 a_n9628_8799.n76 a_n9628_8799.n25 161.3
R384 a_n9628_8799.n75 a_n9628_8799.n74 161.3
R385 a_n9628_8799.n73 a_n9628_8799.n26 161.3
R386 a_n9628_8799.n72 a_n9628_8799.n71 161.3
R387 a_n9628_8799.n70 a_n9628_8799.n27 161.3
R388 a_n9628_8799.n69 a_n9628_8799.n68 161.3
R389 a_n9628_8799.n67 a_n9628_8799.n28 161.3
R390 a_n9628_8799.n66 a_n9628_8799.n65 161.3
R391 a_n9628_8799.n64 a_n9628_8799.n29 161.3
R392 a_n9628_8799.n63 a_n9628_8799.n62 161.3
R393 a_n9628_8799.n61 a_n9628_8799.n30 161.3
R394 a_n9628_8799.n60 a_n9628_8799.n59 161.3
R395 a_n9628_8799.n58 a_n9628_8799.n31 161.3
R396 a_n9628_8799.n57 a_n9628_8799.n56 161.3
R397 a_n9628_8799.n55 a_n9628_8799.n32 161.3
R398 a_n9628_8799.n54 a_n9628_8799.n53 161.3
R399 a_n9628_8799.n52 a_n9628_8799.n33 161.3
R400 a_n9628_8799.n51 a_n9628_8799.n50 161.3
R401 a_n9628_8799.n49 a_n9628_8799.n34 161.3
R402 a_n9628_8799.n48 a_n9628_8799.n47 161.3
R403 a_n9628_8799.n46 a_n9628_8799.n35 161.3
R404 a_n9628_8799.n45 a_n9628_8799.n44 161.3
R405 a_n9628_8799.n43 a_n9628_8799.n36 161.3
R406 a_n9628_8799.n42 a_n9628_8799.n41 161.3
R407 a_n9628_8799.n40 a_n9628_8799.n37 161.3
R408 a_n9628_8799.n146 a_n9628_8799.n145 161.3
R409 a_n9628_8799.n144 a_n9628_8799.n85 161.3
R410 a_n9628_8799.n143 a_n9628_8799.n142 161.3
R411 a_n9628_8799.n141 a_n9628_8799.n86 161.3
R412 a_n9628_8799.n140 a_n9628_8799.n139 161.3
R413 a_n9628_8799.n138 a_n9628_8799.n87 161.3
R414 a_n9628_8799.n137 a_n9628_8799.n136 161.3
R415 a_n9628_8799.n135 a_n9628_8799.n88 161.3
R416 a_n9628_8799.n134 a_n9628_8799.n133 161.3
R417 a_n9628_8799.n132 a_n9628_8799.n89 161.3
R418 a_n9628_8799.n131 a_n9628_8799.n130 161.3
R419 a_n9628_8799.n129 a_n9628_8799.n90 161.3
R420 a_n9628_8799.n128 a_n9628_8799.n127 161.3
R421 a_n9628_8799.n126 a_n9628_8799.n91 161.3
R422 a_n9628_8799.n125 a_n9628_8799.n124 161.3
R423 a_n9628_8799.n123 a_n9628_8799.n92 161.3
R424 a_n9628_8799.n122 a_n9628_8799.n121 161.3
R425 a_n9628_8799.n120 a_n9628_8799.n93 161.3
R426 a_n9628_8799.n119 a_n9628_8799.n118 161.3
R427 a_n9628_8799.n117 a_n9628_8799.n94 161.3
R428 a_n9628_8799.n116 a_n9628_8799.n115 161.3
R429 a_n9628_8799.n114 a_n9628_8799.n95 161.3
R430 a_n9628_8799.n113 a_n9628_8799.n112 161.3
R431 a_n9628_8799.n111 a_n9628_8799.n96 161.3
R432 a_n9628_8799.n110 a_n9628_8799.n109 161.3
R433 a_n9628_8799.n108 a_n9628_8799.n97 161.3
R434 a_n9628_8799.n107 a_n9628_8799.n106 161.3
R435 a_n9628_8799.n105 a_n9628_8799.n98 161.3
R436 a_n9628_8799.n104 a_n9628_8799.n103 161.3
R437 a_n9628_8799.n102 a_n9628_8799.n99 161.3
R438 a_n9628_8799.n209 a_n9628_8799.n208 161.3
R439 a_n9628_8799.n207 a_n9628_8799.n148 161.3
R440 a_n9628_8799.n206 a_n9628_8799.n205 161.3
R441 a_n9628_8799.n204 a_n9628_8799.n149 161.3
R442 a_n9628_8799.n203 a_n9628_8799.n202 161.3
R443 a_n9628_8799.n201 a_n9628_8799.n150 161.3
R444 a_n9628_8799.n200 a_n9628_8799.n199 161.3
R445 a_n9628_8799.n198 a_n9628_8799.n151 161.3
R446 a_n9628_8799.n197 a_n9628_8799.n196 161.3
R447 a_n9628_8799.n195 a_n9628_8799.n152 161.3
R448 a_n9628_8799.n194 a_n9628_8799.n193 161.3
R449 a_n9628_8799.n192 a_n9628_8799.n153 161.3
R450 a_n9628_8799.n191 a_n9628_8799.n190 161.3
R451 a_n9628_8799.n189 a_n9628_8799.n154 161.3
R452 a_n9628_8799.n188 a_n9628_8799.n187 161.3
R453 a_n9628_8799.n186 a_n9628_8799.n155 161.3
R454 a_n9628_8799.n185 a_n9628_8799.n184 161.3
R455 a_n9628_8799.n183 a_n9628_8799.n156 161.3
R456 a_n9628_8799.n182 a_n9628_8799.n181 161.3
R457 a_n9628_8799.n180 a_n9628_8799.n157 161.3
R458 a_n9628_8799.n179 a_n9628_8799.n178 161.3
R459 a_n9628_8799.n177 a_n9628_8799.n158 161.3
R460 a_n9628_8799.n176 a_n9628_8799.n175 161.3
R461 a_n9628_8799.n174 a_n9628_8799.n159 161.3
R462 a_n9628_8799.n173 a_n9628_8799.n172 161.3
R463 a_n9628_8799.n171 a_n9628_8799.n160 161.3
R464 a_n9628_8799.n170 a_n9628_8799.n169 161.3
R465 a_n9628_8799.n168 a_n9628_8799.n161 161.3
R466 a_n9628_8799.n167 a_n9628_8799.n166 161.3
R467 a_n9628_8799.n165 a_n9628_8799.n162 161.3
R468 a_n9628_8799.n13 a_n9628_8799.n11 98.9633
R469 a_n9628_8799.n2 a_n9628_8799.n0 98.9631
R470 a_n9628_8799.n21 a_n9628_8799.n20 98.6055
R471 a_n9628_8799.n19 a_n9628_8799.n18 98.6055
R472 a_n9628_8799.n17 a_n9628_8799.n16 98.6055
R473 a_n9628_8799.n15 a_n9628_8799.n14 98.6055
R474 a_n9628_8799.n13 a_n9628_8799.n12 98.6055
R475 a_n9628_8799.n2 a_n9628_8799.n1 98.6055
R476 a_n9628_8799.n4 a_n9628_8799.n3 98.6055
R477 a_n9628_8799.n6 a_n9628_8799.n5 98.6055
R478 a_n9628_8799.n8 a_n9628_8799.n7 98.6055
R479 a_n9628_8799.n10 a_n9628_8799.n9 98.6055
R480 a_n9628_8799.n415 a_n9628_8799.n414 81.3766
R481 a_n9628_8799.n403 a_n9628_8799.n401 81.3764
R482 a_n9628_8799.n411 a_n9628_8799.n409 81.3764
R483 a_n9628_8799.n408 a_n9628_8799.n407 80.9324
R484 a_n9628_8799.n406 a_n9628_8799.n405 80.9324
R485 a_n9628_8799.n403 a_n9628_8799.n402 80.9324
R486 a_n9628_8799.n411 a_n9628_8799.n410 80.9324
R487 a_n9628_8799.n414 a_n9628_8799.n413 80.9324
R488 a_n9628_8799.n231 a_n9628_8799.n228 70.4033
R489 a_n9628_8799.n293 a_n9628_8799.n290 70.4033
R490 a_n9628_8799.n356 a_n9628_8799.n353 70.4033
R491 a_n9628_8799.n38 a_n9628_8799.n37 70.4033
R492 a_n9628_8799.n100 a_n9628_8799.n99 70.4033
R493 a_n9628_8799.n163 a_n9628_8799.n162 70.4033
R494 a_n9628_8799.n271 a_n9628_8799.n270 48.2005
R495 a_n9628_8799.n264 a_n9628_8799.n263 48.2005
R496 a_n9628_8799.n257 a_n9628_8799.n256 48.2005
R497 a_n9628_8799.n250 a_n9628_8799.n249 48.2005
R498 a_n9628_8799.n243 a_n9628_8799.n242 48.2005
R499 a_n9628_8799.n236 a_n9628_8799.n235 48.2005
R500 a_n9628_8799.n333 a_n9628_8799.n332 48.2005
R501 a_n9628_8799.n326 a_n9628_8799.n325 48.2005
R502 a_n9628_8799.n319 a_n9628_8799.n318 48.2005
R503 a_n9628_8799.n312 a_n9628_8799.n311 48.2005
R504 a_n9628_8799.n305 a_n9628_8799.n304 48.2005
R505 a_n9628_8799.n298 a_n9628_8799.n297 48.2005
R506 a_n9628_8799.n396 a_n9628_8799.n395 48.2005
R507 a_n9628_8799.n389 a_n9628_8799.n388 48.2005
R508 a_n9628_8799.n382 a_n9628_8799.n381 48.2005
R509 a_n9628_8799.n375 a_n9628_8799.n374 48.2005
R510 a_n9628_8799.n368 a_n9628_8799.n367 48.2005
R511 a_n9628_8799.n361 a_n9628_8799.n360 48.2005
R512 a_n9628_8799.n46 a_n9628_8799.n45 48.2005
R513 a_n9628_8799.n53 a_n9628_8799.n52 48.2005
R514 a_n9628_8799.n59 a_n9628_8799.n30 48.2005
R515 a_n9628_8799.n69 a_n9628_8799.n28 48.2005
R516 a_n9628_8799.n76 a_n9628_8799.n75 48.2005
R517 a_n9628_8799.n83 a_n9628_8799.n82 48.2005
R518 a_n9628_8799.n108 a_n9628_8799.n107 48.2005
R519 a_n9628_8799.n115 a_n9628_8799.n114 48.2005
R520 a_n9628_8799.n121 a_n9628_8799.n92 48.2005
R521 a_n9628_8799.n131 a_n9628_8799.n90 48.2005
R522 a_n9628_8799.n138 a_n9628_8799.n137 48.2005
R523 a_n9628_8799.n145 a_n9628_8799.n144 48.2005
R524 a_n9628_8799.n171 a_n9628_8799.n170 48.2005
R525 a_n9628_8799.n178 a_n9628_8799.n177 48.2005
R526 a_n9628_8799.n184 a_n9628_8799.n155 48.2005
R527 a_n9628_8799.n194 a_n9628_8799.n153 48.2005
R528 a_n9628_8799.n201 a_n9628_8799.n200 48.2005
R529 a_n9628_8799.n208 a_n9628_8799.n207 48.2005
R530 a_n9628_8799.n269 a_n9628_8799.n212 40.1672
R531 a_n9628_8799.n230 a_n9628_8799.n227 40.1672
R532 a_n9628_8799.n331 a_n9628_8799.n274 40.1672
R533 a_n9628_8799.n292 a_n9628_8799.n289 40.1672
R534 a_n9628_8799.n394 a_n9628_8799.n337 40.1672
R535 a_n9628_8799.n355 a_n9628_8799.n352 40.1672
R536 a_n9628_8799.n41 a_n9628_8799.n40 40.1672
R537 a_n9628_8799.n81 a_n9628_8799.n24 40.1672
R538 a_n9628_8799.n103 a_n9628_8799.n102 40.1672
R539 a_n9628_8799.n143 a_n9628_8799.n86 40.1672
R540 a_n9628_8799.n166 a_n9628_8799.n165 40.1672
R541 a_n9628_8799.n206 a_n9628_8799.n149 40.1672
R542 a_n9628_8799.n262 a_n9628_8799.n215 38.7066
R543 a_n9628_8799.n237 a_n9628_8799.n224 38.7066
R544 a_n9628_8799.n324 a_n9628_8799.n277 38.7066
R545 a_n9628_8799.n299 a_n9628_8799.n286 38.7066
R546 a_n9628_8799.n387 a_n9628_8799.n340 38.7066
R547 a_n9628_8799.n362 a_n9628_8799.n349 38.7066
R548 a_n9628_8799.n47 a_n9628_8799.n34 38.7066
R549 a_n9628_8799.n71 a_n9628_8799.n26 38.7066
R550 a_n9628_8799.n109 a_n9628_8799.n96 38.7066
R551 a_n9628_8799.n133 a_n9628_8799.n88 38.7066
R552 a_n9628_8799.n172 a_n9628_8799.n159 38.7066
R553 a_n9628_8799.n196 a_n9628_8799.n151 38.7066
R554 a_n9628_8799.n255 a_n9628_8799.n218 37.246
R555 a_n9628_8799.n244 a_n9628_8799.n221 37.246
R556 a_n9628_8799.n317 a_n9628_8799.n280 37.246
R557 a_n9628_8799.n306 a_n9628_8799.n283 37.246
R558 a_n9628_8799.n380 a_n9628_8799.n343 37.246
R559 a_n9628_8799.n369 a_n9628_8799.n346 37.246
R560 a_n9628_8799.n57 a_n9628_8799.n32 37.246
R561 a_n9628_8799.n65 a_n9628_8799.n64 37.246
R562 a_n9628_8799.n119 a_n9628_8799.n94 37.246
R563 a_n9628_8799.n127 a_n9628_8799.n126 37.246
R564 a_n9628_8799.n182 a_n9628_8799.n157 37.246
R565 a_n9628_8799.n190 a_n9628_8799.n189 37.246
R566 a_n9628_8799.n251 a_n9628_8799.n218 35.7853
R567 a_n9628_8799.n248 a_n9628_8799.n221 35.7853
R568 a_n9628_8799.n313 a_n9628_8799.n280 35.7853
R569 a_n9628_8799.n310 a_n9628_8799.n283 35.7853
R570 a_n9628_8799.n376 a_n9628_8799.n343 35.7853
R571 a_n9628_8799.n373 a_n9628_8799.n346 35.7853
R572 a_n9628_8799.n58 a_n9628_8799.n57 35.7853
R573 a_n9628_8799.n64 a_n9628_8799.n63 35.7853
R574 a_n9628_8799.n120 a_n9628_8799.n119 35.7853
R575 a_n9628_8799.n126 a_n9628_8799.n125 35.7853
R576 a_n9628_8799.n183 a_n9628_8799.n182 35.7853
R577 a_n9628_8799.n189 a_n9628_8799.n188 35.7853
R578 a_n9628_8799.n258 a_n9628_8799.n215 34.3247
R579 a_n9628_8799.n241 a_n9628_8799.n224 34.3247
R580 a_n9628_8799.n320 a_n9628_8799.n277 34.3247
R581 a_n9628_8799.n303 a_n9628_8799.n286 34.3247
R582 a_n9628_8799.n383 a_n9628_8799.n340 34.3247
R583 a_n9628_8799.n366 a_n9628_8799.n349 34.3247
R584 a_n9628_8799.n51 a_n9628_8799.n34 34.3247
R585 a_n9628_8799.n71 a_n9628_8799.n70 34.3247
R586 a_n9628_8799.n113 a_n9628_8799.n96 34.3247
R587 a_n9628_8799.n133 a_n9628_8799.n132 34.3247
R588 a_n9628_8799.n176 a_n9628_8799.n159 34.3247
R589 a_n9628_8799.n196 a_n9628_8799.n195 34.3247
R590 a_n9628_8799.n22 a_n9628_8799.n10 33.7114
R591 a_n9628_8799.n265 a_n9628_8799.n212 32.8641
R592 a_n9628_8799.n234 a_n9628_8799.n227 32.8641
R593 a_n9628_8799.n327 a_n9628_8799.n274 32.8641
R594 a_n9628_8799.n296 a_n9628_8799.n289 32.8641
R595 a_n9628_8799.n390 a_n9628_8799.n337 32.8641
R596 a_n9628_8799.n359 a_n9628_8799.n352 32.8641
R597 a_n9628_8799.n41 a_n9628_8799.n36 32.8641
R598 a_n9628_8799.n77 a_n9628_8799.n24 32.8641
R599 a_n9628_8799.n103 a_n9628_8799.n98 32.8641
R600 a_n9628_8799.n139 a_n9628_8799.n86 32.8641
R601 a_n9628_8799.n166 a_n9628_8799.n161 32.8641
R602 a_n9628_8799.n202 a_n9628_8799.n149 32.8641
R603 a_n9628_8799.n412 a_n9628_8799.n408 32.0866
R604 a_n9628_8799.n22 a_n9628_8799.n21 21.1779
R605 a_n9628_8799.n229 a_n9628_8799.n228 20.9576
R606 a_n9628_8799.n291 a_n9628_8799.n290 20.9576
R607 a_n9628_8799.n354 a_n9628_8799.n353 20.9576
R608 a_n9628_8799.n39 a_n9628_8799.n38 20.9576
R609 a_n9628_8799.n101 a_n9628_8799.n100 20.9576
R610 a_n9628_8799.n164 a_n9628_8799.n163 20.9576
R611 a_n9628_8799.n265 a_n9628_8799.n264 15.3369
R612 a_n9628_8799.n235 a_n9628_8799.n234 15.3369
R613 a_n9628_8799.n327 a_n9628_8799.n326 15.3369
R614 a_n9628_8799.n297 a_n9628_8799.n296 15.3369
R615 a_n9628_8799.n390 a_n9628_8799.n389 15.3369
R616 a_n9628_8799.n360 a_n9628_8799.n359 15.3369
R617 a_n9628_8799.n45 a_n9628_8799.n36 15.3369
R618 a_n9628_8799.n77 a_n9628_8799.n76 15.3369
R619 a_n9628_8799.n107 a_n9628_8799.n98 15.3369
R620 a_n9628_8799.n139 a_n9628_8799.n138 15.3369
R621 a_n9628_8799.n170 a_n9628_8799.n161 15.3369
R622 a_n9628_8799.n202 a_n9628_8799.n201 15.3369
R623 a_n9628_8799.n258 a_n9628_8799.n257 13.8763
R624 a_n9628_8799.n242 a_n9628_8799.n241 13.8763
R625 a_n9628_8799.n320 a_n9628_8799.n319 13.8763
R626 a_n9628_8799.n304 a_n9628_8799.n303 13.8763
R627 a_n9628_8799.n383 a_n9628_8799.n382 13.8763
R628 a_n9628_8799.n367 a_n9628_8799.n366 13.8763
R629 a_n9628_8799.n52 a_n9628_8799.n51 13.8763
R630 a_n9628_8799.n70 a_n9628_8799.n69 13.8763
R631 a_n9628_8799.n114 a_n9628_8799.n113 13.8763
R632 a_n9628_8799.n132 a_n9628_8799.n131 13.8763
R633 a_n9628_8799.n177 a_n9628_8799.n176 13.8763
R634 a_n9628_8799.n195 a_n9628_8799.n194 13.8763
R635 a_n9628_8799.n251 a_n9628_8799.n250 12.4157
R636 a_n9628_8799.n249 a_n9628_8799.n248 12.4157
R637 a_n9628_8799.n313 a_n9628_8799.n312 12.4157
R638 a_n9628_8799.n311 a_n9628_8799.n310 12.4157
R639 a_n9628_8799.n376 a_n9628_8799.n375 12.4157
R640 a_n9628_8799.n374 a_n9628_8799.n373 12.4157
R641 a_n9628_8799.n59 a_n9628_8799.n58 12.4157
R642 a_n9628_8799.n63 a_n9628_8799.n30 12.4157
R643 a_n9628_8799.n121 a_n9628_8799.n120 12.4157
R644 a_n9628_8799.n125 a_n9628_8799.n92 12.4157
R645 a_n9628_8799.n184 a_n9628_8799.n183 12.4157
R646 a_n9628_8799.n188 a_n9628_8799.n155 12.4157
R647 a_n9628_8799.n404 a_n9628_8799.n400 12.3339
R648 a_n9628_8799.n400 a_n9628_8799.n22 11.4887
R649 a_n9628_8799.n256 a_n9628_8799.n255 10.955
R650 a_n9628_8799.n244 a_n9628_8799.n243 10.955
R651 a_n9628_8799.n318 a_n9628_8799.n317 10.955
R652 a_n9628_8799.n306 a_n9628_8799.n305 10.955
R653 a_n9628_8799.n381 a_n9628_8799.n380 10.955
R654 a_n9628_8799.n369 a_n9628_8799.n368 10.955
R655 a_n9628_8799.n53 a_n9628_8799.n32 10.955
R656 a_n9628_8799.n65 a_n9628_8799.n28 10.955
R657 a_n9628_8799.n115 a_n9628_8799.n94 10.955
R658 a_n9628_8799.n127 a_n9628_8799.n90 10.955
R659 a_n9628_8799.n178 a_n9628_8799.n157 10.955
R660 a_n9628_8799.n190 a_n9628_8799.n153 10.955
R661 a_n9628_8799.n263 a_n9628_8799.n262 9.49444
R662 a_n9628_8799.n237 a_n9628_8799.n236 9.49444
R663 a_n9628_8799.n325 a_n9628_8799.n324 9.49444
R664 a_n9628_8799.n299 a_n9628_8799.n298 9.49444
R665 a_n9628_8799.n388 a_n9628_8799.n387 9.49444
R666 a_n9628_8799.n362 a_n9628_8799.n361 9.49444
R667 a_n9628_8799.n47 a_n9628_8799.n46 9.49444
R668 a_n9628_8799.n75 a_n9628_8799.n26 9.49444
R669 a_n9628_8799.n109 a_n9628_8799.n108 9.49444
R670 a_n9628_8799.n137 a_n9628_8799.n88 9.49444
R671 a_n9628_8799.n172 a_n9628_8799.n171 9.49444
R672 a_n9628_8799.n200 a_n9628_8799.n151 9.49444
R673 a_n9628_8799.n335 a_n9628_8799.n272 9.04406
R674 a_n9628_8799.n147 a_n9628_8799.n84 9.04406
R675 a_n9628_8799.n270 a_n9628_8799.n269 8.03383
R676 a_n9628_8799.n230 a_n9628_8799.n229 8.03383
R677 a_n9628_8799.n332 a_n9628_8799.n331 8.03383
R678 a_n9628_8799.n292 a_n9628_8799.n291 8.03383
R679 a_n9628_8799.n395 a_n9628_8799.n394 8.03383
R680 a_n9628_8799.n355 a_n9628_8799.n354 8.03383
R681 a_n9628_8799.n40 a_n9628_8799.n39 8.03383
R682 a_n9628_8799.n82 a_n9628_8799.n81 8.03383
R683 a_n9628_8799.n102 a_n9628_8799.n101 8.03383
R684 a_n9628_8799.n144 a_n9628_8799.n143 8.03383
R685 a_n9628_8799.n165 a_n9628_8799.n164 8.03383
R686 a_n9628_8799.n207 a_n9628_8799.n206 8.03383
R687 a_n9628_8799.n399 a_n9628_8799.n210 7.14965
R688 a_n9628_8799.n399 a_n9628_8799.n398 6.85731
R689 a_n9628_8799.n335 a_n9628_8799.n334 4.93611
R690 a_n9628_8799.n398 a_n9628_8799.n397 4.93611
R691 a_n9628_8799.n147 a_n9628_8799.n146 4.93611
R692 a_n9628_8799.n210 a_n9628_8799.n209 4.93611
R693 a_n9628_8799.n398 a_n9628_8799.n335 4.10845
R694 a_n9628_8799.n210 a_n9628_8799.n147 4.10845
R695 a_n9628_8799.n20 a_n9628_8799.t7 3.61217
R696 a_n9628_8799.n20 a_n9628_8799.t1 3.61217
R697 a_n9628_8799.n18 a_n9628_8799.t6 3.61217
R698 a_n9628_8799.n18 a_n9628_8799.t37 3.61217
R699 a_n9628_8799.n16 a_n9628_8799.t35 3.61217
R700 a_n9628_8799.n16 a_n9628_8799.t10 3.61217
R701 a_n9628_8799.n14 a_n9628_8799.t2 3.61217
R702 a_n9628_8799.n14 a_n9628_8799.t16 3.61217
R703 a_n9628_8799.n12 a_n9628_8799.t5 3.61217
R704 a_n9628_8799.n12 a_n9628_8799.t4 3.61217
R705 a_n9628_8799.n11 a_n9628_8799.t17 3.61217
R706 a_n9628_8799.n11 a_n9628_8799.t39 3.61217
R707 a_n9628_8799.n0 a_n9628_8799.t13 3.61217
R708 a_n9628_8799.n0 a_n9628_8799.t12 3.61217
R709 a_n9628_8799.n1 a_n9628_8799.t38 3.61217
R710 a_n9628_8799.n1 a_n9628_8799.t18 3.61217
R711 a_n9628_8799.n3 a_n9628_8799.t0 3.61217
R712 a_n9628_8799.n3 a_n9628_8799.t15 3.61217
R713 a_n9628_8799.n5 a_n9628_8799.t11 3.61217
R714 a_n9628_8799.n5 a_n9628_8799.t14 3.61217
R715 a_n9628_8799.n7 a_n9628_8799.t8 3.61217
R716 a_n9628_8799.n7 a_n9628_8799.t36 3.61217
R717 a_n9628_8799.n9 a_n9628_8799.t3 3.61217
R718 a_n9628_8799.n9 a_n9628_8799.t9 3.61217
R719 a_n9628_8799.n400 a_n9628_8799.n399 3.4105
R720 a_n9628_8799.n409 a_n9628_8799.t29 2.82907
R721 a_n9628_8799.n409 a_n9628_8799.t27 2.82907
R722 a_n9628_8799.n410 a_n9628_8799.t22 2.82907
R723 a_n9628_8799.n410 a_n9628_8799.t26 2.82907
R724 a_n9628_8799.n413 a_n9628_8799.t33 2.82907
R725 a_n9628_8799.n413 a_n9628_8799.t23 2.82907
R726 a_n9628_8799.n407 a_n9628_8799.t32 2.82907
R727 a_n9628_8799.n407 a_n9628_8799.t28 2.82907
R728 a_n9628_8799.n405 a_n9628_8799.t19 2.82907
R729 a_n9628_8799.n405 a_n9628_8799.t31 2.82907
R730 a_n9628_8799.n402 a_n9628_8799.t20 2.82907
R731 a_n9628_8799.n402 a_n9628_8799.t21 2.82907
R732 a_n9628_8799.n401 a_n9628_8799.t24 2.82907
R733 a_n9628_8799.n401 a_n9628_8799.t25 2.82907
R734 a_n9628_8799.n415 a_n9628_8799.t30 2.82907
R735 a_n9628_8799.t34 a_n9628_8799.n415 2.82907
R736 a_n9628_8799.n408 a_n9628_8799.n406 0.444466
R737 a_n9628_8799.n15 a_n9628_8799.n13 0.358259
R738 a_n9628_8799.n17 a_n9628_8799.n15 0.358259
R739 a_n9628_8799.n19 a_n9628_8799.n17 0.358259
R740 a_n9628_8799.n21 a_n9628_8799.n19 0.358259
R741 a_n9628_8799.n10 a_n9628_8799.n8 0.358259
R742 a_n9628_8799.n8 a_n9628_8799.n6 0.358259
R743 a_n9628_8799.n6 a_n9628_8799.n4 0.358259
R744 a_n9628_8799.n4 a_n9628_8799.n2 0.358259
R745 a_n9628_8799.n404 a_n9628_8799.n403 0.222483
R746 a_n9628_8799.n406 a_n9628_8799.n404 0.222483
R747 a_n9628_8799.n414 a_n9628_8799.n412 0.222483
R748 a_n9628_8799.n412 a_n9628_8799.n411 0.222483
R749 a_n9628_8799.n272 a_n9628_8799.n211 0.189894
R750 a_n9628_8799.n268 a_n9628_8799.n211 0.189894
R751 a_n9628_8799.n268 a_n9628_8799.n267 0.189894
R752 a_n9628_8799.n267 a_n9628_8799.n266 0.189894
R753 a_n9628_8799.n266 a_n9628_8799.n213 0.189894
R754 a_n9628_8799.n214 a_n9628_8799.n213 0.189894
R755 a_n9628_8799.n261 a_n9628_8799.n214 0.189894
R756 a_n9628_8799.n261 a_n9628_8799.n260 0.189894
R757 a_n9628_8799.n260 a_n9628_8799.n259 0.189894
R758 a_n9628_8799.n259 a_n9628_8799.n216 0.189894
R759 a_n9628_8799.n217 a_n9628_8799.n216 0.189894
R760 a_n9628_8799.n254 a_n9628_8799.n217 0.189894
R761 a_n9628_8799.n254 a_n9628_8799.n253 0.189894
R762 a_n9628_8799.n253 a_n9628_8799.n252 0.189894
R763 a_n9628_8799.n252 a_n9628_8799.n219 0.189894
R764 a_n9628_8799.n220 a_n9628_8799.n219 0.189894
R765 a_n9628_8799.n247 a_n9628_8799.n220 0.189894
R766 a_n9628_8799.n247 a_n9628_8799.n246 0.189894
R767 a_n9628_8799.n246 a_n9628_8799.n245 0.189894
R768 a_n9628_8799.n245 a_n9628_8799.n222 0.189894
R769 a_n9628_8799.n223 a_n9628_8799.n222 0.189894
R770 a_n9628_8799.n240 a_n9628_8799.n223 0.189894
R771 a_n9628_8799.n240 a_n9628_8799.n239 0.189894
R772 a_n9628_8799.n239 a_n9628_8799.n238 0.189894
R773 a_n9628_8799.n238 a_n9628_8799.n225 0.189894
R774 a_n9628_8799.n226 a_n9628_8799.n225 0.189894
R775 a_n9628_8799.n233 a_n9628_8799.n226 0.189894
R776 a_n9628_8799.n233 a_n9628_8799.n232 0.189894
R777 a_n9628_8799.n232 a_n9628_8799.n231 0.189894
R778 a_n9628_8799.n334 a_n9628_8799.n273 0.189894
R779 a_n9628_8799.n330 a_n9628_8799.n273 0.189894
R780 a_n9628_8799.n330 a_n9628_8799.n329 0.189894
R781 a_n9628_8799.n329 a_n9628_8799.n328 0.189894
R782 a_n9628_8799.n328 a_n9628_8799.n275 0.189894
R783 a_n9628_8799.n276 a_n9628_8799.n275 0.189894
R784 a_n9628_8799.n323 a_n9628_8799.n276 0.189894
R785 a_n9628_8799.n323 a_n9628_8799.n322 0.189894
R786 a_n9628_8799.n322 a_n9628_8799.n321 0.189894
R787 a_n9628_8799.n321 a_n9628_8799.n278 0.189894
R788 a_n9628_8799.n279 a_n9628_8799.n278 0.189894
R789 a_n9628_8799.n316 a_n9628_8799.n279 0.189894
R790 a_n9628_8799.n316 a_n9628_8799.n315 0.189894
R791 a_n9628_8799.n315 a_n9628_8799.n314 0.189894
R792 a_n9628_8799.n314 a_n9628_8799.n281 0.189894
R793 a_n9628_8799.n282 a_n9628_8799.n281 0.189894
R794 a_n9628_8799.n309 a_n9628_8799.n282 0.189894
R795 a_n9628_8799.n309 a_n9628_8799.n308 0.189894
R796 a_n9628_8799.n308 a_n9628_8799.n307 0.189894
R797 a_n9628_8799.n307 a_n9628_8799.n284 0.189894
R798 a_n9628_8799.n285 a_n9628_8799.n284 0.189894
R799 a_n9628_8799.n302 a_n9628_8799.n285 0.189894
R800 a_n9628_8799.n302 a_n9628_8799.n301 0.189894
R801 a_n9628_8799.n301 a_n9628_8799.n300 0.189894
R802 a_n9628_8799.n300 a_n9628_8799.n287 0.189894
R803 a_n9628_8799.n288 a_n9628_8799.n287 0.189894
R804 a_n9628_8799.n295 a_n9628_8799.n288 0.189894
R805 a_n9628_8799.n295 a_n9628_8799.n294 0.189894
R806 a_n9628_8799.n294 a_n9628_8799.n293 0.189894
R807 a_n9628_8799.n397 a_n9628_8799.n336 0.189894
R808 a_n9628_8799.n393 a_n9628_8799.n336 0.189894
R809 a_n9628_8799.n393 a_n9628_8799.n392 0.189894
R810 a_n9628_8799.n392 a_n9628_8799.n391 0.189894
R811 a_n9628_8799.n391 a_n9628_8799.n338 0.189894
R812 a_n9628_8799.n339 a_n9628_8799.n338 0.189894
R813 a_n9628_8799.n386 a_n9628_8799.n339 0.189894
R814 a_n9628_8799.n386 a_n9628_8799.n385 0.189894
R815 a_n9628_8799.n385 a_n9628_8799.n384 0.189894
R816 a_n9628_8799.n384 a_n9628_8799.n341 0.189894
R817 a_n9628_8799.n342 a_n9628_8799.n341 0.189894
R818 a_n9628_8799.n379 a_n9628_8799.n342 0.189894
R819 a_n9628_8799.n379 a_n9628_8799.n378 0.189894
R820 a_n9628_8799.n378 a_n9628_8799.n377 0.189894
R821 a_n9628_8799.n377 a_n9628_8799.n344 0.189894
R822 a_n9628_8799.n345 a_n9628_8799.n344 0.189894
R823 a_n9628_8799.n372 a_n9628_8799.n345 0.189894
R824 a_n9628_8799.n372 a_n9628_8799.n371 0.189894
R825 a_n9628_8799.n371 a_n9628_8799.n370 0.189894
R826 a_n9628_8799.n370 a_n9628_8799.n347 0.189894
R827 a_n9628_8799.n348 a_n9628_8799.n347 0.189894
R828 a_n9628_8799.n365 a_n9628_8799.n348 0.189894
R829 a_n9628_8799.n365 a_n9628_8799.n364 0.189894
R830 a_n9628_8799.n364 a_n9628_8799.n363 0.189894
R831 a_n9628_8799.n363 a_n9628_8799.n350 0.189894
R832 a_n9628_8799.n351 a_n9628_8799.n350 0.189894
R833 a_n9628_8799.n358 a_n9628_8799.n351 0.189894
R834 a_n9628_8799.n358 a_n9628_8799.n357 0.189894
R835 a_n9628_8799.n357 a_n9628_8799.n356 0.189894
R836 a_n9628_8799.n42 a_n9628_8799.n37 0.189894
R837 a_n9628_8799.n43 a_n9628_8799.n42 0.189894
R838 a_n9628_8799.n44 a_n9628_8799.n43 0.189894
R839 a_n9628_8799.n44 a_n9628_8799.n35 0.189894
R840 a_n9628_8799.n48 a_n9628_8799.n35 0.189894
R841 a_n9628_8799.n49 a_n9628_8799.n48 0.189894
R842 a_n9628_8799.n50 a_n9628_8799.n49 0.189894
R843 a_n9628_8799.n50 a_n9628_8799.n33 0.189894
R844 a_n9628_8799.n54 a_n9628_8799.n33 0.189894
R845 a_n9628_8799.n55 a_n9628_8799.n54 0.189894
R846 a_n9628_8799.n56 a_n9628_8799.n55 0.189894
R847 a_n9628_8799.n56 a_n9628_8799.n31 0.189894
R848 a_n9628_8799.n60 a_n9628_8799.n31 0.189894
R849 a_n9628_8799.n61 a_n9628_8799.n60 0.189894
R850 a_n9628_8799.n62 a_n9628_8799.n61 0.189894
R851 a_n9628_8799.n62 a_n9628_8799.n29 0.189894
R852 a_n9628_8799.n66 a_n9628_8799.n29 0.189894
R853 a_n9628_8799.n67 a_n9628_8799.n66 0.189894
R854 a_n9628_8799.n68 a_n9628_8799.n67 0.189894
R855 a_n9628_8799.n68 a_n9628_8799.n27 0.189894
R856 a_n9628_8799.n72 a_n9628_8799.n27 0.189894
R857 a_n9628_8799.n73 a_n9628_8799.n72 0.189894
R858 a_n9628_8799.n74 a_n9628_8799.n73 0.189894
R859 a_n9628_8799.n74 a_n9628_8799.n25 0.189894
R860 a_n9628_8799.n78 a_n9628_8799.n25 0.189894
R861 a_n9628_8799.n79 a_n9628_8799.n78 0.189894
R862 a_n9628_8799.n80 a_n9628_8799.n79 0.189894
R863 a_n9628_8799.n80 a_n9628_8799.n23 0.189894
R864 a_n9628_8799.n84 a_n9628_8799.n23 0.189894
R865 a_n9628_8799.n104 a_n9628_8799.n99 0.189894
R866 a_n9628_8799.n105 a_n9628_8799.n104 0.189894
R867 a_n9628_8799.n106 a_n9628_8799.n105 0.189894
R868 a_n9628_8799.n106 a_n9628_8799.n97 0.189894
R869 a_n9628_8799.n110 a_n9628_8799.n97 0.189894
R870 a_n9628_8799.n111 a_n9628_8799.n110 0.189894
R871 a_n9628_8799.n112 a_n9628_8799.n111 0.189894
R872 a_n9628_8799.n112 a_n9628_8799.n95 0.189894
R873 a_n9628_8799.n116 a_n9628_8799.n95 0.189894
R874 a_n9628_8799.n117 a_n9628_8799.n116 0.189894
R875 a_n9628_8799.n118 a_n9628_8799.n117 0.189894
R876 a_n9628_8799.n118 a_n9628_8799.n93 0.189894
R877 a_n9628_8799.n122 a_n9628_8799.n93 0.189894
R878 a_n9628_8799.n123 a_n9628_8799.n122 0.189894
R879 a_n9628_8799.n124 a_n9628_8799.n123 0.189894
R880 a_n9628_8799.n124 a_n9628_8799.n91 0.189894
R881 a_n9628_8799.n128 a_n9628_8799.n91 0.189894
R882 a_n9628_8799.n129 a_n9628_8799.n128 0.189894
R883 a_n9628_8799.n130 a_n9628_8799.n129 0.189894
R884 a_n9628_8799.n130 a_n9628_8799.n89 0.189894
R885 a_n9628_8799.n134 a_n9628_8799.n89 0.189894
R886 a_n9628_8799.n135 a_n9628_8799.n134 0.189894
R887 a_n9628_8799.n136 a_n9628_8799.n135 0.189894
R888 a_n9628_8799.n136 a_n9628_8799.n87 0.189894
R889 a_n9628_8799.n140 a_n9628_8799.n87 0.189894
R890 a_n9628_8799.n141 a_n9628_8799.n140 0.189894
R891 a_n9628_8799.n142 a_n9628_8799.n141 0.189894
R892 a_n9628_8799.n142 a_n9628_8799.n85 0.189894
R893 a_n9628_8799.n146 a_n9628_8799.n85 0.189894
R894 a_n9628_8799.n167 a_n9628_8799.n162 0.189894
R895 a_n9628_8799.n168 a_n9628_8799.n167 0.189894
R896 a_n9628_8799.n169 a_n9628_8799.n168 0.189894
R897 a_n9628_8799.n169 a_n9628_8799.n160 0.189894
R898 a_n9628_8799.n173 a_n9628_8799.n160 0.189894
R899 a_n9628_8799.n174 a_n9628_8799.n173 0.189894
R900 a_n9628_8799.n175 a_n9628_8799.n174 0.189894
R901 a_n9628_8799.n175 a_n9628_8799.n158 0.189894
R902 a_n9628_8799.n179 a_n9628_8799.n158 0.189894
R903 a_n9628_8799.n180 a_n9628_8799.n179 0.189894
R904 a_n9628_8799.n181 a_n9628_8799.n180 0.189894
R905 a_n9628_8799.n181 a_n9628_8799.n156 0.189894
R906 a_n9628_8799.n185 a_n9628_8799.n156 0.189894
R907 a_n9628_8799.n186 a_n9628_8799.n185 0.189894
R908 a_n9628_8799.n187 a_n9628_8799.n186 0.189894
R909 a_n9628_8799.n187 a_n9628_8799.n154 0.189894
R910 a_n9628_8799.n191 a_n9628_8799.n154 0.189894
R911 a_n9628_8799.n192 a_n9628_8799.n191 0.189894
R912 a_n9628_8799.n193 a_n9628_8799.n192 0.189894
R913 a_n9628_8799.n193 a_n9628_8799.n152 0.189894
R914 a_n9628_8799.n197 a_n9628_8799.n152 0.189894
R915 a_n9628_8799.n198 a_n9628_8799.n197 0.189894
R916 a_n9628_8799.n199 a_n9628_8799.n198 0.189894
R917 a_n9628_8799.n199 a_n9628_8799.n150 0.189894
R918 a_n9628_8799.n203 a_n9628_8799.n150 0.189894
R919 a_n9628_8799.n204 a_n9628_8799.n203 0.189894
R920 a_n9628_8799.n205 a_n9628_8799.n204 0.189894
R921 a_n9628_8799.n205 a_n9628_8799.n148 0.189894
R922 a_n9628_8799.n209 a_n9628_8799.n148 0.189894
R923 gnd.n7021 gnd.n394 1810.87
R924 gnd.n2339 gnd.n2338 927.927
R925 gnd.n7484 gnd.n172 838.452
R926 gnd.n7471 gnd.n170 838.452
R927 gnd.n5010 gnd.n3022 838.452
R928 gnd.n5079 gnd.n3024 838.452
R929 gnd.n6166 gnd.n2575 838.452
R930 gnd.n6086 gnd.n2573 838.452
R931 gnd.n3865 gnd.n2365 838.452
R932 gnd.n3907 gnd.n2367 838.452
R933 gnd.n7486 gnd.n167 783.196
R934 gnd.n7346 gnd.n169 783.196
R935 gnd.n5561 gnd.n3021 783.196
R936 gnd.n5842 gnd.n3025 783.196
R937 gnd.n6168 gnd.n2570 783.196
R938 gnd.n2780 gnd.n2572 783.196
R939 gnd.n4119 gnd.n2364 783.196
R940 gnd.n6295 gnd.n2368 783.196
R941 gnd.n6147 gnd.n2604 771.183
R942 gnd.n5860 gnd.n2999 771.183
R943 gnd.n6151 gnd.n2586 771.183
R944 gnd.n5167 gnd.n3001 771.183
R945 gnd.n2246 gnd.n878 766.379
R946 gnd.n2249 gnd.n2248 766.379
R947 gnd.n1486 gnd.n1389 766.379
R948 gnd.n1482 gnd.n1387 766.379
R949 gnd.n2337 gnd.n900 756.769
R950 gnd.n2240 gnd.n2239 756.769
R951 gnd.n1579 gnd.n1296 756.769
R952 gnd.n1577 gnd.n1299 756.769
R953 gnd.n6499 gnd.n706 737.549
R954 gnd.n7020 gnd.n395 737.549
R955 gnd.n7231 gnd.n267 737.549
R956 gnd.n6323 gnd.n871 737.549
R957 gnd.n6495 gnd.n706 585
R958 gnd.n706 gnd.n705 585
R959 gnd.n6494 gnd.n6493 585
R960 gnd.n6493 gnd.n6492 585
R961 gnd.n709 gnd.n708 585
R962 gnd.n6491 gnd.n709 585
R963 gnd.n6489 gnd.n6488 585
R964 gnd.n6490 gnd.n6489 585
R965 gnd.n6487 gnd.n711 585
R966 gnd.n711 gnd.n710 585
R967 gnd.n6486 gnd.n6485 585
R968 gnd.n6485 gnd.n6484 585
R969 gnd.n717 gnd.n716 585
R970 gnd.n6483 gnd.n717 585
R971 gnd.n6481 gnd.n6480 585
R972 gnd.n6482 gnd.n6481 585
R973 gnd.n6479 gnd.n719 585
R974 gnd.n719 gnd.n718 585
R975 gnd.n6478 gnd.n6477 585
R976 gnd.n6477 gnd.n6476 585
R977 gnd.n725 gnd.n724 585
R978 gnd.n6475 gnd.n725 585
R979 gnd.n6473 gnd.n6472 585
R980 gnd.n6474 gnd.n6473 585
R981 gnd.n6471 gnd.n727 585
R982 gnd.n727 gnd.n726 585
R983 gnd.n6470 gnd.n6469 585
R984 gnd.n6469 gnd.n6468 585
R985 gnd.n733 gnd.n732 585
R986 gnd.n6467 gnd.n733 585
R987 gnd.n6465 gnd.n6464 585
R988 gnd.n6466 gnd.n6465 585
R989 gnd.n6463 gnd.n735 585
R990 gnd.n735 gnd.n734 585
R991 gnd.n6462 gnd.n6461 585
R992 gnd.n6461 gnd.n6460 585
R993 gnd.n741 gnd.n740 585
R994 gnd.n6459 gnd.n741 585
R995 gnd.n6457 gnd.n6456 585
R996 gnd.n6458 gnd.n6457 585
R997 gnd.n6455 gnd.n743 585
R998 gnd.n743 gnd.n742 585
R999 gnd.n6454 gnd.n6453 585
R1000 gnd.n6453 gnd.n6452 585
R1001 gnd.n749 gnd.n748 585
R1002 gnd.n6451 gnd.n749 585
R1003 gnd.n6449 gnd.n6448 585
R1004 gnd.n6450 gnd.n6449 585
R1005 gnd.n6447 gnd.n751 585
R1006 gnd.n751 gnd.n750 585
R1007 gnd.n6446 gnd.n6445 585
R1008 gnd.n6445 gnd.n6444 585
R1009 gnd.n757 gnd.n756 585
R1010 gnd.n6443 gnd.n757 585
R1011 gnd.n6441 gnd.n6440 585
R1012 gnd.n6442 gnd.n6441 585
R1013 gnd.n6439 gnd.n759 585
R1014 gnd.n759 gnd.n758 585
R1015 gnd.n6438 gnd.n6437 585
R1016 gnd.n6437 gnd.n6436 585
R1017 gnd.n765 gnd.n764 585
R1018 gnd.n6435 gnd.n765 585
R1019 gnd.n6433 gnd.n6432 585
R1020 gnd.n6434 gnd.n6433 585
R1021 gnd.n6431 gnd.n767 585
R1022 gnd.n767 gnd.n766 585
R1023 gnd.n6430 gnd.n6429 585
R1024 gnd.n6429 gnd.n6428 585
R1025 gnd.n773 gnd.n772 585
R1026 gnd.n6427 gnd.n773 585
R1027 gnd.n6425 gnd.n6424 585
R1028 gnd.n6426 gnd.n6425 585
R1029 gnd.n6423 gnd.n775 585
R1030 gnd.n775 gnd.n774 585
R1031 gnd.n6422 gnd.n6421 585
R1032 gnd.n6421 gnd.n6420 585
R1033 gnd.n781 gnd.n780 585
R1034 gnd.n6419 gnd.n781 585
R1035 gnd.n6417 gnd.n6416 585
R1036 gnd.n6418 gnd.n6417 585
R1037 gnd.n6415 gnd.n783 585
R1038 gnd.n783 gnd.n782 585
R1039 gnd.n6414 gnd.n6413 585
R1040 gnd.n6413 gnd.n6412 585
R1041 gnd.n789 gnd.n788 585
R1042 gnd.n6411 gnd.n789 585
R1043 gnd.n6409 gnd.n6408 585
R1044 gnd.n6410 gnd.n6409 585
R1045 gnd.n6407 gnd.n791 585
R1046 gnd.n791 gnd.n790 585
R1047 gnd.n6406 gnd.n6405 585
R1048 gnd.n6405 gnd.n6404 585
R1049 gnd.n797 gnd.n796 585
R1050 gnd.n6403 gnd.n797 585
R1051 gnd.n6401 gnd.n6400 585
R1052 gnd.n6402 gnd.n6401 585
R1053 gnd.n6399 gnd.n799 585
R1054 gnd.n799 gnd.n798 585
R1055 gnd.n6398 gnd.n6397 585
R1056 gnd.n6397 gnd.n6396 585
R1057 gnd.n805 gnd.n804 585
R1058 gnd.n6395 gnd.n805 585
R1059 gnd.n6393 gnd.n6392 585
R1060 gnd.n6394 gnd.n6393 585
R1061 gnd.n6391 gnd.n807 585
R1062 gnd.n807 gnd.n806 585
R1063 gnd.n6390 gnd.n6389 585
R1064 gnd.n6389 gnd.n6388 585
R1065 gnd.n813 gnd.n812 585
R1066 gnd.n6387 gnd.n813 585
R1067 gnd.n6385 gnd.n6384 585
R1068 gnd.n6386 gnd.n6385 585
R1069 gnd.n6383 gnd.n815 585
R1070 gnd.n815 gnd.n814 585
R1071 gnd.n6382 gnd.n6381 585
R1072 gnd.n6381 gnd.n6380 585
R1073 gnd.n821 gnd.n820 585
R1074 gnd.n6379 gnd.n821 585
R1075 gnd.n6377 gnd.n6376 585
R1076 gnd.n6378 gnd.n6377 585
R1077 gnd.n6375 gnd.n823 585
R1078 gnd.n823 gnd.n822 585
R1079 gnd.n6374 gnd.n6373 585
R1080 gnd.n6373 gnd.n6372 585
R1081 gnd.n829 gnd.n828 585
R1082 gnd.n6371 gnd.n829 585
R1083 gnd.n6369 gnd.n6368 585
R1084 gnd.n6370 gnd.n6369 585
R1085 gnd.n6367 gnd.n831 585
R1086 gnd.n831 gnd.n830 585
R1087 gnd.n6366 gnd.n6365 585
R1088 gnd.n6365 gnd.n6364 585
R1089 gnd.n837 gnd.n836 585
R1090 gnd.n6363 gnd.n837 585
R1091 gnd.n6361 gnd.n6360 585
R1092 gnd.n6362 gnd.n6361 585
R1093 gnd.n6359 gnd.n839 585
R1094 gnd.n839 gnd.n838 585
R1095 gnd.n6358 gnd.n6357 585
R1096 gnd.n6357 gnd.n6356 585
R1097 gnd.n845 gnd.n844 585
R1098 gnd.n6355 gnd.n845 585
R1099 gnd.n6353 gnd.n6352 585
R1100 gnd.n6354 gnd.n6353 585
R1101 gnd.n6351 gnd.n847 585
R1102 gnd.n847 gnd.n846 585
R1103 gnd.n6350 gnd.n6349 585
R1104 gnd.n6349 gnd.n6348 585
R1105 gnd.n853 gnd.n852 585
R1106 gnd.n6347 gnd.n853 585
R1107 gnd.n6345 gnd.n6344 585
R1108 gnd.n6346 gnd.n6345 585
R1109 gnd.n6343 gnd.n855 585
R1110 gnd.n855 gnd.n854 585
R1111 gnd.n6342 gnd.n6341 585
R1112 gnd.n6341 gnd.n6340 585
R1113 gnd.n861 gnd.n860 585
R1114 gnd.n6339 gnd.n861 585
R1115 gnd.n6337 gnd.n6336 585
R1116 gnd.n6338 gnd.n6337 585
R1117 gnd.n6335 gnd.n863 585
R1118 gnd.n863 gnd.n862 585
R1119 gnd.n6334 gnd.n6333 585
R1120 gnd.n6333 gnd.n6332 585
R1121 gnd.n869 gnd.n868 585
R1122 gnd.n6331 gnd.n869 585
R1123 gnd.n6329 gnd.n6328 585
R1124 gnd.n6330 gnd.n6329 585
R1125 gnd.n6499 gnd.n6498 585
R1126 gnd.n6500 gnd.n6499 585
R1127 gnd.n704 gnd.n703 585
R1128 gnd.n6501 gnd.n704 585
R1129 gnd.n6504 gnd.n6503 585
R1130 gnd.n6503 gnd.n6502 585
R1131 gnd.n701 gnd.n700 585
R1132 gnd.n700 gnd.n699 585
R1133 gnd.n6509 gnd.n6508 585
R1134 gnd.n6510 gnd.n6509 585
R1135 gnd.n698 gnd.n697 585
R1136 gnd.n6511 gnd.n698 585
R1137 gnd.n6514 gnd.n6513 585
R1138 gnd.n6513 gnd.n6512 585
R1139 gnd.n695 gnd.n694 585
R1140 gnd.n694 gnd.n693 585
R1141 gnd.n6519 gnd.n6518 585
R1142 gnd.n6520 gnd.n6519 585
R1143 gnd.n692 gnd.n691 585
R1144 gnd.n6521 gnd.n692 585
R1145 gnd.n6524 gnd.n6523 585
R1146 gnd.n6523 gnd.n6522 585
R1147 gnd.n689 gnd.n688 585
R1148 gnd.n688 gnd.n687 585
R1149 gnd.n6529 gnd.n6528 585
R1150 gnd.n6530 gnd.n6529 585
R1151 gnd.n686 gnd.n685 585
R1152 gnd.n6531 gnd.n686 585
R1153 gnd.n6534 gnd.n6533 585
R1154 gnd.n6533 gnd.n6532 585
R1155 gnd.n683 gnd.n682 585
R1156 gnd.n682 gnd.n681 585
R1157 gnd.n6539 gnd.n6538 585
R1158 gnd.n6540 gnd.n6539 585
R1159 gnd.n680 gnd.n679 585
R1160 gnd.n6541 gnd.n680 585
R1161 gnd.n6544 gnd.n6543 585
R1162 gnd.n6543 gnd.n6542 585
R1163 gnd.n677 gnd.n676 585
R1164 gnd.n676 gnd.n675 585
R1165 gnd.n6549 gnd.n6548 585
R1166 gnd.n6550 gnd.n6549 585
R1167 gnd.n674 gnd.n673 585
R1168 gnd.n6551 gnd.n674 585
R1169 gnd.n6554 gnd.n6553 585
R1170 gnd.n6553 gnd.n6552 585
R1171 gnd.n671 gnd.n670 585
R1172 gnd.n670 gnd.n669 585
R1173 gnd.n6559 gnd.n6558 585
R1174 gnd.n6560 gnd.n6559 585
R1175 gnd.n668 gnd.n667 585
R1176 gnd.n6561 gnd.n668 585
R1177 gnd.n6564 gnd.n6563 585
R1178 gnd.n6563 gnd.n6562 585
R1179 gnd.n665 gnd.n664 585
R1180 gnd.n664 gnd.n663 585
R1181 gnd.n6569 gnd.n6568 585
R1182 gnd.n6570 gnd.n6569 585
R1183 gnd.n662 gnd.n661 585
R1184 gnd.n6571 gnd.n662 585
R1185 gnd.n6574 gnd.n6573 585
R1186 gnd.n6573 gnd.n6572 585
R1187 gnd.n659 gnd.n658 585
R1188 gnd.n658 gnd.n657 585
R1189 gnd.n6579 gnd.n6578 585
R1190 gnd.n6580 gnd.n6579 585
R1191 gnd.n656 gnd.n655 585
R1192 gnd.n6581 gnd.n656 585
R1193 gnd.n6584 gnd.n6583 585
R1194 gnd.n6583 gnd.n6582 585
R1195 gnd.n653 gnd.n652 585
R1196 gnd.n652 gnd.n651 585
R1197 gnd.n6589 gnd.n6588 585
R1198 gnd.n6590 gnd.n6589 585
R1199 gnd.n650 gnd.n649 585
R1200 gnd.n6591 gnd.n650 585
R1201 gnd.n6594 gnd.n6593 585
R1202 gnd.n6593 gnd.n6592 585
R1203 gnd.n647 gnd.n646 585
R1204 gnd.n646 gnd.n645 585
R1205 gnd.n6599 gnd.n6598 585
R1206 gnd.n6600 gnd.n6599 585
R1207 gnd.n644 gnd.n643 585
R1208 gnd.n6601 gnd.n644 585
R1209 gnd.n6604 gnd.n6603 585
R1210 gnd.n6603 gnd.n6602 585
R1211 gnd.n641 gnd.n640 585
R1212 gnd.n640 gnd.n639 585
R1213 gnd.n6609 gnd.n6608 585
R1214 gnd.n6610 gnd.n6609 585
R1215 gnd.n638 gnd.n637 585
R1216 gnd.n6611 gnd.n638 585
R1217 gnd.n6614 gnd.n6613 585
R1218 gnd.n6613 gnd.n6612 585
R1219 gnd.n635 gnd.n634 585
R1220 gnd.n634 gnd.n633 585
R1221 gnd.n6619 gnd.n6618 585
R1222 gnd.n6620 gnd.n6619 585
R1223 gnd.n632 gnd.n631 585
R1224 gnd.n6621 gnd.n632 585
R1225 gnd.n6624 gnd.n6623 585
R1226 gnd.n6623 gnd.n6622 585
R1227 gnd.n629 gnd.n628 585
R1228 gnd.n628 gnd.n627 585
R1229 gnd.n6629 gnd.n6628 585
R1230 gnd.n6630 gnd.n6629 585
R1231 gnd.n626 gnd.n625 585
R1232 gnd.n6631 gnd.n626 585
R1233 gnd.n6634 gnd.n6633 585
R1234 gnd.n6633 gnd.n6632 585
R1235 gnd.n623 gnd.n622 585
R1236 gnd.n622 gnd.n621 585
R1237 gnd.n6639 gnd.n6638 585
R1238 gnd.n6640 gnd.n6639 585
R1239 gnd.n620 gnd.n619 585
R1240 gnd.n6641 gnd.n620 585
R1241 gnd.n6644 gnd.n6643 585
R1242 gnd.n6643 gnd.n6642 585
R1243 gnd.n617 gnd.n616 585
R1244 gnd.n616 gnd.n615 585
R1245 gnd.n6649 gnd.n6648 585
R1246 gnd.n6650 gnd.n6649 585
R1247 gnd.n614 gnd.n613 585
R1248 gnd.n6651 gnd.n614 585
R1249 gnd.n6654 gnd.n6653 585
R1250 gnd.n6653 gnd.n6652 585
R1251 gnd.n611 gnd.n610 585
R1252 gnd.n610 gnd.n609 585
R1253 gnd.n6659 gnd.n6658 585
R1254 gnd.n6660 gnd.n6659 585
R1255 gnd.n608 gnd.n607 585
R1256 gnd.n6661 gnd.n608 585
R1257 gnd.n6664 gnd.n6663 585
R1258 gnd.n6663 gnd.n6662 585
R1259 gnd.n605 gnd.n604 585
R1260 gnd.n604 gnd.n603 585
R1261 gnd.n6669 gnd.n6668 585
R1262 gnd.n6670 gnd.n6669 585
R1263 gnd.n602 gnd.n601 585
R1264 gnd.n6671 gnd.n602 585
R1265 gnd.n6674 gnd.n6673 585
R1266 gnd.n6673 gnd.n6672 585
R1267 gnd.n599 gnd.n598 585
R1268 gnd.n598 gnd.n597 585
R1269 gnd.n6679 gnd.n6678 585
R1270 gnd.n6680 gnd.n6679 585
R1271 gnd.n596 gnd.n595 585
R1272 gnd.n6681 gnd.n596 585
R1273 gnd.n6684 gnd.n6683 585
R1274 gnd.n6683 gnd.n6682 585
R1275 gnd.n593 gnd.n592 585
R1276 gnd.n592 gnd.n591 585
R1277 gnd.n6689 gnd.n6688 585
R1278 gnd.n6690 gnd.n6689 585
R1279 gnd.n590 gnd.n589 585
R1280 gnd.n6691 gnd.n590 585
R1281 gnd.n6694 gnd.n6693 585
R1282 gnd.n6693 gnd.n6692 585
R1283 gnd.n587 gnd.n586 585
R1284 gnd.n586 gnd.n585 585
R1285 gnd.n6699 gnd.n6698 585
R1286 gnd.n6700 gnd.n6699 585
R1287 gnd.n584 gnd.n583 585
R1288 gnd.n6701 gnd.n584 585
R1289 gnd.n6704 gnd.n6703 585
R1290 gnd.n6703 gnd.n6702 585
R1291 gnd.n581 gnd.n580 585
R1292 gnd.n580 gnd.n579 585
R1293 gnd.n6709 gnd.n6708 585
R1294 gnd.n6710 gnd.n6709 585
R1295 gnd.n578 gnd.n577 585
R1296 gnd.n6711 gnd.n578 585
R1297 gnd.n6714 gnd.n6713 585
R1298 gnd.n6713 gnd.n6712 585
R1299 gnd.n575 gnd.n574 585
R1300 gnd.n574 gnd.n573 585
R1301 gnd.n6719 gnd.n6718 585
R1302 gnd.n6720 gnd.n6719 585
R1303 gnd.n572 gnd.n571 585
R1304 gnd.n6721 gnd.n572 585
R1305 gnd.n6724 gnd.n6723 585
R1306 gnd.n6723 gnd.n6722 585
R1307 gnd.n569 gnd.n568 585
R1308 gnd.n568 gnd.n567 585
R1309 gnd.n6729 gnd.n6728 585
R1310 gnd.n6730 gnd.n6729 585
R1311 gnd.n566 gnd.n565 585
R1312 gnd.n6731 gnd.n566 585
R1313 gnd.n6734 gnd.n6733 585
R1314 gnd.n6733 gnd.n6732 585
R1315 gnd.n563 gnd.n562 585
R1316 gnd.n562 gnd.n561 585
R1317 gnd.n6739 gnd.n6738 585
R1318 gnd.n6740 gnd.n6739 585
R1319 gnd.n560 gnd.n559 585
R1320 gnd.n6741 gnd.n560 585
R1321 gnd.n6744 gnd.n6743 585
R1322 gnd.n6743 gnd.n6742 585
R1323 gnd.n557 gnd.n556 585
R1324 gnd.n556 gnd.n555 585
R1325 gnd.n6749 gnd.n6748 585
R1326 gnd.n6750 gnd.n6749 585
R1327 gnd.n554 gnd.n553 585
R1328 gnd.n6751 gnd.n554 585
R1329 gnd.n6754 gnd.n6753 585
R1330 gnd.n6753 gnd.n6752 585
R1331 gnd.n551 gnd.n550 585
R1332 gnd.n550 gnd.n549 585
R1333 gnd.n6759 gnd.n6758 585
R1334 gnd.n6760 gnd.n6759 585
R1335 gnd.n548 gnd.n547 585
R1336 gnd.n6761 gnd.n548 585
R1337 gnd.n6764 gnd.n6763 585
R1338 gnd.n6763 gnd.n6762 585
R1339 gnd.n545 gnd.n544 585
R1340 gnd.n544 gnd.n543 585
R1341 gnd.n6769 gnd.n6768 585
R1342 gnd.n6770 gnd.n6769 585
R1343 gnd.n542 gnd.n541 585
R1344 gnd.n6771 gnd.n542 585
R1345 gnd.n6774 gnd.n6773 585
R1346 gnd.n6773 gnd.n6772 585
R1347 gnd.n539 gnd.n538 585
R1348 gnd.n538 gnd.n537 585
R1349 gnd.n6779 gnd.n6778 585
R1350 gnd.n6780 gnd.n6779 585
R1351 gnd.n536 gnd.n535 585
R1352 gnd.n6781 gnd.n536 585
R1353 gnd.n6784 gnd.n6783 585
R1354 gnd.n6783 gnd.n6782 585
R1355 gnd.n533 gnd.n532 585
R1356 gnd.n532 gnd.n531 585
R1357 gnd.n6789 gnd.n6788 585
R1358 gnd.n6790 gnd.n6789 585
R1359 gnd.n530 gnd.n529 585
R1360 gnd.n6791 gnd.n530 585
R1361 gnd.n6794 gnd.n6793 585
R1362 gnd.n6793 gnd.n6792 585
R1363 gnd.n527 gnd.n526 585
R1364 gnd.n526 gnd.n525 585
R1365 gnd.n6799 gnd.n6798 585
R1366 gnd.n6800 gnd.n6799 585
R1367 gnd.n524 gnd.n523 585
R1368 gnd.n6801 gnd.n524 585
R1369 gnd.n6804 gnd.n6803 585
R1370 gnd.n6803 gnd.n6802 585
R1371 gnd.n521 gnd.n520 585
R1372 gnd.n520 gnd.n519 585
R1373 gnd.n6809 gnd.n6808 585
R1374 gnd.n6810 gnd.n6809 585
R1375 gnd.n518 gnd.n517 585
R1376 gnd.n6811 gnd.n518 585
R1377 gnd.n6814 gnd.n6813 585
R1378 gnd.n6813 gnd.n6812 585
R1379 gnd.n515 gnd.n514 585
R1380 gnd.n514 gnd.n513 585
R1381 gnd.n6819 gnd.n6818 585
R1382 gnd.n6820 gnd.n6819 585
R1383 gnd.n512 gnd.n511 585
R1384 gnd.n6821 gnd.n512 585
R1385 gnd.n6824 gnd.n6823 585
R1386 gnd.n6823 gnd.n6822 585
R1387 gnd.n509 gnd.n508 585
R1388 gnd.n508 gnd.n507 585
R1389 gnd.n6829 gnd.n6828 585
R1390 gnd.n6830 gnd.n6829 585
R1391 gnd.n506 gnd.n505 585
R1392 gnd.n6831 gnd.n506 585
R1393 gnd.n6834 gnd.n6833 585
R1394 gnd.n6833 gnd.n6832 585
R1395 gnd.n503 gnd.n502 585
R1396 gnd.n502 gnd.n501 585
R1397 gnd.n6839 gnd.n6838 585
R1398 gnd.n6840 gnd.n6839 585
R1399 gnd.n500 gnd.n499 585
R1400 gnd.n6841 gnd.n500 585
R1401 gnd.n6844 gnd.n6843 585
R1402 gnd.n6843 gnd.n6842 585
R1403 gnd.n497 gnd.n496 585
R1404 gnd.n496 gnd.n495 585
R1405 gnd.n6849 gnd.n6848 585
R1406 gnd.n6850 gnd.n6849 585
R1407 gnd.n494 gnd.n493 585
R1408 gnd.n6851 gnd.n494 585
R1409 gnd.n6854 gnd.n6853 585
R1410 gnd.n6853 gnd.n6852 585
R1411 gnd.n491 gnd.n490 585
R1412 gnd.n490 gnd.n489 585
R1413 gnd.n6859 gnd.n6858 585
R1414 gnd.n6860 gnd.n6859 585
R1415 gnd.n488 gnd.n487 585
R1416 gnd.n6861 gnd.n488 585
R1417 gnd.n6864 gnd.n6863 585
R1418 gnd.n6863 gnd.n6862 585
R1419 gnd.n485 gnd.n484 585
R1420 gnd.n484 gnd.n483 585
R1421 gnd.n6869 gnd.n6868 585
R1422 gnd.n6870 gnd.n6869 585
R1423 gnd.n482 gnd.n481 585
R1424 gnd.n6871 gnd.n482 585
R1425 gnd.n6874 gnd.n6873 585
R1426 gnd.n6873 gnd.n6872 585
R1427 gnd.n479 gnd.n478 585
R1428 gnd.n478 gnd.n477 585
R1429 gnd.n6879 gnd.n6878 585
R1430 gnd.n6880 gnd.n6879 585
R1431 gnd.n476 gnd.n475 585
R1432 gnd.n6881 gnd.n476 585
R1433 gnd.n6884 gnd.n6883 585
R1434 gnd.n6883 gnd.n6882 585
R1435 gnd.n473 gnd.n472 585
R1436 gnd.n472 gnd.n471 585
R1437 gnd.n6889 gnd.n6888 585
R1438 gnd.n6890 gnd.n6889 585
R1439 gnd.n470 gnd.n469 585
R1440 gnd.n6891 gnd.n470 585
R1441 gnd.n6894 gnd.n6893 585
R1442 gnd.n6893 gnd.n6892 585
R1443 gnd.n467 gnd.n466 585
R1444 gnd.n466 gnd.n465 585
R1445 gnd.n6899 gnd.n6898 585
R1446 gnd.n6900 gnd.n6899 585
R1447 gnd.n464 gnd.n463 585
R1448 gnd.n6901 gnd.n464 585
R1449 gnd.n6904 gnd.n6903 585
R1450 gnd.n6903 gnd.n6902 585
R1451 gnd.n461 gnd.n460 585
R1452 gnd.n460 gnd.n459 585
R1453 gnd.n6909 gnd.n6908 585
R1454 gnd.n6910 gnd.n6909 585
R1455 gnd.n458 gnd.n457 585
R1456 gnd.n6911 gnd.n458 585
R1457 gnd.n6914 gnd.n6913 585
R1458 gnd.n6913 gnd.n6912 585
R1459 gnd.n455 gnd.n454 585
R1460 gnd.n454 gnd.n453 585
R1461 gnd.n6919 gnd.n6918 585
R1462 gnd.n6920 gnd.n6919 585
R1463 gnd.n452 gnd.n451 585
R1464 gnd.n6921 gnd.n452 585
R1465 gnd.n6924 gnd.n6923 585
R1466 gnd.n6923 gnd.n6922 585
R1467 gnd.n449 gnd.n448 585
R1468 gnd.n448 gnd.n447 585
R1469 gnd.n6929 gnd.n6928 585
R1470 gnd.n6930 gnd.n6929 585
R1471 gnd.n446 gnd.n445 585
R1472 gnd.n6931 gnd.n446 585
R1473 gnd.n6934 gnd.n6933 585
R1474 gnd.n6933 gnd.n6932 585
R1475 gnd.n443 gnd.n442 585
R1476 gnd.n442 gnd.n441 585
R1477 gnd.n6939 gnd.n6938 585
R1478 gnd.n6940 gnd.n6939 585
R1479 gnd.n440 gnd.n439 585
R1480 gnd.n6941 gnd.n440 585
R1481 gnd.n6944 gnd.n6943 585
R1482 gnd.n6943 gnd.n6942 585
R1483 gnd.n437 gnd.n436 585
R1484 gnd.n436 gnd.n435 585
R1485 gnd.n6949 gnd.n6948 585
R1486 gnd.n6950 gnd.n6949 585
R1487 gnd.n434 gnd.n433 585
R1488 gnd.n6951 gnd.n434 585
R1489 gnd.n6954 gnd.n6953 585
R1490 gnd.n6953 gnd.n6952 585
R1491 gnd.n431 gnd.n430 585
R1492 gnd.n430 gnd.n429 585
R1493 gnd.n6959 gnd.n6958 585
R1494 gnd.n6960 gnd.n6959 585
R1495 gnd.n428 gnd.n427 585
R1496 gnd.n6961 gnd.n428 585
R1497 gnd.n6964 gnd.n6963 585
R1498 gnd.n6963 gnd.n6962 585
R1499 gnd.n425 gnd.n424 585
R1500 gnd.n424 gnd.n423 585
R1501 gnd.n6969 gnd.n6968 585
R1502 gnd.n6970 gnd.n6969 585
R1503 gnd.n422 gnd.n421 585
R1504 gnd.n6971 gnd.n422 585
R1505 gnd.n6974 gnd.n6973 585
R1506 gnd.n6973 gnd.n6972 585
R1507 gnd.n419 gnd.n418 585
R1508 gnd.n418 gnd.n417 585
R1509 gnd.n6979 gnd.n6978 585
R1510 gnd.n6980 gnd.n6979 585
R1511 gnd.n416 gnd.n415 585
R1512 gnd.n6981 gnd.n416 585
R1513 gnd.n6984 gnd.n6983 585
R1514 gnd.n6983 gnd.n6982 585
R1515 gnd.n413 gnd.n412 585
R1516 gnd.n412 gnd.n411 585
R1517 gnd.n6989 gnd.n6988 585
R1518 gnd.n6990 gnd.n6989 585
R1519 gnd.n410 gnd.n409 585
R1520 gnd.n6991 gnd.n410 585
R1521 gnd.n6994 gnd.n6993 585
R1522 gnd.n6993 gnd.n6992 585
R1523 gnd.n407 gnd.n406 585
R1524 gnd.n406 gnd.n405 585
R1525 gnd.n6999 gnd.n6998 585
R1526 gnd.n7000 gnd.n6999 585
R1527 gnd.n404 gnd.n403 585
R1528 gnd.n7001 gnd.n404 585
R1529 gnd.n7004 gnd.n7003 585
R1530 gnd.n7003 gnd.n7002 585
R1531 gnd.n401 gnd.n400 585
R1532 gnd.n400 gnd.n399 585
R1533 gnd.n7010 gnd.n7009 585
R1534 gnd.n7011 gnd.n7010 585
R1535 gnd.n398 gnd.n397 585
R1536 gnd.n7012 gnd.n398 585
R1537 gnd.n7015 gnd.n7014 585
R1538 gnd.n7014 gnd.n7013 585
R1539 gnd.n7016 gnd.n395 585
R1540 gnd.n395 gnd.n394 585
R1541 gnd.n270 gnd.n269 585
R1542 gnd.n269 gnd.n268 585
R1543 gnd.n7225 gnd.n7224 585
R1544 gnd.n7224 gnd.n7223 585
R1545 gnd.n273 gnd.n272 585
R1546 gnd.n7222 gnd.n273 585
R1547 gnd.n7220 gnd.n7219 585
R1548 gnd.n7221 gnd.n7220 585
R1549 gnd.n276 gnd.n275 585
R1550 gnd.n275 gnd.n274 585
R1551 gnd.n7215 gnd.n7214 585
R1552 gnd.n7214 gnd.n7213 585
R1553 gnd.n279 gnd.n278 585
R1554 gnd.n7212 gnd.n279 585
R1555 gnd.n7210 gnd.n7209 585
R1556 gnd.n7211 gnd.n7210 585
R1557 gnd.n282 gnd.n281 585
R1558 gnd.n281 gnd.n280 585
R1559 gnd.n7205 gnd.n7204 585
R1560 gnd.n7204 gnd.n7203 585
R1561 gnd.n285 gnd.n284 585
R1562 gnd.n7202 gnd.n285 585
R1563 gnd.n7200 gnd.n7199 585
R1564 gnd.n7201 gnd.n7200 585
R1565 gnd.n288 gnd.n287 585
R1566 gnd.n287 gnd.n286 585
R1567 gnd.n7195 gnd.n7194 585
R1568 gnd.n7194 gnd.n7193 585
R1569 gnd.n291 gnd.n290 585
R1570 gnd.n7192 gnd.n291 585
R1571 gnd.n7190 gnd.n7189 585
R1572 gnd.n7191 gnd.n7190 585
R1573 gnd.n294 gnd.n293 585
R1574 gnd.n293 gnd.n292 585
R1575 gnd.n7185 gnd.n7184 585
R1576 gnd.n7184 gnd.n7183 585
R1577 gnd.n297 gnd.n296 585
R1578 gnd.n7182 gnd.n297 585
R1579 gnd.n7180 gnd.n7179 585
R1580 gnd.n7181 gnd.n7180 585
R1581 gnd.n300 gnd.n299 585
R1582 gnd.n299 gnd.n298 585
R1583 gnd.n7175 gnd.n7174 585
R1584 gnd.n7174 gnd.n7173 585
R1585 gnd.n303 gnd.n302 585
R1586 gnd.n7172 gnd.n303 585
R1587 gnd.n7170 gnd.n7169 585
R1588 gnd.n7171 gnd.n7170 585
R1589 gnd.n306 gnd.n305 585
R1590 gnd.n305 gnd.n304 585
R1591 gnd.n7165 gnd.n7164 585
R1592 gnd.n7164 gnd.n7163 585
R1593 gnd.n309 gnd.n308 585
R1594 gnd.n7162 gnd.n309 585
R1595 gnd.n7160 gnd.n7159 585
R1596 gnd.n7161 gnd.n7160 585
R1597 gnd.n312 gnd.n311 585
R1598 gnd.n311 gnd.n310 585
R1599 gnd.n7155 gnd.n7154 585
R1600 gnd.n7154 gnd.n7153 585
R1601 gnd.n315 gnd.n314 585
R1602 gnd.n7152 gnd.n315 585
R1603 gnd.n7150 gnd.n7149 585
R1604 gnd.n7151 gnd.n7150 585
R1605 gnd.n318 gnd.n317 585
R1606 gnd.n317 gnd.n316 585
R1607 gnd.n7145 gnd.n7144 585
R1608 gnd.n7144 gnd.n7143 585
R1609 gnd.n321 gnd.n320 585
R1610 gnd.n7142 gnd.n321 585
R1611 gnd.n7140 gnd.n7139 585
R1612 gnd.n7141 gnd.n7140 585
R1613 gnd.n324 gnd.n323 585
R1614 gnd.n323 gnd.n322 585
R1615 gnd.n7135 gnd.n7134 585
R1616 gnd.n7134 gnd.n7133 585
R1617 gnd.n327 gnd.n326 585
R1618 gnd.n7132 gnd.n327 585
R1619 gnd.n7130 gnd.n7129 585
R1620 gnd.n7131 gnd.n7130 585
R1621 gnd.n330 gnd.n329 585
R1622 gnd.n329 gnd.n328 585
R1623 gnd.n7125 gnd.n7124 585
R1624 gnd.n7124 gnd.n7123 585
R1625 gnd.n333 gnd.n332 585
R1626 gnd.n7122 gnd.n333 585
R1627 gnd.n7120 gnd.n7119 585
R1628 gnd.n7121 gnd.n7120 585
R1629 gnd.n336 gnd.n335 585
R1630 gnd.n335 gnd.n334 585
R1631 gnd.n7115 gnd.n7114 585
R1632 gnd.n7114 gnd.n7113 585
R1633 gnd.n339 gnd.n338 585
R1634 gnd.n7112 gnd.n339 585
R1635 gnd.n7110 gnd.n7109 585
R1636 gnd.n7111 gnd.n7110 585
R1637 gnd.n342 gnd.n341 585
R1638 gnd.n341 gnd.n340 585
R1639 gnd.n7105 gnd.n7104 585
R1640 gnd.n7104 gnd.n7103 585
R1641 gnd.n345 gnd.n344 585
R1642 gnd.n7102 gnd.n345 585
R1643 gnd.n7100 gnd.n7099 585
R1644 gnd.n7101 gnd.n7100 585
R1645 gnd.n348 gnd.n347 585
R1646 gnd.n347 gnd.n346 585
R1647 gnd.n7095 gnd.n7094 585
R1648 gnd.n7094 gnd.n7093 585
R1649 gnd.n351 gnd.n350 585
R1650 gnd.n7092 gnd.n351 585
R1651 gnd.n7090 gnd.n7089 585
R1652 gnd.n7091 gnd.n7090 585
R1653 gnd.n354 gnd.n353 585
R1654 gnd.n353 gnd.n352 585
R1655 gnd.n7085 gnd.n7084 585
R1656 gnd.n7084 gnd.n7083 585
R1657 gnd.n357 gnd.n356 585
R1658 gnd.n7082 gnd.n357 585
R1659 gnd.n7080 gnd.n7079 585
R1660 gnd.n7081 gnd.n7080 585
R1661 gnd.n360 gnd.n359 585
R1662 gnd.n359 gnd.n358 585
R1663 gnd.n7075 gnd.n7074 585
R1664 gnd.n7074 gnd.n7073 585
R1665 gnd.n363 gnd.n362 585
R1666 gnd.n7072 gnd.n363 585
R1667 gnd.n7070 gnd.n7069 585
R1668 gnd.n7071 gnd.n7070 585
R1669 gnd.n366 gnd.n365 585
R1670 gnd.n365 gnd.n364 585
R1671 gnd.n7065 gnd.n7064 585
R1672 gnd.n7064 gnd.n7063 585
R1673 gnd.n369 gnd.n368 585
R1674 gnd.n7062 gnd.n369 585
R1675 gnd.n7060 gnd.n7059 585
R1676 gnd.n7061 gnd.n7060 585
R1677 gnd.n372 gnd.n371 585
R1678 gnd.n371 gnd.n370 585
R1679 gnd.n7055 gnd.n7054 585
R1680 gnd.n7054 gnd.n7053 585
R1681 gnd.n375 gnd.n374 585
R1682 gnd.n7052 gnd.n375 585
R1683 gnd.n7050 gnd.n7049 585
R1684 gnd.n7051 gnd.n7050 585
R1685 gnd.n378 gnd.n377 585
R1686 gnd.n377 gnd.n376 585
R1687 gnd.n7045 gnd.n7044 585
R1688 gnd.n7044 gnd.n7043 585
R1689 gnd.n381 gnd.n380 585
R1690 gnd.n7042 gnd.n381 585
R1691 gnd.n7040 gnd.n7039 585
R1692 gnd.n7041 gnd.n7040 585
R1693 gnd.n384 gnd.n383 585
R1694 gnd.n383 gnd.n382 585
R1695 gnd.n7035 gnd.n7034 585
R1696 gnd.n7034 gnd.n7033 585
R1697 gnd.n387 gnd.n386 585
R1698 gnd.n7032 gnd.n387 585
R1699 gnd.n7030 gnd.n7029 585
R1700 gnd.n7031 gnd.n7030 585
R1701 gnd.n390 gnd.n389 585
R1702 gnd.n389 gnd.n388 585
R1703 gnd.n7025 gnd.n7024 585
R1704 gnd.n7024 gnd.n7023 585
R1705 gnd.n393 gnd.n392 585
R1706 gnd.n7022 gnd.n393 585
R1707 gnd.n7020 gnd.n7019 585
R1708 gnd.n7021 gnd.n7020 585
R1709 gnd.n6166 gnd.n6165 585
R1710 gnd.n6167 gnd.n6166 585
R1711 gnd.n2560 gnd.n2559 585
R1712 gnd.n6160 gnd.n2560 585
R1713 gnd.n6175 gnd.n6174 585
R1714 gnd.n6174 gnd.n6173 585
R1715 gnd.n6176 gnd.n2555 585
R1716 gnd.n4314 gnd.n2555 585
R1717 gnd.n6178 gnd.n6177 585
R1718 gnd.n6179 gnd.n6178 585
R1719 gnd.n2540 gnd.n2539 585
R1720 gnd.n4308 gnd.n2540 585
R1721 gnd.n6187 gnd.n6186 585
R1722 gnd.n6186 gnd.n6185 585
R1723 gnd.n6188 gnd.n2535 585
R1724 gnd.n4303 gnd.n2535 585
R1725 gnd.n6190 gnd.n6189 585
R1726 gnd.n6191 gnd.n6190 585
R1727 gnd.n2519 gnd.n2518 585
R1728 gnd.n4298 gnd.n2519 585
R1729 gnd.n6199 gnd.n6198 585
R1730 gnd.n6198 gnd.n6197 585
R1731 gnd.n6200 gnd.n2514 585
R1732 gnd.n4331 gnd.n2514 585
R1733 gnd.n6202 gnd.n6201 585
R1734 gnd.n6203 gnd.n6202 585
R1735 gnd.n2500 gnd.n2499 585
R1736 gnd.n4291 gnd.n2500 585
R1737 gnd.n6211 gnd.n6210 585
R1738 gnd.n6210 gnd.n6209 585
R1739 gnd.n6212 gnd.n2495 585
R1740 gnd.n4283 gnd.n2495 585
R1741 gnd.n6214 gnd.n6213 585
R1742 gnd.n6215 gnd.n6214 585
R1743 gnd.n2482 gnd.n2481 585
R1744 gnd.n4251 gnd.n2482 585
R1745 gnd.n6224 gnd.n6223 585
R1746 gnd.n6223 gnd.n6222 585
R1747 gnd.n6225 gnd.n2477 585
R1748 gnd.n4242 gnd.n2477 585
R1749 gnd.n6227 gnd.n6226 585
R1750 gnd.n6228 gnd.n6227 585
R1751 gnd.n2466 gnd.n2465 585
R1752 gnd.n4227 gnd.n2466 585
R1753 gnd.n6237 gnd.n6236 585
R1754 gnd.n6236 gnd.n6235 585
R1755 gnd.n6238 gnd.n2461 585
R1756 gnd.n4264 gnd.n2461 585
R1757 gnd.n6240 gnd.n6239 585
R1758 gnd.n6241 gnd.n6240 585
R1759 gnd.n2447 gnd.n2446 585
R1760 gnd.n4220 gnd.n2447 585
R1761 gnd.n6250 gnd.n6249 585
R1762 gnd.n6249 gnd.n6248 585
R1763 gnd.n6251 gnd.n2442 585
R1764 gnd.n4211 gnd.n2442 585
R1765 gnd.n6253 gnd.n6252 585
R1766 gnd.n6254 gnd.n6253 585
R1767 gnd.n2427 gnd.n2426 585
R1768 gnd.n4205 gnd.n2427 585
R1769 gnd.n6262 gnd.n6261 585
R1770 gnd.n6261 gnd.n6260 585
R1771 gnd.n6263 gnd.n2422 585
R1772 gnd.n4197 gnd.n2422 585
R1773 gnd.n6265 gnd.n6264 585
R1774 gnd.n6266 gnd.n6265 585
R1775 gnd.n2406 gnd.n2405 585
R1776 gnd.n4142 gnd.n2406 585
R1777 gnd.n6274 gnd.n6273 585
R1778 gnd.n6273 gnd.n6272 585
R1779 gnd.n6275 gnd.n2401 585
R1780 gnd.n4148 gnd.n2401 585
R1781 gnd.n6277 gnd.n6276 585
R1782 gnd.n6278 gnd.n6277 585
R1783 gnd.n2385 gnd.n2384 585
R1784 gnd.n4154 gnd.n2385 585
R1785 gnd.n6286 gnd.n6285 585
R1786 gnd.n6285 gnd.n6284 585
R1787 gnd.n6287 gnd.n2379 585
R1788 gnd.n4160 gnd.n2379 585
R1789 gnd.n6289 gnd.n6288 585
R1790 gnd.n6290 gnd.n6289 585
R1791 gnd.n2380 gnd.n2378 585
R1792 gnd.n4166 gnd.n2378 585
R1793 gnd.n4123 gnd.n2367 585
R1794 gnd.n6296 gnd.n2367 585
R1795 gnd.n3908 gnd.n3907 585
R1796 gnd.n3905 gnd.n3842 585
R1797 gnd.n3904 gnd.n3903 585
R1798 gnd.n3902 gnd.n3901 585
R1799 gnd.n3900 gnd.n3846 585
R1800 gnd.n3898 gnd.n3897 585
R1801 gnd.n3896 gnd.n3847 585
R1802 gnd.n3895 gnd.n3894 585
R1803 gnd.n3892 gnd.n3852 585
R1804 gnd.n3890 gnd.n3889 585
R1805 gnd.n3888 gnd.n3853 585
R1806 gnd.n3887 gnd.n3886 585
R1807 gnd.n3884 gnd.n3858 585
R1808 gnd.n3882 gnd.n3881 585
R1809 gnd.n3880 gnd.n3859 585
R1810 gnd.n3879 gnd.n3878 585
R1811 gnd.n3876 gnd.n3864 585
R1812 gnd.n3874 gnd.n3873 585
R1813 gnd.n3866 gnd.n3865 585
R1814 gnd.n3865 gnd.n2363 585
R1815 gnd.n6087 gnd.n6086 585
R1816 gnd.n6088 gnd.n2675 585
R1817 gnd.n6089 gnd.n2670 585
R1818 gnd.n2688 gnd.n2659 585
R1819 gnd.n6096 gnd.n2658 585
R1820 gnd.n6097 gnd.n2657 585
R1821 gnd.n2685 gnd.n2651 585
R1822 gnd.n6104 gnd.n2650 585
R1823 gnd.n6105 gnd.n2649 585
R1824 gnd.n2683 gnd.n2641 585
R1825 gnd.n6112 gnd.n2640 585
R1826 gnd.n6113 gnd.n2639 585
R1827 gnd.n2680 gnd.n2633 585
R1828 gnd.n6120 gnd.n2632 585
R1829 gnd.n6121 gnd.n2631 585
R1830 gnd.n2678 gnd.n2623 585
R1831 gnd.n6128 gnd.n2622 585
R1832 gnd.n6129 gnd.n2621 585
R1833 gnd.n2620 gnd.n2575 585
R1834 gnd.n6084 gnd.n2575 585
R1835 gnd.n2580 gnd.n2573 585
R1836 gnd.n6167 gnd.n2573 585
R1837 gnd.n6159 gnd.n6158 585
R1838 gnd.n6160 gnd.n6159 585
R1839 gnd.n2579 gnd.n2563 585
R1840 gnd.n6173 gnd.n2563 585
R1841 gnd.n4317 gnd.n4315 585
R1842 gnd.n4315 gnd.n4314 585
R1843 gnd.n4318 gnd.n2553 585
R1844 gnd.n6179 gnd.n2553 585
R1845 gnd.n4319 gnd.n3778 585
R1846 gnd.n4308 gnd.n3778 585
R1847 gnd.n3776 gnd.n2542 585
R1848 gnd.n6185 gnd.n2542 585
R1849 gnd.n4323 gnd.n3775 585
R1850 gnd.n4303 gnd.n3775 585
R1851 gnd.n4324 gnd.n2533 585
R1852 gnd.n6191 gnd.n2533 585
R1853 gnd.n4325 gnd.n3774 585
R1854 gnd.n4298 gnd.n3774 585
R1855 gnd.n3771 gnd.n2522 585
R1856 gnd.n6197 gnd.n2522 585
R1857 gnd.n4330 gnd.n4329 585
R1858 gnd.n4331 gnd.n4330 585
R1859 gnd.n3770 gnd.n2513 585
R1860 gnd.n6203 gnd.n2513 585
R1861 gnd.n4290 gnd.n4289 585
R1862 gnd.n4291 gnd.n4290 585
R1863 gnd.n3781 gnd.n2502 585
R1864 gnd.n6209 gnd.n2502 585
R1865 gnd.n4285 gnd.n4284 585
R1866 gnd.n4284 gnd.n4283 585
R1867 gnd.n3783 gnd.n2493 585
R1868 gnd.n6215 gnd.n2493 585
R1869 gnd.n4254 gnd.n4252 585
R1870 gnd.n4252 gnd.n4251 585
R1871 gnd.n4255 gnd.n2485 585
R1872 gnd.n6222 gnd.n2485 585
R1873 gnd.n4256 gnd.n3807 585
R1874 gnd.n4242 gnd.n3807 585
R1875 gnd.n3805 gnd.n2476 585
R1876 gnd.n6228 gnd.n2476 585
R1877 gnd.n4260 gnd.n3804 585
R1878 gnd.n4227 gnd.n3804 585
R1879 gnd.n4261 gnd.n2468 585
R1880 gnd.n6235 gnd.n2468 585
R1881 gnd.n4263 gnd.n4262 585
R1882 gnd.n4264 gnd.n4263 585
R1883 gnd.n3801 gnd.n2459 585
R1884 gnd.n6241 gnd.n2459 585
R1885 gnd.n4219 gnd.n4218 585
R1886 gnd.n4220 gnd.n4219 585
R1887 gnd.n3810 gnd.n2450 585
R1888 gnd.n6248 gnd.n2450 585
R1889 gnd.n4213 gnd.n4212 585
R1890 gnd.n4212 gnd.n4211 585
R1891 gnd.n3812 gnd.n2440 585
R1892 gnd.n6254 gnd.n2440 585
R1893 gnd.n4204 gnd.n4203 585
R1894 gnd.n4205 gnd.n4204 585
R1895 gnd.n3815 gnd.n2429 585
R1896 gnd.n6260 gnd.n2429 585
R1897 gnd.n4199 gnd.n4198 585
R1898 gnd.n4198 gnd.n4197 585
R1899 gnd.n3817 gnd.n2420 585
R1900 gnd.n6266 gnd.n2420 585
R1901 gnd.n4141 gnd.n4140 585
R1902 gnd.n4142 gnd.n4141 585
R1903 gnd.n4134 gnd.n2409 585
R1904 gnd.n6272 gnd.n2409 585
R1905 gnd.n4150 gnd.n4149 585
R1906 gnd.n4149 gnd.n4148 585
R1907 gnd.n4151 gnd.n2399 585
R1908 gnd.n6278 gnd.n2399 585
R1909 gnd.n4153 gnd.n4152 585
R1910 gnd.n4154 gnd.n4153 585
R1911 gnd.n3839 gnd.n2388 585
R1912 gnd.n6284 gnd.n2388 585
R1913 gnd.n4162 gnd.n4161 585
R1914 gnd.n4161 gnd.n4160 585
R1915 gnd.n4163 gnd.n2376 585
R1916 gnd.n6290 gnd.n2376 585
R1917 gnd.n4165 gnd.n4164 585
R1918 gnd.n4166 gnd.n4165 585
R1919 gnd.n3835 gnd.n2365 585
R1920 gnd.n6296 gnd.n2365 585
R1921 gnd.n2246 gnd.n2245 585
R1922 gnd.n2247 gnd.n2246 585
R1923 gnd.n953 gnd.n952 585
R1924 gnd.n959 gnd.n952 585
R1925 gnd.n2221 gnd.n971 585
R1926 gnd.n971 gnd.n958 585
R1927 gnd.n2223 gnd.n2222 585
R1928 gnd.n2224 gnd.n2223 585
R1929 gnd.n972 gnd.n970 585
R1930 gnd.n970 gnd.n966 585
R1931 gnd.n1955 gnd.n1954 585
R1932 gnd.n1954 gnd.n1953 585
R1933 gnd.n977 gnd.n976 585
R1934 gnd.n1924 gnd.n977 585
R1935 gnd.n1944 gnd.n1943 585
R1936 gnd.n1943 gnd.n1942 585
R1937 gnd.n984 gnd.n983 585
R1938 gnd.n1930 gnd.n984 585
R1939 gnd.n1900 gnd.n1004 585
R1940 gnd.n1004 gnd.n1003 585
R1941 gnd.n1902 gnd.n1901 585
R1942 gnd.n1903 gnd.n1902 585
R1943 gnd.n1005 gnd.n1002 585
R1944 gnd.n1013 gnd.n1002 585
R1945 gnd.n1878 gnd.n1025 585
R1946 gnd.n1025 gnd.n1012 585
R1947 gnd.n1880 gnd.n1879 585
R1948 gnd.n1881 gnd.n1880 585
R1949 gnd.n1026 gnd.n1024 585
R1950 gnd.n1024 gnd.n1020 585
R1951 gnd.n1866 gnd.n1865 585
R1952 gnd.n1865 gnd.n1864 585
R1953 gnd.n1031 gnd.n1030 585
R1954 gnd.n1040 gnd.n1031 585
R1955 gnd.n1855 gnd.n1854 585
R1956 gnd.n1854 gnd.n1853 585
R1957 gnd.n1038 gnd.n1037 585
R1958 gnd.n1841 gnd.n1038 585
R1959 gnd.n1813 gnd.n1057 585
R1960 gnd.n1057 gnd.n1047 585
R1961 gnd.n1815 gnd.n1814 585
R1962 gnd.n1816 gnd.n1815 585
R1963 gnd.n1058 gnd.n1056 585
R1964 gnd.n1066 gnd.n1056 585
R1965 gnd.n1791 gnd.n1078 585
R1966 gnd.n1078 gnd.n1065 585
R1967 gnd.n1793 gnd.n1792 585
R1968 gnd.n1794 gnd.n1793 585
R1969 gnd.n1079 gnd.n1077 585
R1970 gnd.n1077 gnd.n1073 585
R1971 gnd.n1779 gnd.n1778 585
R1972 gnd.n1778 gnd.n1777 585
R1973 gnd.n1084 gnd.n1083 585
R1974 gnd.n1093 gnd.n1084 585
R1975 gnd.n1768 gnd.n1767 585
R1976 gnd.n1767 gnd.n1766 585
R1977 gnd.n1091 gnd.n1090 585
R1978 gnd.n1754 gnd.n1091 585
R1979 gnd.n1192 gnd.n1191 585
R1980 gnd.n1192 gnd.n1100 585
R1981 gnd.n1711 gnd.n1710 585
R1982 gnd.n1710 gnd.n1709 585
R1983 gnd.n1712 gnd.n1186 585
R1984 gnd.n1197 gnd.n1186 585
R1985 gnd.n1714 gnd.n1713 585
R1986 gnd.n1715 gnd.n1714 585
R1987 gnd.n1187 gnd.n1185 585
R1988 gnd.n1210 gnd.n1185 585
R1989 gnd.n1170 gnd.n1169 585
R1990 gnd.n1173 gnd.n1170 585
R1991 gnd.n1725 gnd.n1724 585
R1992 gnd.n1724 gnd.n1723 585
R1993 gnd.n1726 gnd.n1164 585
R1994 gnd.n1685 gnd.n1164 585
R1995 gnd.n1728 gnd.n1727 585
R1996 gnd.n1729 gnd.n1728 585
R1997 gnd.n1165 gnd.n1163 585
R1998 gnd.n1224 gnd.n1163 585
R1999 gnd.n1677 gnd.n1676 585
R2000 gnd.n1676 gnd.n1675 585
R2001 gnd.n1221 gnd.n1220 585
R2002 gnd.n1659 gnd.n1221 585
R2003 gnd.n1646 gnd.n1240 585
R2004 gnd.n1240 gnd.n1239 585
R2005 gnd.n1648 gnd.n1647 585
R2006 gnd.n1649 gnd.n1648 585
R2007 gnd.n1241 gnd.n1238 585
R2008 gnd.n1247 gnd.n1238 585
R2009 gnd.n1627 gnd.n1626 585
R2010 gnd.n1628 gnd.n1627 585
R2011 gnd.n1258 gnd.n1257 585
R2012 gnd.n1257 gnd.n1253 585
R2013 gnd.n1617 gnd.n1616 585
R2014 gnd.n1618 gnd.n1617 585
R2015 gnd.n1268 gnd.n1267 585
R2016 gnd.n1273 gnd.n1267 585
R2017 gnd.n1595 gnd.n1286 585
R2018 gnd.n1286 gnd.n1272 585
R2019 gnd.n1597 gnd.n1596 585
R2020 gnd.n1598 gnd.n1597 585
R2021 gnd.n1287 gnd.n1285 585
R2022 gnd.n1285 gnd.n1281 585
R2023 gnd.n1586 gnd.n1585 585
R2024 gnd.n1587 gnd.n1586 585
R2025 gnd.n1294 gnd.n1293 585
R2026 gnd.n1298 gnd.n1293 585
R2027 gnd.n1563 gnd.n1315 585
R2028 gnd.n1315 gnd.n1297 585
R2029 gnd.n1565 gnd.n1564 585
R2030 gnd.n1566 gnd.n1565 585
R2031 gnd.n1316 gnd.n1314 585
R2032 gnd.n1314 gnd.n1305 585
R2033 gnd.n1558 gnd.n1557 585
R2034 gnd.n1557 gnd.n1556 585
R2035 gnd.n1363 gnd.n1362 585
R2036 gnd.n1364 gnd.n1363 585
R2037 gnd.n1517 gnd.n1516 585
R2038 gnd.n1518 gnd.n1517 585
R2039 gnd.n1373 gnd.n1372 585
R2040 gnd.n1372 gnd.n1371 585
R2041 gnd.n1512 gnd.n1511 585
R2042 gnd.n1511 gnd.n1510 585
R2043 gnd.n1376 gnd.n1375 585
R2044 gnd.n1377 gnd.n1376 585
R2045 gnd.n1501 gnd.n1500 585
R2046 gnd.n1502 gnd.n1501 585
R2047 gnd.n1384 gnd.n1383 585
R2048 gnd.n1493 gnd.n1383 585
R2049 gnd.n1496 gnd.n1495 585
R2050 gnd.n1495 gnd.n1494 585
R2051 gnd.n1387 gnd.n1386 585
R2052 gnd.n1388 gnd.n1387 585
R2053 gnd.n1482 gnd.n1481 585
R2054 gnd.n1480 gnd.n1406 585
R2055 gnd.n1479 gnd.n1405 585
R2056 gnd.n1484 gnd.n1405 585
R2057 gnd.n1478 gnd.n1477 585
R2058 gnd.n1476 gnd.n1475 585
R2059 gnd.n1474 gnd.n1473 585
R2060 gnd.n1472 gnd.n1471 585
R2061 gnd.n1470 gnd.n1469 585
R2062 gnd.n1468 gnd.n1467 585
R2063 gnd.n1466 gnd.n1465 585
R2064 gnd.n1464 gnd.n1463 585
R2065 gnd.n1462 gnd.n1461 585
R2066 gnd.n1460 gnd.n1459 585
R2067 gnd.n1458 gnd.n1457 585
R2068 gnd.n1456 gnd.n1455 585
R2069 gnd.n1454 gnd.n1453 585
R2070 gnd.n1452 gnd.n1451 585
R2071 gnd.n1450 gnd.n1449 585
R2072 gnd.n1448 gnd.n1447 585
R2073 gnd.n1446 gnd.n1445 585
R2074 gnd.n1444 gnd.n1443 585
R2075 gnd.n1442 gnd.n1441 585
R2076 gnd.n1440 gnd.n1439 585
R2077 gnd.n1438 gnd.n1437 585
R2078 gnd.n1436 gnd.n1435 585
R2079 gnd.n1393 gnd.n1392 585
R2080 gnd.n1487 gnd.n1486 585
R2081 gnd.n2250 gnd.n2249 585
R2082 gnd.n2252 gnd.n2251 585
R2083 gnd.n2254 gnd.n2253 585
R2084 gnd.n2256 gnd.n2255 585
R2085 gnd.n2258 gnd.n2257 585
R2086 gnd.n2260 gnd.n2259 585
R2087 gnd.n2262 gnd.n2261 585
R2088 gnd.n2264 gnd.n2263 585
R2089 gnd.n2266 gnd.n2265 585
R2090 gnd.n2268 gnd.n2267 585
R2091 gnd.n2270 gnd.n2269 585
R2092 gnd.n2272 gnd.n2271 585
R2093 gnd.n2274 gnd.n2273 585
R2094 gnd.n2276 gnd.n2275 585
R2095 gnd.n2278 gnd.n2277 585
R2096 gnd.n2280 gnd.n2279 585
R2097 gnd.n2282 gnd.n2281 585
R2098 gnd.n2284 gnd.n2283 585
R2099 gnd.n2286 gnd.n2285 585
R2100 gnd.n2288 gnd.n2287 585
R2101 gnd.n2290 gnd.n2289 585
R2102 gnd.n2292 gnd.n2291 585
R2103 gnd.n2294 gnd.n2293 585
R2104 gnd.n2296 gnd.n2295 585
R2105 gnd.n2298 gnd.n2297 585
R2106 gnd.n2299 gnd.n920 585
R2107 gnd.n2300 gnd.n878 585
R2108 gnd.n2338 gnd.n878 585
R2109 gnd.n2248 gnd.n950 585
R2110 gnd.n2248 gnd.n2247 585
R2111 gnd.n1917 gnd.n949 585
R2112 gnd.n959 gnd.n949 585
R2113 gnd.n1919 gnd.n1918 585
R2114 gnd.n1918 gnd.n958 585
R2115 gnd.n1920 gnd.n968 585
R2116 gnd.n2224 gnd.n968 585
R2117 gnd.n1922 gnd.n1921 585
R2118 gnd.n1921 gnd.n966 585
R2119 gnd.n1923 gnd.n979 585
R2120 gnd.n1953 gnd.n979 585
R2121 gnd.n1926 gnd.n1925 585
R2122 gnd.n1925 gnd.n1924 585
R2123 gnd.n1927 gnd.n986 585
R2124 gnd.n1942 gnd.n986 585
R2125 gnd.n1929 gnd.n1928 585
R2126 gnd.n1930 gnd.n1929 585
R2127 gnd.n996 gnd.n995 585
R2128 gnd.n1003 gnd.n995 585
R2129 gnd.n1905 gnd.n1904 585
R2130 gnd.n1904 gnd.n1903 585
R2131 gnd.n999 gnd.n998 585
R2132 gnd.n1013 gnd.n999 585
R2133 gnd.n1829 gnd.n1828 585
R2134 gnd.n1828 gnd.n1012 585
R2135 gnd.n1830 gnd.n1022 585
R2136 gnd.n1881 gnd.n1022 585
R2137 gnd.n1832 gnd.n1831 585
R2138 gnd.n1831 gnd.n1020 585
R2139 gnd.n1833 gnd.n1033 585
R2140 gnd.n1864 gnd.n1033 585
R2141 gnd.n1835 gnd.n1834 585
R2142 gnd.n1834 gnd.n1040 585
R2143 gnd.n1836 gnd.n1039 585
R2144 gnd.n1853 gnd.n1039 585
R2145 gnd.n1838 gnd.n1837 585
R2146 gnd.n1841 gnd.n1838 585
R2147 gnd.n1050 gnd.n1049 585
R2148 gnd.n1049 gnd.n1047 585
R2149 gnd.n1818 gnd.n1817 585
R2150 gnd.n1817 gnd.n1816 585
R2151 gnd.n1053 gnd.n1052 585
R2152 gnd.n1066 gnd.n1053 585
R2153 gnd.n1742 gnd.n1741 585
R2154 gnd.n1741 gnd.n1065 585
R2155 gnd.n1743 gnd.n1075 585
R2156 gnd.n1794 gnd.n1075 585
R2157 gnd.n1745 gnd.n1744 585
R2158 gnd.n1744 gnd.n1073 585
R2159 gnd.n1746 gnd.n1086 585
R2160 gnd.n1777 gnd.n1086 585
R2161 gnd.n1748 gnd.n1747 585
R2162 gnd.n1747 gnd.n1093 585
R2163 gnd.n1749 gnd.n1092 585
R2164 gnd.n1766 gnd.n1092 585
R2165 gnd.n1751 gnd.n1750 585
R2166 gnd.n1754 gnd.n1751 585
R2167 gnd.n1103 gnd.n1102 585
R2168 gnd.n1102 gnd.n1100 585
R2169 gnd.n1194 gnd.n1193 585
R2170 gnd.n1709 gnd.n1193 585
R2171 gnd.n1196 gnd.n1195 585
R2172 gnd.n1197 gnd.n1196 585
R2173 gnd.n1207 gnd.n1183 585
R2174 gnd.n1715 gnd.n1183 585
R2175 gnd.n1209 gnd.n1208 585
R2176 gnd.n1210 gnd.n1209 585
R2177 gnd.n1206 gnd.n1205 585
R2178 gnd.n1206 gnd.n1173 585
R2179 gnd.n1204 gnd.n1171 585
R2180 gnd.n1723 gnd.n1171 585
R2181 gnd.n1160 gnd.n1158 585
R2182 gnd.n1685 gnd.n1160 585
R2183 gnd.n1731 gnd.n1730 585
R2184 gnd.n1730 gnd.n1729 585
R2185 gnd.n1159 gnd.n1157 585
R2186 gnd.n1224 gnd.n1159 585
R2187 gnd.n1656 gnd.n1223 585
R2188 gnd.n1675 gnd.n1223 585
R2189 gnd.n1658 gnd.n1657 585
R2190 gnd.n1659 gnd.n1658 585
R2191 gnd.n1233 gnd.n1232 585
R2192 gnd.n1239 gnd.n1232 585
R2193 gnd.n1651 gnd.n1650 585
R2194 gnd.n1650 gnd.n1649 585
R2195 gnd.n1236 gnd.n1235 585
R2196 gnd.n1247 gnd.n1236 585
R2197 gnd.n1536 gnd.n1255 585
R2198 gnd.n1628 gnd.n1255 585
R2199 gnd.n1538 gnd.n1537 585
R2200 gnd.n1537 gnd.n1253 585
R2201 gnd.n1539 gnd.n1266 585
R2202 gnd.n1618 gnd.n1266 585
R2203 gnd.n1541 gnd.n1540 585
R2204 gnd.n1541 gnd.n1273 585
R2205 gnd.n1543 gnd.n1542 585
R2206 gnd.n1542 gnd.n1272 585
R2207 gnd.n1544 gnd.n1283 585
R2208 gnd.n1598 gnd.n1283 585
R2209 gnd.n1546 gnd.n1545 585
R2210 gnd.n1545 gnd.n1281 585
R2211 gnd.n1547 gnd.n1292 585
R2212 gnd.n1587 gnd.n1292 585
R2213 gnd.n1549 gnd.n1548 585
R2214 gnd.n1549 gnd.n1298 585
R2215 gnd.n1551 gnd.n1550 585
R2216 gnd.n1550 gnd.n1297 585
R2217 gnd.n1552 gnd.n1313 585
R2218 gnd.n1566 gnd.n1313 585
R2219 gnd.n1553 gnd.n1366 585
R2220 gnd.n1366 gnd.n1305 585
R2221 gnd.n1555 gnd.n1554 585
R2222 gnd.n1556 gnd.n1555 585
R2223 gnd.n1367 gnd.n1365 585
R2224 gnd.n1365 gnd.n1364 585
R2225 gnd.n1520 gnd.n1519 585
R2226 gnd.n1519 gnd.n1518 585
R2227 gnd.n1370 gnd.n1369 585
R2228 gnd.n1371 gnd.n1370 585
R2229 gnd.n1509 gnd.n1508 585
R2230 gnd.n1510 gnd.n1509 585
R2231 gnd.n1379 gnd.n1378 585
R2232 gnd.n1378 gnd.n1377 585
R2233 gnd.n1504 gnd.n1503 585
R2234 gnd.n1503 gnd.n1502 585
R2235 gnd.n1382 gnd.n1381 585
R2236 gnd.n1493 gnd.n1382 585
R2237 gnd.n1492 gnd.n1491 585
R2238 gnd.n1494 gnd.n1492 585
R2239 gnd.n1390 gnd.n1389 585
R2240 gnd.n1389 gnd.n1388 585
R2241 gnd.n7484 gnd.n7483 585
R2242 gnd.n7485 gnd.n7484 585
R2243 gnd.n158 gnd.n157 585
R2244 gnd.n7478 gnd.n158 585
R2245 gnd.n7493 gnd.n7492 585
R2246 gnd.n7492 gnd.n7491 585
R2247 gnd.n7494 gnd.n153 585
R2248 gnd.n5731 gnd.n153 585
R2249 gnd.n7496 gnd.n7495 585
R2250 gnd.n7497 gnd.n7496 585
R2251 gnd.n137 gnd.n136 585
R2252 gnd.n5737 gnd.n137 585
R2253 gnd.n7505 gnd.n7504 585
R2254 gnd.n7504 gnd.n7503 585
R2255 gnd.n7506 gnd.n132 585
R2256 gnd.n5743 gnd.n132 585
R2257 gnd.n7508 gnd.n7507 585
R2258 gnd.n7509 gnd.n7508 585
R2259 gnd.n116 gnd.n115 585
R2260 gnd.n5749 gnd.n116 585
R2261 gnd.n7517 gnd.n7516 585
R2262 gnd.n7516 gnd.n7515 585
R2263 gnd.n7518 gnd.n111 585
R2264 gnd.n5755 gnd.n111 585
R2265 gnd.n7520 gnd.n7519 585
R2266 gnd.n7521 gnd.n7520 585
R2267 gnd.n97 gnd.n96 585
R2268 gnd.n5712 gnd.n97 585
R2269 gnd.n7529 gnd.n7528 585
R2270 gnd.n7528 gnd.n7527 585
R2271 gnd.n7530 gnd.n91 585
R2272 gnd.n5703 gnd.n91 585
R2273 gnd.n7532 gnd.n7531 585
R2274 gnd.n7533 gnd.n7532 585
R2275 gnd.n92 gnd.n90 585
R2276 gnd.n5697 gnd.n90 585
R2277 gnd.n5772 gnd.n5771 585
R2278 gnd.n5771 gnd.n5770 585
R2279 gnd.n5773 gnd.n72 585
R2280 gnd.n7541 gnd.n72 585
R2281 gnd.n5774 gnd.n3131 585
R2282 gnd.n5687 gnd.n3131 585
R2283 gnd.n5776 gnd.n5775 585
R2284 gnd.n5777 gnd.n5776 585
R2285 gnd.n3132 gnd.n3124 585
R2286 gnd.n5782 gnd.n3124 585
R2287 gnd.n5682 gnd.n5681 585
R2288 gnd.n5681 gnd.n3120 585
R2289 gnd.n5680 gnd.n5679 585
R2290 gnd.n5680 gnd.n3113 585
R2291 gnd.n3103 gnd.n3102 585
R2292 gnd.n5791 gnd.n3103 585
R2293 gnd.n5797 gnd.n5796 585
R2294 gnd.n5796 gnd.n5795 585
R2295 gnd.n5798 gnd.n3098 585
R2296 gnd.n5670 gnd.n3098 585
R2297 gnd.n5800 gnd.n5799 585
R2298 gnd.n5801 gnd.n5800 585
R2299 gnd.n3084 gnd.n3083 585
R2300 gnd.n5652 gnd.n3084 585
R2301 gnd.n5809 gnd.n5808 585
R2302 gnd.n5808 gnd.n5807 585
R2303 gnd.n5810 gnd.n3079 585
R2304 gnd.n5645 gnd.n3079 585
R2305 gnd.n5812 gnd.n5811 585
R2306 gnd.n5813 gnd.n5812 585
R2307 gnd.n3063 gnd.n3062 585
R2308 gnd.n5589 gnd.n3063 585
R2309 gnd.n5821 gnd.n5820 585
R2310 gnd.n5820 gnd.n5819 585
R2311 gnd.n5822 gnd.n3058 585
R2312 gnd.n5600 gnd.n3058 585
R2313 gnd.n5824 gnd.n5823 585
R2314 gnd.n5825 gnd.n5824 585
R2315 gnd.n3043 gnd.n3042 585
R2316 gnd.n5580 gnd.n3043 585
R2317 gnd.n5833 gnd.n5832 585
R2318 gnd.n5832 gnd.n5831 585
R2319 gnd.n5834 gnd.n3037 585
R2320 gnd.n5572 gnd.n3037 585
R2321 gnd.n5836 gnd.n5835 585
R2322 gnd.n5837 gnd.n5836 585
R2323 gnd.n3038 gnd.n3036 585
R2324 gnd.n4993 gnd.n3036 585
R2325 gnd.n5565 gnd.n3024 585
R2326 gnd.n5843 gnd.n3024 585
R2327 gnd.n5080 gnd.n5079 585
R2328 gnd.n5043 gnd.n5042 585
R2329 gnd.n5094 gnd.n5093 585
R2330 gnd.n5096 gnd.n5041 585
R2331 gnd.n5099 gnd.n5098 585
R2332 gnd.n5034 gnd.n5033 585
R2333 gnd.n5113 gnd.n5112 585
R2334 gnd.n5115 gnd.n5032 585
R2335 gnd.n5118 gnd.n5117 585
R2336 gnd.n5025 gnd.n5024 585
R2337 gnd.n5132 gnd.n5131 585
R2338 gnd.n5134 gnd.n5023 585
R2339 gnd.n5137 gnd.n5136 585
R2340 gnd.n5016 gnd.n5015 585
R2341 gnd.n5152 gnd.n5151 585
R2342 gnd.n5154 gnd.n5014 585
R2343 gnd.n5157 gnd.n5156 585
R2344 gnd.n5158 gnd.n5011 585
R2345 gnd.n5010 gnd.n5009 585
R2346 gnd.n5010 gnd.n3012 585
R2347 gnd.n7472 gnd.n7471 585
R2348 gnd.n183 gnd.n182 585
R2349 gnd.n241 gnd.n240 585
R2350 gnd.n193 gnd.n192 585
R2351 gnd.n236 gnd.n235 585
R2352 gnd.n234 gnd.n233 585
R2353 gnd.n232 gnd.n231 585
R2354 gnd.n225 gnd.n195 585
R2355 gnd.n227 gnd.n226 585
R2356 gnd.n224 gnd.n223 585
R2357 gnd.n222 gnd.n221 585
R2358 gnd.n215 gnd.n197 585
R2359 gnd.n217 gnd.n216 585
R2360 gnd.n214 gnd.n213 585
R2361 gnd.n212 gnd.n211 585
R2362 gnd.n205 gnd.n199 585
R2363 gnd.n207 gnd.n206 585
R2364 gnd.n204 gnd.n203 585
R2365 gnd.n202 gnd.n172 585
R2366 gnd.n7469 gnd.n172 585
R2367 gnd.n7475 gnd.n170 585
R2368 gnd.n7485 gnd.n170 585
R2369 gnd.n7477 gnd.n7476 585
R2370 gnd.n7478 gnd.n7477 585
R2371 gnd.n177 gnd.n161 585
R2372 gnd.n7491 gnd.n161 585
R2373 gnd.n5730 gnd.n5729 585
R2374 gnd.n5731 gnd.n5730 585
R2375 gnd.n5724 gnd.n151 585
R2376 gnd.n7497 gnd.n151 585
R2377 gnd.n5739 gnd.n5738 585
R2378 gnd.n5738 gnd.n5737 585
R2379 gnd.n5740 gnd.n140 585
R2380 gnd.n7503 gnd.n140 585
R2381 gnd.n5742 gnd.n5741 585
R2382 gnd.n5743 gnd.n5742 585
R2383 gnd.n3196 gnd.n130 585
R2384 gnd.n7509 gnd.n130 585
R2385 gnd.n5751 gnd.n5750 585
R2386 gnd.n5750 gnd.n5749 585
R2387 gnd.n5752 gnd.n119 585
R2388 gnd.n7515 gnd.n119 585
R2389 gnd.n5754 gnd.n5753 585
R2390 gnd.n5755 gnd.n5754 585
R2391 gnd.n3192 gnd.n110 585
R2392 gnd.n7521 gnd.n110 585
R2393 gnd.n5711 gnd.n5710 585
R2394 gnd.n5712 gnd.n5711 585
R2395 gnd.n3199 gnd.n100 585
R2396 gnd.n7527 gnd.n100 585
R2397 gnd.n5705 gnd.n5704 585
R2398 gnd.n5704 gnd.n5703 585
R2399 gnd.n3201 gnd.n88 585
R2400 gnd.n7533 gnd.n88 585
R2401 gnd.n5696 gnd.n5695 585
R2402 gnd.n5697 gnd.n5696 585
R2403 gnd.n68 gnd.n67 585
R2404 gnd.n5770 gnd.n68 585
R2405 gnd.n7543 gnd.n7542 585
R2406 gnd.n7542 gnd.n7541 585
R2407 gnd.n7544 gnd.n66 585
R2408 gnd.n5687 gnd.n66 585
R2409 gnd.n3129 gnd.n64 585
R2410 gnd.n5777 gnd.n3129 585
R2411 gnd.n5660 gnd.n3122 585
R2412 gnd.n5782 gnd.n3122 585
R2413 gnd.n5662 gnd.n5659 585
R2414 gnd.n5659 gnd.n3120 585
R2415 gnd.n5663 gnd.n5658 585
R2416 gnd.n5658 gnd.n3113 585
R2417 gnd.n5664 gnd.n3112 585
R2418 gnd.n5791 gnd.n3112 585
R2419 gnd.n3207 gnd.n3106 585
R2420 gnd.n5795 gnd.n3106 585
R2421 gnd.n5669 gnd.n5668 585
R2422 gnd.n5670 gnd.n5669 585
R2423 gnd.n3206 gnd.n3097 585
R2424 gnd.n5801 gnd.n3097 585
R2425 gnd.n5654 gnd.n5653 585
R2426 gnd.n5653 gnd.n5652 585
R2427 gnd.n3209 gnd.n3086 585
R2428 gnd.n5807 gnd.n3086 585
R2429 gnd.n5592 gnd.n3211 585
R2430 gnd.n5645 gnd.n3211 585
R2431 gnd.n5593 gnd.n3077 585
R2432 gnd.n5813 gnd.n3077 585
R2433 gnd.n5594 gnd.n5590 585
R2434 gnd.n5590 gnd.n5589 585
R2435 gnd.n3219 gnd.n3066 585
R2436 gnd.n5819 gnd.n3066 585
R2437 gnd.n5599 gnd.n5598 585
R2438 gnd.n5600 gnd.n5599 585
R2439 gnd.n3218 gnd.n3057 585
R2440 gnd.n5825 gnd.n3057 585
R2441 gnd.n5579 gnd.n5578 585
R2442 gnd.n5580 gnd.n5579 585
R2443 gnd.n3224 gnd.n3046 585
R2444 gnd.n5831 gnd.n3046 585
R2445 gnd.n5574 gnd.n5573 585
R2446 gnd.n5573 gnd.n5572 585
R2447 gnd.n3226 gnd.n3034 585
R2448 gnd.n5837 gnd.n3034 585
R2449 gnd.n4995 gnd.n4994 585
R2450 gnd.n4994 gnd.n4993 585
R2451 gnd.n4996 gnd.n3022 585
R2452 gnd.n5843 gnd.n3022 585
R2453 gnd.n2233 gnd.n900 585
R2454 gnd.n900 gnd.n877 585
R2455 gnd.n2234 gnd.n961 585
R2456 gnd.n961 gnd.n951 585
R2457 gnd.n2236 gnd.n2235 585
R2458 gnd.n2237 gnd.n2236 585
R2459 gnd.n962 gnd.n960 585
R2460 gnd.n969 gnd.n960 585
R2461 gnd.n2227 gnd.n2226 585
R2462 gnd.n2226 gnd.n2225 585
R2463 gnd.n965 gnd.n964 585
R2464 gnd.n1952 gnd.n965 585
R2465 gnd.n1938 gnd.n988 585
R2466 gnd.n988 gnd.n978 585
R2467 gnd.n1940 gnd.n1939 585
R2468 gnd.n1941 gnd.n1940 585
R2469 gnd.n989 gnd.n987 585
R2470 gnd.n987 gnd.n985 585
R2471 gnd.n1933 gnd.n1932 585
R2472 gnd.n1932 gnd.n1931 585
R2473 gnd.n992 gnd.n991 585
R2474 gnd.n1001 gnd.n992 585
R2475 gnd.n1889 gnd.n1015 585
R2476 gnd.n1015 gnd.n1000 585
R2477 gnd.n1891 gnd.n1890 585
R2478 gnd.n1892 gnd.n1891 585
R2479 gnd.n1016 gnd.n1014 585
R2480 gnd.n1023 gnd.n1014 585
R2481 gnd.n1884 gnd.n1883 585
R2482 gnd.n1883 gnd.n1882 585
R2483 gnd.n1019 gnd.n1018 585
R2484 gnd.n1863 gnd.n1019 585
R2485 gnd.n1849 gnd.n1042 585
R2486 gnd.n1042 gnd.n1032 585
R2487 gnd.n1851 gnd.n1850 585
R2488 gnd.n1852 gnd.n1851 585
R2489 gnd.n1043 gnd.n1041 585
R2490 gnd.n1840 gnd.n1041 585
R2491 gnd.n1844 gnd.n1843 585
R2492 gnd.n1843 gnd.n1842 585
R2493 gnd.n1046 gnd.n1045 585
R2494 gnd.n1055 gnd.n1046 585
R2495 gnd.n1802 gnd.n1068 585
R2496 gnd.n1068 gnd.n1054 585
R2497 gnd.n1804 gnd.n1803 585
R2498 gnd.n1805 gnd.n1804 585
R2499 gnd.n1069 gnd.n1067 585
R2500 gnd.n1076 gnd.n1067 585
R2501 gnd.n1797 gnd.n1796 585
R2502 gnd.n1796 gnd.n1795 585
R2503 gnd.n1072 gnd.n1071 585
R2504 gnd.n1776 gnd.n1072 585
R2505 gnd.n1762 gnd.n1095 585
R2506 gnd.n1095 gnd.n1085 585
R2507 gnd.n1764 gnd.n1763 585
R2508 gnd.n1765 gnd.n1764 585
R2509 gnd.n1096 gnd.n1094 585
R2510 gnd.n1753 gnd.n1094 585
R2511 gnd.n1757 gnd.n1756 585
R2512 gnd.n1756 gnd.n1755 585
R2513 gnd.n1099 gnd.n1098 585
R2514 gnd.n1708 gnd.n1099 585
R2515 gnd.n1201 gnd.n1200 585
R2516 gnd.n1202 gnd.n1201 585
R2517 gnd.n1181 gnd.n1180 585
R2518 gnd.n1184 gnd.n1181 585
R2519 gnd.n1718 gnd.n1717 585
R2520 gnd.n1717 gnd.n1716 585
R2521 gnd.n1719 gnd.n1175 585
R2522 gnd.n1211 gnd.n1175 585
R2523 gnd.n1721 gnd.n1720 585
R2524 gnd.n1722 gnd.n1721 585
R2525 gnd.n1176 gnd.n1174 585
R2526 gnd.n1686 gnd.n1174 585
R2527 gnd.n1670 gnd.n1669 585
R2528 gnd.n1669 gnd.n1162 585
R2529 gnd.n1671 gnd.n1226 585
R2530 gnd.n1226 gnd.n1161 585
R2531 gnd.n1673 gnd.n1672 585
R2532 gnd.n1674 gnd.n1673 585
R2533 gnd.n1227 gnd.n1225 585
R2534 gnd.n1225 gnd.n1222 585
R2535 gnd.n1662 gnd.n1661 585
R2536 gnd.n1661 gnd.n1660 585
R2537 gnd.n1230 gnd.n1229 585
R2538 gnd.n1237 gnd.n1230 585
R2539 gnd.n1636 gnd.n1635 585
R2540 gnd.n1637 gnd.n1636 585
R2541 gnd.n1249 gnd.n1248 585
R2542 gnd.n1256 gnd.n1248 585
R2543 gnd.n1631 gnd.n1630 585
R2544 gnd.n1630 gnd.n1629 585
R2545 gnd.n1252 gnd.n1251 585
R2546 gnd.n1619 gnd.n1252 585
R2547 gnd.n1606 gnd.n1276 585
R2548 gnd.n1276 gnd.n1275 585
R2549 gnd.n1608 gnd.n1607 585
R2550 gnd.n1609 gnd.n1608 585
R2551 gnd.n1277 gnd.n1274 585
R2552 gnd.n1284 gnd.n1274 585
R2553 gnd.n1601 gnd.n1600 585
R2554 gnd.n1600 gnd.n1599 585
R2555 gnd.n1280 gnd.n1279 585
R2556 gnd.n1588 gnd.n1280 585
R2557 gnd.n1575 gnd.n1301 585
R2558 gnd.n1301 gnd.n1300 585
R2559 gnd.n1577 gnd.n1576 585
R2560 gnd.n1578 gnd.n1577 585
R2561 gnd.n1571 gnd.n1299 585
R2562 gnd.n1570 gnd.n1569 585
R2563 gnd.n1304 gnd.n1303 585
R2564 gnd.n1567 gnd.n1304 585
R2565 gnd.n1326 gnd.n1325 585
R2566 gnd.n1329 gnd.n1328 585
R2567 gnd.n1327 gnd.n1322 585
R2568 gnd.n1334 gnd.n1333 585
R2569 gnd.n1336 gnd.n1335 585
R2570 gnd.n1339 gnd.n1338 585
R2571 gnd.n1337 gnd.n1320 585
R2572 gnd.n1344 gnd.n1343 585
R2573 gnd.n1346 gnd.n1345 585
R2574 gnd.n1349 gnd.n1348 585
R2575 gnd.n1347 gnd.n1318 585
R2576 gnd.n1354 gnd.n1353 585
R2577 gnd.n1358 gnd.n1355 585
R2578 gnd.n1359 gnd.n1296 585
R2579 gnd.n2239 gnd.n915 585
R2580 gnd.n2306 gnd.n2305 585
R2581 gnd.n2308 gnd.n2307 585
R2582 gnd.n2310 gnd.n2309 585
R2583 gnd.n2312 gnd.n2311 585
R2584 gnd.n2314 gnd.n2313 585
R2585 gnd.n2316 gnd.n2315 585
R2586 gnd.n2318 gnd.n2317 585
R2587 gnd.n2320 gnd.n2319 585
R2588 gnd.n2322 gnd.n2321 585
R2589 gnd.n2324 gnd.n2323 585
R2590 gnd.n2326 gnd.n2325 585
R2591 gnd.n2328 gnd.n2327 585
R2592 gnd.n2331 gnd.n2330 585
R2593 gnd.n2329 gnd.n903 585
R2594 gnd.n2335 gnd.n901 585
R2595 gnd.n2337 gnd.n2336 585
R2596 gnd.n2338 gnd.n2337 585
R2597 gnd.n2240 gnd.n956 585
R2598 gnd.n2240 gnd.n877 585
R2599 gnd.n2242 gnd.n2241 585
R2600 gnd.n2241 gnd.n951 585
R2601 gnd.n2238 gnd.n955 585
R2602 gnd.n2238 gnd.n2237 585
R2603 gnd.n2217 gnd.n957 585
R2604 gnd.n969 gnd.n957 585
R2605 gnd.n2216 gnd.n967 585
R2606 gnd.n2225 gnd.n967 585
R2607 gnd.n1951 gnd.n974 585
R2608 gnd.n1952 gnd.n1951 585
R2609 gnd.n1950 gnd.n1949 585
R2610 gnd.n1950 gnd.n978 585
R2611 gnd.n1948 gnd.n980 585
R2612 gnd.n1941 gnd.n980 585
R2613 gnd.n993 gnd.n981 585
R2614 gnd.n993 gnd.n985 585
R2615 gnd.n1897 gnd.n994 585
R2616 gnd.n1931 gnd.n994 585
R2617 gnd.n1896 gnd.n1895 585
R2618 gnd.n1895 gnd.n1001 585
R2619 gnd.n1894 gnd.n1009 585
R2620 gnd.n1894 gnd.n1000 585
R2621 gnd.n1893 gnd.n1011 585
R2622 gnd.n1893 gnd.n1892 585
R2623 gnd.n1872 gnd.n1010 585
R2624 gnd.n1023 gnd.n1010 585
R2625 gnd.n1871 gnd.n1021 585
R2626 gnd.n1882 gnd.n1021 585
R2627 gnd.n1862 gnd.n1028 585
R2628 gnd.n1863 gnd.n1862 585
R2629 gnd.n1861 gnd.n1860 585
R2630 gnd.n1861 gnd.n1032 585
R2631 gnd.n1859 gnd.n1034 585
R2632 gnd.n1852 gnd.n1034 585
R2633 gnd.n1839 gnd.n1035 585
R2634 gnd.n1840 gnd.n1839 585
R2635 gnd.n1810 gnd.n1048 585
R2636 gnd.n1842 gnd.n1048 585
R2637 gnd.n1809 gnd.n1808 585
R2638 gnd.n1808 gnd.n1055 585
R2639 gnd.n1807 gnd.n1062 585
R2640 gnd.n1807 gnd.n1054 585
R2641 gnd.n1806 gnd.n1064 585
R2642 gnd.n1806 gnd.n1805 585
R2643 gnd.n1785 gnd.n1063 585
R2644 gnd.n1076 gnd.n1063 585
R2645 gnd.n1784 gnd.n1074 585
R2646 gnd.n1795 gnd.n1074 585
R2647 gnd.n1775 gnd.n1081 585
R2648 gnd.n1776 gnd.n1775 585
R2649 gnd.n1774 gnd.n1773 585
R2650 gnd.n1774 gnd.n1085 585
R2651 gnd.n1772 gnd.n1087 585
R2652 gnd.n1765 gnd.n1087 585
R2653 gnd.n1752 gnd.n1088 585
R2654 gnd.n1753 gnd.n1752 585
R2655 gnd.n1705 gnd.n1101 585
R2656 gnd.n1755 gnd.n1101 585
R2657 gnd.n1707 gnd.n1706 585
R2658 gnd.n1708 gnd.n1707 585
R2659 gnd.n1700 gnd.n1203 585
R2660 gnd.n1203 gnd.n1202 585
R2661 gnd.n1698 gnd.n1697 585
R2662 gnd.n1697 gnd.n1184 585
R2663 gnd.n1695 gnd.n1182 585
R2664 gnd.n1716 gnd.n1182 585
R2665 gnd.n1213 gnd.n1212 585
R2666 gnd.n1212 gnd.n1211 585
R2667 gnd.n1689 gnd.n1172 585
R2668 gnd.n1722 gnd.n1172 585
R2669 gnd.n1688 gnd.n1687 585
R2670 gnd.n1687 gnd.n1686 585
R2671 gnd.n1684 gnd.n1215 585
R2672 gnd.n1684 gnd.n1162 585
R2673 gnd.n1683 gnd.n1682 585
R2674 gnd.n1683 gnd.n1161 585
R2675 gnd.n1218 gnd.n1217 585
R2676 gnd.n1674 gnd.n1217 585
R2677 gnd.n1642 gnd.n1641 585
R2678 gnd.n1641 gnd.n1222 585
R2679 gnd.n1643 gnd.n1231 585
R2680 gnd.n1660 gnd.n1231 585
R2681 gnd.n1640 gnd.n1639 585
R2682 gnd.n1639 gnd.n1237 585
R2683 gnd.n1638 gnd.n1245 585
R2684 gnd.n1638 gnd.n1637 585
R2685 gnd.n1623 gnd.n1246 585
R2686 gnd.n1256 gnd.n1246 585
R2687 gnd.n1622 gnd.n1254 585
R2688 gnd.n1629 gnd.n1254 585
R2689 gnd.n1621 gnd.n1620 585
R2690 gnd.n1620 gnd.n1619 585
R2691 gnd.n1265 gnd.n1262 585
R2692 gnd.n1275 gnd.n1265 585
R2693 gnd.n1611 gnd.n1610 585
R2694 gnd.n1610 gnd.n1609 585
R2695 gnd.n1271 gnd.n1270 585
R2696 gnd.n1284 gnd.n1271 585
R2697 gnd.n1591 gnd.n1282 585
R2698 gnd.n1599 gnd.n1282 585
R2699 gnd.n1590 gnd.n1589 585
R2700 gnd.n1589 gnd.n1588 585
R2701 gnd.n1291 gnd.n1289 585
R2702 gnd.n1300 gnd.n1291 585
R2703 gnd.n1580 gnd.n1579 585
R2704 gnd.n1579 gnd.n1578 585
R2705 gnd.n5316 gnd.n5315 585
R2706 gnd.n5317 gnd.n5316 585
R2707 gnd.n5230 gnd.n3306 585
R2708 gnd.n5225 gnd.n3306 585
R2709 gnd.n5229 gnd.n5228 585
R2710 gnd.n5228 gnd.n5227 585
R2711 gnd.n3309 gnd.n3308 585
R2712 gnd.n4953 gnd.n3309 585
R2713 gnd.n4942 gnd.n3380 585
R2714 gnd.n3380 gnd.n3379 585
R2715 gnd.n4944 gnd.n4943 585
R2716 gnd.n4945 gnd.n4944 585
R2717 gnd.n4941 gnd.n3377 585
R2718 gnd.n3385 gnd.n3377 585
R2719 gnd.n4940 gnd.n4939 585
R2720 gnd.n4939 gnd.n4938 585
R2721 gnd.n3382 gnd.n3381 585
R2722 gnd.n4820 gnd.n3382 585
R2723 gnd.n4919 gnd.n4918 585
R2724 gnd.n4920 gnd.n4919 585
R2725 gnd.n4917 gnd.n3397 585
R2726 gnd.n3397 gnd.n3393 585
R2727 gnd.n4916 gnd.n4915 585
R2728 gnd.n4915 gnd.n4914 585
R2729 gnd.n3399 gnd.n3398 585
R2730 gnd.n4829 gnd.n3399 585
R2731 gnd.n4896 gnd.n4895 585
R2732 gnd.n4897 gnd.n4896 585
R2733 gnd.n4894 gnd.n3410 585
R2734 gnd.n3410 gnd.n3407 585
R2735 gnd.n4893 gnd.n4892 585
R2736 gnd.n4892 gnd.n4891 585
R2737 gnd.n3412 gnd.n3411 585
R2738 gnd.n4836 gnd.n3412 585
R2739 gnd.n4876 gnd.n4875 585
R2740 gnd.n4877 gnd.n4876 585
R2741 gnd.n4874 gnd.n3423 585
R2742 gnd.n4869 gnd.n3423 585
R2743 gnd.n4873 gnd.n4872 585
R2744 gnd.n4872 gnd.n4871 585
R2745 gnd.n3425 gnd.n3424 585
R2746 gnd.n3437 gnd.n3425 585
R2747 gnd.n4806 gnd.n4805 585
R2748 gnd.n4806 gnd.n3436 585
R2749 gnd.n4810 gnd.n4809 585
R2750 gnd.n4809 gnd.n4808 585
R2751 gnd.n4811 gnd.n3443 585
R2752 gnd.n4849 gnd.n3443 585
R2753 gnd.n4812 gnd.n3452 585
R2754 gnd.n4737 gnd.n3452 585
R2755 gnd.n4814 gnd.n4813 585
R2756 gnd.n4815 gnd.n4814 585
R2757 gnd.n4804 gnd.n3451 585
R2758 gnd.n4798 gnd.n3451 585
R2759 gnd.n4803 gnd.n4802 585
R2760 gnd.n4802 gnd.n4801 585
R2761 gnd.n3454 gnd.n3453 585
R2762 gnd.n4787 gnd.n3454 585
R2763 gnd.n4777 gnd.n3471 585
R2764 gnd.n3471 gnd.n3463 585
R2765 gnd.n4779 gnd.n4778 585
R2766 gnd.n4780 gnd.n4779 585
R2767 gnd.n4776 gnd.n3470 585
R2768 gnd.n3475 gnd.n3470 585
R2769 gnd.n4775 gnd.n4774 585
R2770 gnd.n4774 gnd.n4773 585
R2771 gnd.n3473 gnd.n3472 585
R2772 gnd.n4728 gnd.n3473 585
R2773 gnd.n4761 gnd.n4760 585
R2774 gnd.n4762 gnd.n4761 585
R2775 gnd.n4759 gnd.n3486 585
R2776 gnd.n3486 gnd.n3482 585
R2777 gnd.n4758 gnd.n4757 585
R2778 gnd.n4757 gnd.n4756 585
R2779 gnd.n3488 gnd.n3487 585
R2780 gnd.n4718 gnd.n3488 585
R2781 gnd.n4703 gnd.n4702 585
R2782 gnd.n4702 gnd.n3498 585
R2783 gnd.n4704 gnd.n3508 585
R2784 gnd.n4687 gnd.n3508 585
R2785 gnd.n4706 gnd.n4705 585
R2786 gnd.n4707 gnd.n4706 585
R2787 gnd.n4701 gnd.n3507 585
R2788 gnd.n3507 gnd.n3504 585
R2789 gnd.n4700 gnd.n4699 585
R2790 gnd.n4699 gnd.n4698 585
R2791 gnd.n3510 gnd.n3509 585
R2792 gnd.n4678 gnd.n3510 585
R2793 gnd.n4663 gnd.n4662 585
R2794 gnd.n4662 gnd.n3521 585
R2795 gnd.n4664 gnd.n3531 585
R2796 gnd.n4651 gnd.n3531 585
R2797 gnd.n4666 gnd.n4665 585
R2798 gnd.n4667 gnd.n4666 585
R2799 gnd.n4661 gnd.n3530 585
R2800 gnd.n3530 gnd.n3527 585
R2801 gnd.n4660 gnd.n4659 585
R2802 gnd.n4659 gnd.n4658 585
R2803 gnd.n3533 gnd.n3532 585
R2804 gnd.n3546 gnd.n3533 585
R2805 gnd.n4635 gnd.n4634 585
R2806 gnd.n4636 gnd.n4635 585
R2807 gnd.n4633 gnd.n3548 585
R2808 gnd.n4628 gnd.n3548 585
R2809 gnd.n4632 gnd.n4631 585
R2810 gnd.n4631 gnd.n4630 585
R2811 gnd.n3550 gnd.n3549 585
R2812 gnd.n4615 gnd.n3550 585
R2813 gnd.n4603 gnd.n3568 585
R2814 gnd.n3568 gnd.n3560 585
R2815 gnd.n4605 gnd.n4604 585
R2816 gnd.n4606 gnd.n4605 585
R2817 gnd.n4602 gnd.n3567 585
R2818 gnd.n4546 gnd.n3567 585
R2819 gnd.n4601 gnd.n4600 585
R2820 gnd.n4600 gnd.n4599 585
R2821 gnd.n3570 gnd.n3569 585
R2822 gnd.n4574 gnd.n3570 585
R2823 gnd.n4587 gnd.n4586 585
R2824 gnd.n4588 gnd.n4587 585
R2825 gnd.n4585 gnd.n3581 585
R2826 gnd.n4580 gnd.n3581 585
R2827 gnd.n4584 gnd.n4583 585
R2828 gnd.n4583 gnd.n4582 585
R2829 gnd.n3583 gnd.n3582 585
R2830 gnd.n4569 gnd.n3583 585
R2831 gnd.n4520 gnd.n4517 585
R2832 gnd.n4520 gnd.n4519 585
R2833 gnd.n4521 gnd.n4516 585
R2834 gnd.n4521 gnd.n3597 585
R2835 gnd.n4523 gnd.n4522 585
R2836 gnd.n4522 gnd.n3596 585
R2837 gnd.n4524 gnd.n4514 585
R2838 gnd.n4514 gnd.n4513 585
R2839 gnd.n4526 gnd.n4525 585
R2840 gnd.n4527 gnd.n4526 585
R2841 gnd.n4515 gnd.n3607 585
R2842 gnd.n4503 gnd.n3607 585
R2843 gnd.n2910 gnd.n2909 585
R2844 gnd.n2914 gnd.n2910 585
R2845 gnd.n5962 gnd.n5961 585
R2846 gnd.n5961 gnd.n5960 585
R2847 gnd.n5963 gnd.n2888 585
R2848 gnd.n4496 gnd.n2888 585
R2849 gnd.n6028 gnd.n6027 585
R2850 gnd.n6026 gnd.n2887 585
R2851 gnd.n6025 gnd.n2886 585
R2852 gnd.n6030 gnd.n2886 585
R2853 gnd.n6024 gnd.n6023 585
R2854 gnd.n6022 gnd.n6021 585
R2855 gnd.n6020 gnd.n6019 585
R2856 gnd.n6018 gnd.n6017 585
R2857 gnd.n6016 gnd.n6015 585
R2858 gnd.n6014 gnd.n6013 585
R2859 gnd.n6012 gnd.n6011 585
R2860 gnd.n6010 gnd.n6009 585
R2861 gnd.n6008 gnd.n6007 585
R2862 gnd.n6006 gnd.n6005 585
R2863 gnd.n6004 gnd.n6003 585
R2864 gnd.n6002 gnd.n6001 585
R2865 gnd.n6000 gnd.n5999 585
R2866 gnd.n5998 gnd.n5997 585
R2867 gnd.n5996 gnd.n5995 585
R2868 gnd.n5994 gnd.n5993 585
R2869 gnd.n5992 gnd.n5991 585
R2870 gnd.n5990 gnd.n5989 585
R2871 gnd.n5988 gnd.n5987 585
R2872 gnd.n5986 gnd.n5985 585
R2873 gnd.n5984 gnd.n5983 585
R2874 gnd.n5982 gnd.n5981 585
R2875 gnd.n5980 gnd.n5979 585
R2876 gnd.n5978 gnd.n5977 585
R2877 gnd.n5976 gnd.n5975 585
R2878 gnd.n5974 gnd.n5973 585
R2879 gnd.n5972 gnd.n5971 585
R2880 gnd.n5970 gnd.n5969 585
R2881 gnd.n5968 gnd.n2851 585
R2882 gnd.n6033 gnd.n6032 585
R2883 gnd.n2853 gnd.n2850 585
R2884 gnd.n3612 gnd.n3611 585
R2885 gnd.n3614 gnd.n3613 585
R2886 gnd.n3617 gnd.n3616 585
R2887 gnd.n3619 gnd.n3618 585
R2888 gnd.n3621 gnd.n3620 585
R2889 gnd.n3623 gnd.n3622 585
R2890 gnd.n3625 gnd.n3624 585
R2891 gnd.n3627 gnd.n3626 585
R2892 gnd.n3629 gnd.n3628 585
R2893 gnd.n3631 gnd.n3630 585
R2894 gnd.n3633 gnd.n3632 585
R2895 gnd.n3635 gnd.n3634 585
R2896 gnd.n3637 gnd.n3636 585
R2897 gnd.n3639 gnd.n3638 585
R2898 gnd.n3641 gnd.n3640 585
R2899 gnd.n3643 gnd.n3642 585
R2900 gnd.n3645 gnd.n3644 585
R2901 gnd.n3647 gnd.n3646 585
R2902 gnd.n3649 gnd.n3648 585
R2903 gnd.n3651 gnd.n3650 585
R2904 gnd.n3653 gnd.n3652 585
R2905 gnd.n3655 gnd.n3654 585
R2906 gnd.n3657 gnd.n3656 585
R2907 gnd.n3659 gnd.n3658 585
R2908 gnd.n3661 gnd.n3660 585
R2909 gnd.n3663 gnd.n3662 585
R2910 gnd.n3665 gnd.n3664 585
R2911 gnd.n3667 gnd.n3666 585
R2912 gnd.n3669 gnd.n3668 585
R2913 gnd.n3671 gnd.n3670 585
R2914 gnd.n3673 gnd.n3672 585
R2915 gnd.n5320 gnd.n5319 585
R2916 gnd.n5322 gnd.n5321 585
R2917 gnd.n5324 gnd.n5323 585
R2918 gnd.n5326 gnd.n5325 585
R2919 gnd.n5328 gnd.n5327 585
R2920 gnd.n5330 gnd.n5329 585
R2921 gnd.n5332 gnd.n5331 585
R2922 gnd.n5334 gnd.n5333 585
R2923 gnd.n5336 gnd.n5335 585
R2924 gnd.n5338 gnd.n5337 585
R2925 gnd.n5340 gnd.n5339 585
R2926 gnd.n5342 gnd.n5341 585
R2927 gnd.n5344 gnd.n5343 585
R2928 gnd.n5346 gnd.n5345 585
R2929 gnd.n5348 gnd.n5347 585
R2930 gnd.n5350 gnd.n5349 585
R2931 gnd.n5352 gnd.n5351 585
R2932 gnd.n5354 gnd.n5353 585
R2933 gnd.n5356 gnd.n5355 585
R2934 gnd.n5358 gnd.n5357 585
R2935 gnd.n5360 gnd.n5359 585
R2936 gnd.n5362 gnd.n5361 585
R2937 gnd.n5364 gnd.n5363 585
R2938 gnd.n5366 gnd.n5365 585
R2939 gnd.n5368 gnd.n5367 585
R2940 gnd.n5370 gnd.n5369 585
R2941 gnd.n5372 gnd.n5371 585
R2942 gnd.n5374 gnd.n5373 585
R2943 gnd.n5376 gnd.n5375 585
R2944 gnd.n5378 gnd.n3299 585
R2945 gnd.n5380 gnd.n5379 585
R2946 gnd.n5382 gnd.n3263 585
R2947 gnd.n5384 gnd.n5383 585
R2948 gnd.n5387 gnd.n5386 585
R2949 gnd.n3266 gnd.n3264 585
R2950 gnd.n5253 gnd.n5252 585
R2951 gnd.n5255 gnd.n5254 585
R2952 gnd.n5258 gnd.n5257 585
R2953 gnd.n5260 gnd.n5259 585
R2954 gnd.n5262 gnd.n5261 585
R2955 gnd.n5264 gnd.n5263 585
R2956 gnd.n5266 gnd.n5265 585
R2957 gnd.n5268 gnd.n5267 585
R2958 gnd.n5270 gnd.n5269 585
R2959 gnd.n5272 gnd.n5271 585
R2960 gnd.n5274 gnd.n5273 585
R2961 gnd.n5276 gnd.n5275 585
R2962 gnd.n5278 gnd.n5277 585
R2963 gnd.n5280 gnd.n5279 585
R2964 gnd.n5282 gnd.n5281 585
R2965 gnd.n5284 gnd.n5283 585
R2966 gnd.n5286 gnd.n5285 585
R2967 gnd.n5288 gnd.n5287 585
R2968 gnd.n5290 gnd.n5289 585
R2969 gnd.n5292 gnd.n5291 585
R2970 gnd.n5294 gnd.n5293 585
R2971 gnd.n5296 gnd.n5295 585
R2972 gnd.n5298 gnd.n5297 585
R2973 gnd.n5300 gnd.n5299 585
R2974 gnd.n5302 gnd.n5301 585
R2975 gnd.n5304 gnd.n5303 585
R2976 gnd.n5306 gnd.n5305 585
R2977 gnd.n5308 gnd.n5307 585
R2978 gnd.n5310 gnd.n5309 585
R2979 gnd.n5312 gnd.n5311 585
R2980 gnd.n5313 gnd.n3307 585
R2981 gnd.n5318 gnd.n3302 585
R2982 gnd.n5318 gnd.n5317 585
R2983 gnd.n4949 gnd.n3303 585
R2984 gnd.n5225 gnd.n3303 585
R2985 gnd.n4950 gnd.n3311 585
R2986 gnd.n5227 gnd.n3311 585
R2987 gnd.n4952 gnd.n4951 585
R2988 gnd.n4953 gnd.n4952 585
R2989 gnd.n4948 gnd.n3373 585
R2990 gnd.n3379 gnd.n3373 585
R2991 gnd.n4947 gnd.n4946 585
R2992 gnd.n4946 gnd.n4945 585
R2993 gnd.n3375 gnd.n3374 585
R2994 gnd.n3385 gnd.n3375 585
R2995 gnd.n4819 gnd.n3384 585
R2996 gnd.n4938 gnd.n3384 585
R2997 gnd.n4822 gnd.n4821 585
R2998 gnd.n4821 gnd.n4820 585
R2999 gnd.n4823 gnd.n3395 585
R3000 gnd.n4920 gnd.n3395 585
R3001 gnd.n4825 gnd.n4824 585
R3002 gnd.n4824 gnd.n3393 585
R3003 gnd.n4826 gnd.n3400 585
R3004 gnd.n4914 gnd.n3400 585
R3005 gnd.n4831 gnd.n4830 585
R3006 gnd.n4830 gnd.n4829 585
R3007 gnd.n4832 gnd.n3408 585
R3008 gnd.n4897 gnd.n3408 585
R3009 gnd.n4834 gnd.n4833 585
R3010 gnd.n4833 gnd.n3407 585
R3011 gnd.n4835 gnd.n3414 585
R3012 gnd.n4891 gnd.n3414 585
R3013 gnd.n4838 gnd.n4837 585
R3014 gnd.n4837 gnd.n4836 585
R3015 gnd.n4839 gnd.n3421 585
R3016 gnd.n4877 gnd.n3421 585
R3017 gnd.n4840 gnd.n3428 585
R3018 gnd.n4869 gnd.n3428 585
R3019 gnd.n4841 gnd.n3427 585
R3020 gnd.n4871 gnd.n3427 585
R3021 gnd.n4843 gnd.n4842 585
R3022 gnd.n4843 gnd.n3437 585
R3023 gnd.n4845 gnd.n4844 585
R3024 gnd.n4844 gnd.n3436 585
R3025 gnd.n4846 gnd.n3446 585
R3026 gnd.n4808 gnd.n3446 585
R3027 gnd.n4848 gnd.n4847 585
R3028 gnd.n4849 gnd.n4848 585
R3029 gnd.n4818 gnd.n3445 585
R3030 gnd.n4737 gnd.n3445 585
R3031 gnd.n4817 gnd.n4816 585
R3032 gnd.n4816 gnd.n4815 585
R3033 gnd.n3448 gnd.n3447 585
R3034 gnd.n4798 gnd.n3448 585
R3035 gnd.n4784 gnd.n3456 585
R3036 gnd.n4801 gnd.n3456 585
R3037 gnd.n4786 gnd.n4785 585
R3038 gnd.n4787 gnd.n4786 585
R3039 gnd.n4783 gnd.n3465 585
R3040 gnd.n3465 gnd.n3463 585
R3041 gnd.n4782 gnd.n4781 585
R3042 gnd.n4781 gnd.n4780 585
R3043 gnd.n3467 gnd.n3466 585
R3044 gnd.n3475 gnd.n3467 585
R3045 gnd.n4725 gnd.n3474 585
R3046 gnd.n4773 gnd.n3474 585
R3047 gnd.n4727 gnd.n4726 585
R3048 gnd.n4728 gnd.n4727 585
R3049 gnd.n4724 gnd.n3484 585
R3050 gnd.n4762 gnd.n3484 585
R3051 gnd.n4723 gnd.n4722 585
R3052 gnd.n4722 gnd.n3482 585
R3053 gnd.n4721 gnd.n3490 585
R3054 gnd.n4756 gnd.n3490 585
R3055 gnd.n4720 gnd.n4719 585
R3056 gnd.n4719 gnd.n4718 585
R3057 gnd.n3497 gnd.n3496 585
R3058 gnd.n3498 gnd.n3497 585
R3059 gnd.n4686 gnd.n4685 585
R3060 gnd.n4687 gnd.n4686 585
R3061 gnd.n4684 gnd.n3505 585
R3062 gnd.n4707 gnd.n3505 585
R3063 gnd.n4683 gnd.n4682 585
R3064 gnd.n4682 gnd.n3504 585
R3065 gnd.n4681 gnd.n3512 585
R3066 gnd.n4698 gnd.n3512 585
R3067 gnd.n4680 gnd.n4679 585
R3068 gnd.n4679 gnd.n4678 585
R3069 gnd.n3520 gnd.n3519 585
R3070 gnd.n3521 gnd.n3520 585
R3071 gnd.n4653 gnd.n4652 585
R3072 gnd.n4652 gnd.n4651 585
R3073 gnd.n4654 gnd.n3528 585
R3074 gnd.n4667 gnd.n3528 585
R3075 gnd.n4655 gnd.n3536 585
R3076 gnd.n3536 gnd.n3527 585
R3077 gnd.n4657 gnd.n4656 585
R3078 gnd.n4658 gnd.n4657 585
R3079 gnd.n3537 gnd.n3535 585
R3080 gnd.n3546 gnd.n3535 585
R3081 gnd.n4610 gnd.n3545 585
R3082 gnd.n4636 gnd.n3545 585
R3083 gnd.n4611 gnd.n3553 585
R3084 gnd.n4628 gnd.n3553 585
R3085 gnd.n4612 gnd.n3552 585
R3086 gnd.n4630 gnd.n3552 585
R3087 gnd.n4614 gnd.n4613 585
R3088 gnd.n4615 gnd.n4614 585
R3089 gnd.n4609 gnd.n3562 585
R3090 gnd.n3562 gnd.n3560 585
R3091 gnd.n4608 gnd.n4607 585
R3092 gnd.n4607 gnd.n4606 585
R3093 gnd.n3564 gnd.n3563 585
R3094 gnd.n4546 gnd.n3564 585
R3095 gnd.n4573 gnd.n3572 585
R3096 gnd.n4599 gnd.n3572 585
R3097 gnd.n4576 gnd.n4575 585
R3098 gnd.n4575 gnd.n4574 585
R3099 gnd.n4577 gnd.n3579 585
R3100 gnd.n4588 gnd.n3579 585
R3101 gnd.n4579 gnd.n4578 585
R3102 gnd.n4580 gnd.n4579 585
R3103 gnd.n4572 gnd.n3585 585
R3104 gnd.n4582 gnd.n3585 585
R3105 gnd.n4571 gnd.n4570 585
R3106 gnd.n4570 gnd.n4569 585
R3107 gnd.n3588 gnd.n3587 585
R3108 gnd.n4519 gnd.n3588 585
R3109 gnd.n4508 gnd.n4507 585
R3110 gnd.n4507 gnd.n3597 585
R3111 gnd.n4509 gnd.n3608 585
R3112 gnd.n3608 gnd.n3596 585
R3113 gnd.n4511 gnd.n4510 585
R3114 gnd.n4513 gnd.n4511 585
R3115 gnd.n4506 gnd.n3605 585
R3116 gnd.n4527 gnd.n3605 585
R3117 gnd.n4505 gnd.n4504 585
R3118 gnd.n4504 gnd.n4503 585
R3119 gnd.n4501 gnd.n4500 585
R3120 gnd.n4501 gnd.n2914 585
R3121 gnd.n4499 gnd.n2912 585
R3122 gnd.n5960 gnd.n2912 585
R3123 gnd.n4498 gnd.n4497 585
R3124 gnd.n4497 gnd.n4496 585
R3125 gnd.n6169 gnd.n6168 585
R3126 gnd.n6168 gnd.n6167 585
R3127 gnd.n6170 gnd.n2565 585
R3128 gnd.n6160 gnd.n2565 585
R3129 gnd.n6172 gnd.n6171 585
R3130 gnd.n6173 gnd.n6172 585
R3131 gnd.n2550 gnd.n2549 585
R3132 gnd.n4314 gnd.n2550 585
R3133 gnd.n6181 gnd.n6180 585
R3134 gnd.n6180 gnd.n6179 585
R3135 gnd.n6182 gnd.n2544 585
R3136 gnd.n4308 gnd.n2544 585
R3137 gnd.n6184 gnd.n6183 585
R3138 gnd.n6185 gnd.n6184 585
R3139 gnd.n2530 gnd.n2529 585
R3140 gnd.n4303 gnd.n2530 585
R3141 gnd.n6193 gnd.n6192 585
R3142 gnd.n6192 gnd.n6191 585
R3143 gnd.n6194 gnd.n2524 585
R3144 gnd.n4298 gnd.n2524 585
R3145 gnd.n6196 gnd.n6195 585
R3146 gnd.n6197 gnd.n6196 585
R3147 gnd.n2510 gnd.n2509 585
R3148 gnd.n4331 gnd.n2510 585
R3149 gnd.n6205 gnd.n6204 585
R3150 gnd.n6204 gnd.n6203 585
R3151 gnd.n6206 gnd.n2504 585
R3152 gnd.n4291 gnd.n2504 585
R3153 gnd.n6208 gnd.n6207 585
R3154 gnd.n6209 gnd.n6208 585
R3155 gnd.n2490 gnd.n2489 585
R3156 gnd.n4283 gnd.n2490 585
R3157 gnd.n6217 gnd.n6216 585
R3158 gnd.n6216 gnd.n6215 585
R3159 gnd.n6218 gnd.n2487 585
R3160 gnd.n4251 gnd.n2487 585
R3161 gnd.n6221 gnd.n6220 585
R3162 gnd.n6222 gnd.n6221 585
R3163 gnd.n2488 gnd.n2473 585
R3164 gnd.n4242 gnd.n2473 585
R3165 gnd.n6230 gnd.n6229 585
R3166 gnd.n6229 gnd.n6228 585
R3167 gnd.n6231 gnd.n2470 585
R3168 gnd.n4227 gnd.n2470 585
R3169 gnd.n6234 gnd.n6233 585
R3170 gnd.n6235 gnd.n6234 585
R3171 gnd.n2471 gnd.n2456 585
R3172 gnd.n4264 gnd.n2456 585
R3173 gnd.n6243 gnd.n6242 585
R3174 gnd.n6242 gnd.n6241 585
R3175 gnd.n6244 gnd.n2452 585
R3176 gnd.n4220 gnd.n2452 585
R3177 gnd.n6247 gnd.n6246 585
R3178 gnd.n6248 gnd.n6247 585
R3179 gnd.n2437 gnd.n2436 585
R3180 gnd.n4211 gnd.n2437 585
R3181 gnd.n6256 gnd.n6255 585
R3182 gnd.n6255 gnd.n6254 585
R3183 gnd.n6257 gnd.n2431 585
R3184 gnd.n4205 gnd.n2431 585
R3185 gnd.n6259 gnd.n6258 585
R3186 gnd.n6260 gnd.n6259 585
R3187 gnd.n2417 gnd.n2416 585
R3188 gnd.n4197 gnd.n2417 585
R3189 gnd.n6268 gnd.n6267 585
R3190 gnd.n6267 gnd.n6266 585
R3191 gnd.n6269 gnd.n2411 585
R3192 gnd.n4142 gnd.n2411 585
R3193 gnd.n6271 gnd.n6270 585
R3194 gnd.n6272 gnd.n6271 585
R3195 gnd.n2396 gnd.n2395 585
R3196 gnd.n4148 gnd.n2396 585
R3197 gnd.n6280 gnd.n6279 585
R3198 gnd.n6279 gnd.n6278 585
R3199 gnd.n6281 gnd.n2390 585
R3200 gnd.n4154 gnd.n2390 585
R3201 gnd.n6283 gnd.n6282 585
R3202 gnd.n6284 gnd.n6283 585
R3203 gnd.n2374 gnd.n2373 585
R3204 gnd.n4160 gnd.n2374 585
R3205 gnd.n6292 gnd.n6291 585
R3206 gnd.n6291 gnd.n6290 585
R3207 gnd.n6293 gnd.n2369 585
R3208 gnd.n4166 gnd.n2369 585
R3209 gnd.n6295 gnd.n6294 585
R3210 gnd.n6296 gnd.n6295 585
R3211 gnd.n3973 gnd.n2368 585
R3212 gnd.n3976 gnd.n3975 585
R3213 gnd.n3971 gnd.n3970 585
R3214 gnd.n3970 gnd.n2363 585
R3215 gnd.n3981 gnd.n3980 585
R3216 gnd.n3983 gnd.n3969 585
R3217 gnd.n3986 gnd.n3985 585
R3218 gnd.n3967 gnd.n3966 585
R3219 gnd.n3991 gnd.n3990 585
R3220 gnd.n3993 gnd.n3965 585
R3221 gnd.n3996 gnd.n3995 585
R3222 gnd.n3963 gnd.n3962 585
R3223 gnd.n4001 gnd.n4000 585
R3224 gnd.n4003 gnd.n3961 585
R3225 gnd.n4006 gnd.n4005 585
R3226 gnd.n3959 gnd.n3958 585
R3227 gnd.n4011 gnd.n4010 585
R3228 gnd.n4013 gnd.n3954 585
R3229 gnd.n4016 gnd.n4015 585
R3230 gnd.n3952 gnd.n3951 585
R3231 gnd.n4021 gnd.n4020 585
R3232 gnd.n4023 gnd.n3950 585
R3233 gnd.n4026 gnd.n4025 585
R3234 gnd.n3948 gnd.n3947 585
R3235 gnd.n4031 gnd.n4030 585
R3236 gnd.n4033 gnd.n3946 585
R3237 gnd.n4036 gnd.n4035 585
R3238 gnd.n3944 gnd.n3943 585
R3239 gnd.n4041 gnd.n4040 585
R3240 gnd.n4043 gnd.n3942 585
R3241 gnd.n4046 gnd.n4045 585
R3242 gnd.n3940 gnd.n3939 585
R3243 gnd.n4051 gnd.n4050 585
R3244 gnd.n4053 gnd.n3938 585
R3245 gnd.n4056 gnd.n4055 585
R3246 gnd.n3936 gnd.n3935 585
R3247 gnd.n4061 gnd.n4060 585
R3248 gnd.n4063 gnd.n3934 585
R3249 gnd.n4068 gnd.n4065 585
R3250 gnd.n3932 gnd.n3931 585
R3251 gnd.n4073 gnd.n4072 585
R3252 gnd.n4075 gnd.n3930 585
R3253 gnd.n4078 gnd.n4077 585
R3254 gnd.n3928 gnd.n3927 585
R3255 gnd.n4083 gnd.n4082 585
R3256 gnd.n4085 gnd.n3926 585
R3257 gnd.n4088 gnd.n4087 585
R3258 gnd.n3924 gnd.n3923 585
R3259 gnd.n4093 gnd.n4092 585
R3260 gnd.n4095 gnd.n3922 585
R3261 gnd.n4098 gnd.n4097 585
R3262 gnd.n3920 gnd.n3919 585
R3263 gnd.n4103 gnd.n4102 585
R3264 gnd.n4105 gnd.n3918 585
R3265 gnd.n4108 gnd.n4107 585
R3266 gnd.n3916 gnd.n3915 585
R3267 gnd.n4114 gnd.n4113 585
R3268 gnd.n4116 gnd.n3914 585
R3269 gnd.n4117 gnd.n3913 585
R3270 gnd.n4120 gnd.n4119 585
R3271 gnd.n2781 gnd.n2780 585
R3272 gnd.n2787 gnd.n2786 585
R3273 gnd.n2789 gnd.n2788 585
R3274 gnd.n2791 gnd.n2790 585
R3275 gnd.n2793 gnd.n2792 585
R3276 gnd.n2795 gnd.n2794 585
R3277 gnd.n2797 gnd.n2796 585
R3278 gnd.n2799 gnd.n2798 585
R3279 gnd.n2801 gnd.n2800 585
R3280 gnd.n2803 gnd.n2802 585
R3281 gnd.n2805 gnd.n2804 585
R3282 gnd.n2807 gnd.n2806 585
R3283 gnd.n2809 gnd.n2808 585
R3284 gnd.n2811 gnd.n2810 585
R3285 gnd.n2813 gnd.n2812 585
R3286 gnd.n2815 gnd.n2814 585
R3287 gnd.n2817 gnd.n2816 585
R3288 gnd.n2819 gnd.n2818 585
R3289 gnd.n2821 gnd.n2820 585
R3290 gnd.n2824 gnd.n2823 585
R3291 gnd.n2822 gnd.n2760 585
R3292 gnd.n2829 gnd.n2828 585
R3293 gnd.n2831 gnd.n2830 585
R3294 gnd.n2833 gnd.n2832 585
R3295 gnd.n2835 gnd.n2834 585
R3296 gnd.n2837 gnd.n2836 585
R3297 gnd.n2839 gnd.n2838 585
R3298 gnd.n2841 gnd.n2840 585
R3299 gnd.n2843 gnd.n2842 585
R3300 gnd.n2846 gnd.n2845 585
R3301 gnd.n2844 gnd.n2751 585
R3302 gnd.n6036 gnd.n6035 585
R3303 gnd.n6038 gnd.n6037 585
R3304 gnd.n6040 gnd.n6039 585
R3305 gnd.n6042 gnd.n6041 585
R3306 gnd.n6044 gnd.n6043 585
R3307 gnd.n6046 gnd.n6045 585
R3308 gnd.n6048 gnd.n6047 585
R3309 gnd.n6050 gnd.n6049 585
R3310 gnd.n6053 gnd.n6052 585
R3311 gnd.n6055 gnd.n6054 585
R3312 gnd.n6057 gnd.n6056 585
R3313 gnd.n6059 gnd.n6058 585
R3314 gnd.n6061 gnd.n6060 585
R3315 gnd.n6063 gnd.n6062 585
R3316 gnd.n6065 gnd.n6064 585
R3317 gnd.n6067 gnd.n6066 585
R3318 gnd.n6069 gnd.n6068 585
R3319 gnd.n6071 gnd.n6070 585
R3320 gnd.n6073 gnd.n6072 585
R3321 gnd.n6075 gnd.n6074 585
R3322 gnd.n6077 gnd.n6076 585
R3323 gnd.n6079 gnd.n6078 585
R3324 gnd.n6080 gnd.n2720 585
R3325 gnd.n6082 gnd.n6081 585
R3326 gnd.n2721 gnd.n2719 585
R3327 gnd.n2722 gnd.n2570 585
R3328 gnd.n6084 gnd.n2570 585
R3329 gnd.n6163 gnd.n2572 585
R3330 gnd.n6167 gnd.n2572 585
R3331 gnd.n6162 gnd.n6161 585
R3332 gnd.n6161 gnd.n6160 585
R3333 gnd.n2578 gnd.n2562 585
R3334 gnd.n6173 gnd.n2562 585
R3335 gnd.n4313 gnd.n4312 585
R3336 gnd.n4314 gnd.n4313 585
R3337 gnd.n4311 gnd.n2552 585
R3338 gnd.n6179 gnd.n2552 585
R3339 gnd.n4310 gnd.n4309 585
R3340 gnd.n4309 gnd.n4308 585
R3341 gnd.n4306 gnd.n2541 585
R3342 gnd.n6185 gnd.n2541 585
R3343 gnd.n4305 gnd.n4304 585
R3344 gnd.n4304 gnd.n4303 585
R3345 gnd.n4301 gnd.n2532 585
R3346 gnd.n6191 gnd.n2532 585
R3347 gnd.n4300 gnd.n4299 585
R3348 gnd.n4299 gnd.n4298 585
R3349 gnd.n4296 gnd.n2521 585
R3350 gnd.n6197 gnd.n2521 585
R3351 gnd.n4295 gnd.n3769 585
R3352 gnd.n4331 gnd.n3769 585
R3353 gnd.n4294 gnd.n2512 585
R3354 gnd.n6203 gnd.n2512 585
R3355 gnd.n4293 gnd.n4292 585
R3356 gnd.n4292 gnd.n4291 585
R3357 gnd.n3779 gnd.n2501 585
R3358 gnd.n6209 gnd.n2501 585
R3359 gnd.n4247 gnd.n3784 585
R3360 gnd.n4283 gnd.n3784 585
R3361 gnd.n4248 gnd.n2492 585
R3362 gnd.n6215 gnd.n2492 585
R3363 gnd.n4250 gnd.n4249 585
R3364 gnd.n4251 gnd.n4250 585
R3365 gnd.n4245 gnd.n2484 585
R3366 gnd.n6222 gnd.n2484 585
R3367 gnd.n4244 gnd.n4243 585
R3368 gnd.n4243 gnd.n4242 585
R3369 gnd.n4230 gnd.n2475 585
R3370 gnd.n6228 gnd.n2475 585
R3371 gnd.n4229 gnd.n4228 585
R3372 gnd.n4228 gnd.n4227 585
R3373 gnd.n4225 gnd.n2467 585
R3374 gnd.n6235 gnd.n2467 585
R3375 gnd.n4224 gnd.n3800 585
R3376 gnd.n4264 gnd.n3800 585
R3377 gnd.n4223 gnd.n2458 585
R3378 gnd.n6241 gnd.n2458 585
R3379 gnd.n4222 gnd.n4221 585
R3380 gnd.n4221 gnd.n4220 585
R3381 gnd.n3808 gnd.n2449 585
R3382 gnd.n6248 gnd.n2449 585
R3383 gnd.n4210 gnd.n4209 585
R3384 gnd.n4211 gnd.n4210 585
R3385 gnd.n4208 gnd.n2439 585
R3386 gnd.n6254 gnd.n2439 585
R3387 gnd.n4207 gnd.n4206 585
R3388 gnd.n4206 gnd.n4205 585
R3389 gnd.n3813 gnd.n2428 585
R3390 gnd.n6260 gnd.n2428 585
R3391 gnd.n4136 gnd.n3818 585
R3392 gnd.n4197 gnd.n3818 585
R3393 gnd.n4137 gnd.n2419 585
R3394 gnd.n6266 gnd.n2419 585
R3395 gnd.n4144 gnd.n4143 585
R3396 gnd.n4143 gnd.n4142 585
R3397 gnd.n4145 gnd.n2408 585
R3398 gnd.n6272 gnd.n2408 585
R3399 gnd.n4147 gnd.n4146 585
R3400 gnd.n4148 gnd.n4147 585
R3401 gnd.n4129 gnd.n2398 585
R3402 gnd.n6278 gnd.n2398 585
R3403 gnd.n4156 gnd.n4155 585
R3404 gnd.n4155 gnd.n4154 585
R3405 gnd.n4157 gnd.n2387 585
R3406 gnd.n6284 gnd.n2387 585
R3407 gnd.n4159 gnd.n4158 585
R3408 gnd.n4160 gnd.n4159 585
R3409 gnd.n4127 gnd.n2375 585
R3410 gnd.n6290 gnd.n2375 585
R3411 gnd.n4126 gnd.n3834 585
R3412 gnd.n4166 gnd.n3834 585
R3413 gnd.n3840 gnd.n2364 585
R3414 gnd.n6296 gnd.n2364 585
R3415 gnd.n7487 gnd.n7486 585
R3416 gnd.n7486 gnd.n7485 585
R3417 gnd.n7488 gnd.n162 585
R3418 gnd.n7478 gnd.n162 585
R3419 gnd.n7490 gnd.n7489 585
R3420 gnd.n7491 gnd.n7490 585
R3421 gnd.n148 gnd.n147 585
R3422 gnd.n5731 gnd.n148 585
R3423 gnd.n7499 gnd.n7498 585
R3424 gnd.n7498 gnd.n7497 585
R3425 gnd.n7500 gnd.n142 585
R3426 gnd.n5737 gnd.n142 585
R3427 gnd.n7502 gnd.n7501 585
R3428 gnd.n7503 gnd.n7502 585
R3429 gnd.n127 gnd.n126 585
R3430 gnd.n5743 gnd.n127 585
R3431 gnd.n7511 gnd.n7510 585
R3432 gnd.n7510 gnd.n7509 585
R3433 gnd.n7512 gnd.n121 585
R3434 gnd.n5749 gnd.n121 585
R3435 gnd.n7514 gnd.n7513 585
R3436 gnd.n7515 gnd.n7514 585
R3437 gnd.n107 gnd.n106 585
R3438 gnd.n5755 gnd.n107 585
R3439 gnd.n7523 gnd.n7522 585
R3440 gnd.n7522 gnd.n7521 585
R3441 gnd.n7524 gnd.n102 585
R3442 gnd.n5712 gnd.n102 585
R3443 gnd.n7526 gnd.n7525 585
R3444 gnd.n7527 gnd.n7526 585
R3445 gnd.n85 gnd.n83 585
R3446 gnd.n5703 gnd.n85 585
R3447 gnd.n7535 gnd.n7534 585
R3448 gnd.n7534 gnd.n7533 585
R3449 gnd.n84 gnd.n76 585
R3450 gnd.n5697 gnd.n84 585
R3451 gnd.n7538 gnd.n74 585
R3452 gnd.n5770 gnd.n74 585
R3453 gnd.n7540 gnd.n7539 585
R3454 gnd.n7541 gnd.n7540 585
R3455 gnd.n3126 gnd.n73 585
R3456 gnd.n5687 gnd.n73 585
R3457 gnd.n5778 gnd.n3127 585
R3458 gnd.n5778 gnd.n5777 585
R3459 gnd.n5781 gnd.n5780 585
R3460 gnd.n5782 gnd.n5781 585
R3461 gnd.n5779 gnd.n3125 585
R3462 gnd.n3125 gnd.n3120 585
R3463 gnd.n3109 gnd.n3108 585
R3464 gnd.n3113 gnd.n3108 585
R3465 gnd.n5792 gnd.n3110 585
R3466 gnd.n5792 gnd.n5791 585
R3467 gnd.n5794 gnd.n5793 585
R3468 gnd.n5795 gnd.n5794 585
R3469 gnd.n3094 gnd.n3093 585
R3470 gnd.n5670 gnd.n3094 585
R3471 gnd.n5803 gnd.n5802 585
R3472 gnd.n5802 gnd.n5801 585
R3473 gnd.n5804 gnd.n3088 585
R3474 gnd.n5652 gnd.n3088 585
R3475 gnd.n5806 gnd.n5805 585
R3476 gnd.n5807 gnd.n5806 585
R3477 gnd.n3074 gnd.n3073 585
R3478 gnd.n5645 gnd.n3074 585
R3479 gnd.n5815 gnd.n5814 585
R3480 gnd.n5814 gnd.n5813 585
R3481 gnd.n5816 gnd.n3068 585
R3482 gnd.n5589 gnd.n3068 585
R3483 gnd.n5818 gnd.n5817 585
R3484 gnd.n5819 gnd.n5818 585
R3485 gnd.n3054 gnd.n3053 585
R3486 gnd.n5600 gnd.n3054 585
R3487 gnd.n5827 gnd.n5826 585
R3488 gnd.n5826 gnd.n5825 585
R3489 gnd.n5828 gnd.n3048 585
R3490 gnd.n5580 gnd.n3048 585
R3491 gnd.n5830 gnd.n5829 585
R3492 gnd.n5831 gnd.n5830 585
R3493 gnd.n3031 gnd.n3030 585
R3494 gnd.n5572 gnd.n3031 585
R3495 gnd.n5839 gnd.n5838 585
R3496 gnd.n5838 gnd.n5837 585
R3497 gnd.n5840 gnd.n3026 585
R3498 gnd.n4993 gnd.n3026 585
R3499 gnd.n5842 gnd.n5841 585
R3500 gnd.n5843 gnd.n5842 585
R3501 gnd.n5413 gnd.n3025 585
R3502 gnd.n5418 gnd.n5416 585
R3503 gnd.n5419 gnd.n5412 585
R3504 gnd.n5419 gnd.n3012 585
R3505 gnd.n5422 gnd.n5421 585
R3506 gnd.n5410 gnd.n5409 585
R3507 gnd.n5427 gnd.n5426 585
R3508 gnd.n5429 gnd.n5408 585
R3509 gnd.n5432 gnd.n5431 585
R3510 gnd.n5406 gnd.n5405 585
R3511 gnd.n5437 gnd.n5436 585
R3512 gnd.n5439 gnd.n5404 585
R3513 gnd.n5442 gnd.n5441 585
R3514 gnd.n5402 gnd.n5401 585
R3515 gnd.n5447 gnd.n5446 585
R3516 gnd.n5449 gnd.n5400 585
R3517 gnd.n5452 gnd.n5451 585
R3518 gnd.n5398 gnd.n5397 585
R3519 gnd.n5460 gnd.n5459 585
R3520 gnd.n5462 gnd.n5396 585
R3521 gnd.n5465 gnd.n5464 585
R3522 gnd.n5394 gnd.n5393 585
R3523 gnd.n5470 gnd.n5469 585
R3524 gnd.n5472 gnd.n5392 585
R3525 gnd.n5475 gnd.n5474 585
R3526 gnd.n5390 gnd.n5389 585
R3527 gnd.n5481 gnd.n5480 585
R3528 gnd.n5485 gnd.n3262 585
R3529 gnd.n5488 gnd.n5487 585
R3530 gnd.n3260 gnd.n3259 585
R3531 gnd.n5493 gnd.n5492 585
R3532 gnd.n5495 gnd.n3258 585
R3533 gnd.n5498 gnd.n5497 585
R3534 gnd.n3256 gnd.n3255 585
R3535 gnd.n5503 gnd.n5502 585
R3536 gnd.n5505 gnd.n3254 585
R3537 gnd.n5510 gnd.n5507 585
R3538 gnd.n3252 gnd.n3251 585
R3539 gnd.n5515 gnd.n5514 585
R3540 gnd.n5517 gnd.n3250 585
R3541 gnd.n5520 gnd.n5519 585
R3542 gnd.n3248 gnd.n3247 585
R3543 gnd.n5525 gnd.n5524 585
R3544 gnd.n5527 gnd.n3246 585
R3545 gnd.n5530 gnd.n5529 585
R3546 gnd.n3244 gnd.n3243 585
R3547 gnd.n5535 gnd.n5534 585
R3548 gnd.n5537 gnd.n3242 585
R3549 gnd.n5540 gnd.n5539 585
R3550 gnd.n3240 gnd.n3239 585
R3551 gnd.n5545 gnd.n5544 585
R3552 gnd.n5547 gnd.n3238 585
R3553 gnd.n5550 gnd.n5549 585
R3554 gnd.n3236 gnd.n3235 585
R3555 gnd.n5556 gnd.n5555 585
R3556 gnd.n5558 gnd.n3234 585
R3557 gnd.n5559 gnd.n3233 585
R3558 gnd.n5562 gnd.n5561 585
R3559 gnd.n7347 gnd.n7346 585
R3560 gnd.n7353 gnd.n7352 585
R3561 gnd.n7355 gnd.n7354 585
R3562 gnd.n7357 gnd.n7356 585
R3563 gnd.n7359 gnd.n7358 585
R3564 gnd.n7361 gnd.n7360 585
R3565 gnd.n7363 gnd.n7362 585
R3566 gnd.n7365 gnd.n7364 585
R3567 gnd.n7367 gnd.n7366 585
R3568 gnd.n7369 gnd.n7368 585
R3569 gnd.n7371 gnd.n7370 585
R3570 gnd.n7373 gnd.n7372 585
R3571 gnd.n7375 gnd.n7374 585
R3572 gnd.n7377 gnd.n7376 585
R3573 gnd.n7379 gnd.n7378 585
R3574 gnd.n7381 gnd.n7380 585
R3575 gnd.n7383 gnd.n7382 585
R3576 gnd.n7385 gnd.n7384 585
R3577 gnd.n7387 gnd.n7386 585
R3578 gnd.n7390 gnd.n7389 585
R3579 gnd.n7388 gnd.n7326 585
R3580 gnd.n7395 gnd.n7394 585
R3581 gnd.n7397 gnd.n7396 585
R3582 gnd.n7399 gnd.n7398 585
R3583 gnd.n7401 gnd.n7400 585
R3584 gnd.n7403 gnd.n7402 585
R3585 gnd.n7405 gnd.n7404 585
R3586 gnd.n7407 gnd.n7406 585
R3587 gnd.n7409 gnd.n7408 585
R3588 gnd.n7411 gnd.n7410 585
R3589 gnd.n7413 gnd.n7412 585
R3590 gnd.n7415 gnd.n7414 585
R3591 gnd.n7417 gnd.n7416 585
R3592 gnd.n7419 gnd.n7418 585
R3593 gnd.n7421 gnd.n7420 585
R3594 gnd.n7423 gnd.n7422 585
R3595 gnd.n7425 gnd.n7424 585
R3596 gnd.n7427 gnd.n7426 585
R3597 gnd.n7429 gnd.n7428 585
R3598 gnd.n7431 gnd.n7430 585
R3599 gnd.n7433 gnd.n7432 585
R3600 gnd.n7438 gnd.n7437 585
R3601 gnd.n7440 gnd.n7439 585
R3602 gnd.n7442 gnd.n7441 585
R3603 gnd.n7444 gnd.n7443 585
R3604 gnd.n7446 gnd.n7445 585
R3605 gnd.n7448 gnd.n7447 585
R3606 gnd.n7450 gnd.n7449 585
R3607 gnd.n7452 gnd.n7451 585
R3608 gnd.n7454 gnd.n7453 585
R3609 gnd.n7456 gnd.n7455 585
R3610 gnd.n7458 gnd.n7457 585
R3611 gnd.n7460 gnd.n7459 585
R3612 gnd.n7462 gnd.n7461 585
R3613 gnd.n7464 gnd.n7463 585
R3614 gnd.n7465 gnd.n7286 585
R3615 gnd.n7467 gnd.n7466 585
R3616 gnd.n7287 gnd.n7285 585
R3617 gnd.n7288 gnd.n167 585
R3618 gnd.n7469 gnd.n167 585
R3619 gnd.n7481 gnd.n169 585
R3620 gnd.n7485 gnd.n169 585
R3621 gnd.n7480 gnd.n7479 585
R3622 gnd.n7479 gnd.n7478 585
R3623 gnd.n175 gnd.n160 585
R3624 gnd.n7491 gnd.n160 585
R3625 gnd.n5733 gnd.n5732 585
R3626 gnd.n5732 gnd.n5731 585
R3627 gnd.n5734 gnd.n150 585
R3628 gnd.n7497 gnd.n150 585
R3629 gnd.n5736 gnd.n5735 585
R3630 gnd.n5737 gnd.n5736 585
R3631 gnd.n5719 gnd.n139 585
R3632 gnd.n7503 gnd.n139 585
R3633 gnd.n5745 gnd.n5744 585
R3634 gnd.n5744 gnd.n5743 585
R3635 gnd.n5746 gnd.n129 585
R3636 gnd.n7509 gnd.n129 585
R3637 gnd.n5748 gnd.n5747 585
R3638 gnd.n5749 gnd.n5748 585
R3639 gnd.n5717 gnd.n118 585
R3640 gnd.n7515 gnd.n118 585
R3641 gnd.n5716 gnd.n3191 585
R3642 gnd.n5755 gnd.n3191 585
R3643 gnd.n5715 gnd.n109 585
R3644 gnd.n7521 gnd.n109 585
R3645 gnd.n5714 gnd.n5713 585
R3646 gnd.n5713 gnd.n5712 585
R3647 gnd.n3197 gnd.n99 585
R3648 gnd.n7527 gnd.n99 585
R3649 gnd.n5702 gnd.n5701 585
R3650 gnd.n5703 gnd.n5702 585
R3651 gnd.n5700 gnd.n87 585
R3652 gnd.n7533 gnd.n87 585
R3653 gnd.n5699 gnd.n5698 585
R3654 gnd.n5698 gnd.n5697 585
R3655 gnd.n5691 gnd.n3137 585
R3656 gnd.n5770 gnd.n3137 585
R3657 gnd.n5690 gnd.n70 585
R3658 gnd.n7541 gnd.n70 585
R3659 gnd.n5689 gnd.n5688 585
R3660 gnd.n5688 gnd.n5687 585
R3661 gnd.n5686 gnd.n3128 585
R3662 gnd.n5777 gnd.n3128 585
R3663 gnd.n5685 gnd.n3121 585
R3664 gnd.n5782 gnd.n3121 585
R3665 gnd.n5675 gnd.n3202 585
R3666 gnd.n5675 gnd.n3120 585
R3667 gnd.n5677 gnd.n5676 585
R3668 gnd.n5676 gnd.n3113 585
R3669 gnd.n5674 gnd.n3111 585
R3670 gnd.n5791 gnd.n3111 585
R3671 gnd.n5673 gnd.n3105 585
R3672 gnd.n5795 gnd.n3105 585
R3673 gnd.n5672 gnd.n5671 585
R3674 gnd.n5671 gnd.n5670 585
R3675 gnd.n3204 gnd.n3096 585
R3676 gnd.n5801 gnd.n3096 585
R3677 gnd.n5651 gnd.n5650 585
R3678 gnd.n5652 gnd.n5651 585
R3679 gnd.n5648 gnd.n3085 585
R3680 gnd.n5807 gnd.n3085 585
R3681 gnd.n5647 gnd.n5646 585
R3682 gnd.n5646 gnd.n5645 585
R3683 gnd.n3210 gnd.n3076 585
R3684 gnd.n5813 gnd.n3076 585
R3685 gnd.n5588 gnd.n5587 585
R3686 gnd.n5589 gnd.n5588 585
R3687 gnd.n5585 gnd.n3065 585
R3688 gnd.n5819 gnd.n3065 585
R3689 gnd.n5584 gnd.n3217 585
R3690 gnd.n5600 gnd.n3217 585
R3691 gnd.n5583 gnd.n3056 585
R3692 gnd.n5825 gnd.n3056 585
R3693 gnd.n5582 gnd.n5581 585
R3694 gnd.n5581 gnd.n5580 585
R3695 gnd.n3222 gnd.n3045 585
R3696 gnd.n5831 gnd.n3045 585
R3697 gnd.n5571 gnd.n5570 585
R3698 gnd.n5572 gnd.n5571 585
R3699 gnd.n5569 gnd.n3033 585
R3700 gnd.n5837 gnd.n3033 585
R3701 gnd.n5568 gnd.n3228 585
R3702 gnd.n4993 gnd.n3228 585
R3703 gnd.n3227 gnd.n3021 585
R3704 gnd.n5843 gnd.n3021 585
R3705 gnd.n6327 gnd.n871 585
R3706 gnd.n2339 gnd.n871 585
R3707 gnd.n7231 gnd.n7230 585
R3708 gnd.n7232 gnd.n7231 585
R3709 gnd.n267 gnd.n266 585
R3710 gnd.n7233 gnd.n267 585
R3711 gnd.n7236 gnd.n7235 585
R3712 gnd.n7235 gnd.n7234 585
R3713 gnd.n7237 gnd.n261 585
R3714 gnd.n261 gnd.n260 585
R3715 gnd.n7239 gnd.n7238 585
R3716 gnd.n7240 gnd.n7239 585
R3717 gnd.n259 gnd.n258 585
R3718 gnd.n7241 gnd.n259 585
R3719 gnd.n7244 gnd.n7243 585
R3720 gnd.n7243 gnd.n7242 585
R3721 gnd.n7245 gnd.n253 585
R3722 gnd.n253 gnd.n252 585
R3723 gnd.n7247 gnd.n7246 585
R3724 gnd.n7248 gnd.n7247 585
R3725 gnd.n251 gnd.n250 585
R3726 gnd.n7249 gnd.n251 585
R3727 gnd.n7252 gnd.n7251 585
R3728 gnd.n7251 gnd.n7250 585
R3729 gnd.n7253 gnd.n245 585
R3730 gnd.n245 gnd.n243 585
R3731 gnd.n7255 gnd.n7254 585
R3732 gnd.n7256 gnd.n7255 585
R3733 gnd.n246 gnd.n244 585
R3734 gnd.n244 gnd.n184 585
R3735 gnd.n3174 gnd.n3173 585
R3736 gnd.n3173 gnd.n171 585
R3737 gnd.n3175 gnd.n3167 585
R3738 gnd.n3167 gnd.n168 585
R3739 gnd.n3177 gnd.n3176 585
R3740 gnd.n3177 gnd.n176 585
R3741 gnd.n3178 gnd.n3166 585
R3742 gnd.n3178 gnd.n159 585
R3743 gnd.n3180 gnd.n3179 585
R3744 gnd.n3179 gnd.n152 585
R3745 gnd.n3181 gnd.n3161 585
R3746 gnd.n3161 gnd.n149 585
R3747 gnd.n3183 gnd.n3182 585
R3748 gnd.n3183 gnd.n141 585
R3749 gnd.n3184 gnd.n3160 585
R3750 gnd.n3184 gnd.n138 585
R3751 gnd.n3186 gnd.n3185 585
R3752 gnd.n3185 gnd.n131 585
R3753 gnd.n3187 gnd.n3155 585
R3754 gnd.n3155 gnd.n128 585
R3755 gnd.n3189 gnd.n3188 585
R3756 gnd.n3189 gnd.n120 585
R3757 gnd.n3190 gnd.n3154 585
R3758 gnd.n3190 gnd.n117 585
R3759 gnd.n5758 gnd.n5757 585
R3760 gnd.n5757 gnd.n5756 585
R3761 gnd.n5759 gnd.n3149 585
R3762 gnd.n3149 gnd.n108 585
R3763 gnd.n5761 gnd.n5760 585
R3764 gnd.n5761 gnd.n101 585
R3765 gnd.n5762 gnd.n3148 585
R3766 gnd.n5762 gnd.n98 585
R3767 gnd.n5764 gnd.n5763 585
R3768 gnd.n5763 gnd.n89 585
R3769 gnd.n5765 gnd.n3139 585
R3770 gnd.n3139 gnd.n86 585
R3771 gnd.n5768 gnd.n5767 585
R3772 gnd.n5769 gnd.n5768 585
R3773 gnd.n3146 gnd.n3138 585
R3774 gnd.n3138 gnd.n71 585
R3775 gnd.n3144 gnd.n3143 585
R3776 gnd.n3143 gnd.n69 585
R3777 gnd.n3142 gnd.n3141 585
R3778 gnd.n3142 gnd.n3130 585
R3779 gnd.n3118 gnd.n3117 585
R3780 gnd.n3123 gnd.n3118 585
R3781 gnd.n5785 gnd.n5784 585
R3782 gnd.n5784 gnd.n5783 585
R3783 gnd.n5787 gnd.n3115 585
R3784 gnd.n3119 gnd.n3115 585
R3785 gnd.n5789 gnd.n5788 585
R3786 gnd.n5790 gnd.n5789 585
R3787 gnd.n5635 gnd.n3114 585
R3788 gnd.n3114 gnd.n3107 585
R3789 gnd.n5637 gnd.n5636 585
R3790 gnd.n5637 gnd.n3104 585
R3791 gnd.n5638 gnd.n5632 585
R3792 gnd.n5638 gnd.n3205 585
R3793 gnd.n5640 gnd.n5639 585
R3794 gnd.n5639 gnd.n3095 585
R3795 gnd.n5641 gnd.n3213 585
R3796 gnd.n3213 gnd.n3087 585
R3797 gnd.n5643 gnd.n5642 585
R3798 gnd.n5644 gnd.n5643 585
R3799 gnd.n3214 gnd.n3212 585
R3800 gnd.n3212 gnd.n3078 585
R3801 gnd.n5626 gnd.n5625 585
R3802 gnd.n5625 gnd.n3075 585
R3803 gnd.n5624 gnd.n3216 585
R3804 gnd.n5624 gnd.n3067 585
R3805 gnd.n5623 gnd.n5622 585
R3806 gnd.n5623 gnd.n3064 585
R3807 gnd.n5603 gnd.n5602 585
R3808 gnd.n5602 gnd.n5601 585
R3809 gnd.n5618 gnd.n5617 585
R3810 gnd.n5617 gnd.n3055 585
R3811 gnd.n5616 gnd.n5605 585
R3812 gnd.n5616 gnd.n3047 585
R3813 gnd.n5615 gnd.n5614 585
R3814 gnd.n5615 gnd.n3044 585
R3815 gnd.n5607 gnd.n5606 585
R3816 gnd.n5606 gnd.n3035 585
R3817 gnd.n5610 gnd.n5609 585
R3818 gnd.n5609 gnd.n3032 585
R3819 gnd.n3019 gnd.n3018 585
R3820 gnd.n3023 gnd.n3019 585
R3821 gnd.n5846 gnd.n5845 585
R3822 gnd.n5845 gnd.n5844 585
R3823 gnd.n5847 gnd.n3013 585
R3824 gnd.n3020 gnd.n3013 585
R3825 gnd.n5849 gnd.n5848 585
R3826 gnd.n5850 gnd.n5849 585
R3827 gnd.n3010 gnd.n3009 585
R3828 gnd.n5851 gnd.n3010 585
R3829 gnd.n5854 gnd.n5853 585
R3830 gnd.n5853 gnd.n5852 585
R3831 gnd.n5855 gnd.n3004 585
R3832 gnd.n3004 gnd.n3002 585
R3833 gnd.n5857 gnd.n5856 585
R3834 gnd.n5858 gnd.n5857 585
R3835 gnd.n3005 gnd.n3003 585
R3836 gnd.n3003 gnd.n3000 585
R3837 gnd.n5179 gnd.n5178 585
R3838 gnd.n5180 gnd.n5179 585
R3839 gnd.n3354 gnd.n3353 585
R3840 gnd.n5182 gnd.n3354 585
R3841 gnd.n5187 gnd.n5186 585
R3842 gnd.n5186 gnd.n5185 585
R3843 gnd.n5188 gnd.n3348 585
R3844 gnd.n3355 gnd.n3348 585
R3845 gnd.n5190 gnd.n5189 585
R3846 gnd.n5191 gnd.n5190 585
R3847 gnd.n3342 gnd.n3341 585
R3848 gnd.n5193 gnd.n3342 585
R3849 gnd.n5198 gnd.n5197 585
R3850 gnd.n5197 gnd.n5196 585
R3851 gnd.n5199 gnd.n3336 585
R3852 gnd.n3343 gnd.n3336 585
R3853 gnd.n5201 gnd.n5200 585
R3854 gnd.n5202 gnd.n5201 585
R3855 gnd.n3330 gnd.n3329 585
R3856 gnd.n5204 gnd.n3330 585
R3857 gnd.n5209 gnd.n5208 585
R3858 gnd.n5208 gnd.n5207 585
R3859 gnd.n5210 gnd.n3324 585
R3860 gnd.n3331 gnd.n3324 585
R3861 gnd.n5212 gnd.n5211 585
R3862 gnd.n5213 gnd.n5212 585
R3863 gnd.n3320 gnd.n3319 585
R3864 gnd.n5215 gnd.n3320 585
R3865 gnd.n5220 gnd.n5219 585
R3866 gnd.n5219 gnd.n5218 585
R3867 gnd.n5221 gnd.n3314 585
R3868 gnd.n3314 gnd.n3305 585
R3869 gnd.n5223 gnd.n5222 585
R3870 gnd.n5224 gnd.n5223 585
R3871 gnd.n3315 gnd.n3313 585
R3872 gnd.n3313 gnd.n3310 585
R3873 gnd.n4933 gnd.n4932 585
R3874 gnd.n4932 gnd.n3372 585
R3875 gnd.n4934 gnd.n3388 585
R3876 gnd.n3388 gnd.n3376 585
R3877 gnd.n4936 gnd.n4935 585
R3878 gnd.n4937 gnd.n4936 585
R3879 gnd.n3389 gnd.n3387 585
R3880 gnd.n3396 gnd.n3387 585
R3881 gnd.n4925 gnd.n4924 585
R3882 gnd.n4924 gnd.n4923 585
R3883 gnd.n3392 gnd.n3391 585
R3884 gnd.n4827 gnd.n3392 585
R3885 gnd.n4885 gnd.n3416 585
R3886 gnd.n3416 gnd.n3409 585
R3887 gnd.n4887 gnd.n4886 585
R3888 gnd.n4888 gnd.n4887 585
R3889 gnd.n3417 gnd.n3415 585
R3890 gnd.n3415 gnd.n3413 585
R3891 gnd.n4880 gnd.n4879 585
R3892 gnd.n4879 gnd.n4878 585
R3893 gnd.n3420 gnd.n3419 585
R3894 gnd.n4870 gnd.n3420 585
R3895 gnd.n4856 gnd.n4855 585
R3896 gnd.n4857 gnd.n4856 585
R3897 gnd.n3439 gnd.n3438 585
R3898 gnd.n4807 gnd.n3438 585
R3899 gnd.n4851 gnd.n4850 585
R3900 gnd.n4850 gnd.n4849 585
R3901 gnd.n3442 gnd.n3441 585
R3902 gnd.n3450 gnd.n3442 585
R3903 gnd.n4796 gnd.n4795 585
R3904 gnd.n4797 gnd.n4796 585
R3905 gnd.n3459 gnd.n3458 585
R3906 gnd.n3458 gnd.n3455 585
R3907 gnd.n4791 gnd.n4790 585
R3908 gnd.n4790 gnd.n4789 585
R3909 gnd.n3462 gnd.n3461 585
R3910 gnd.n3468 gnd.n3462 585
R3911 gnd.n4771 gnd.n4770 585
R3912 gnd.n4772 gnd.n4771 585
R3913 gnd.n3478 gnd.n3477 585
R3914 gnd.n3485 gnd.n3477 585
R3915 gnd.n4766 gnd.n4765 585
R3916 gnd.n4765 gnd.n4764 585
R3917 gnd.n3481 gnd.n3480 585
R3918 gnd.n3489 gnd.n3481 585
R3919 gnd.n4715 gnd.n4714 585
R3920 gnd.n4716 gnd.n4715 585
R3921 gnd.n3500 gnd.n3499 585
R3922 gnd.n3518 gnd.n3499 585
R3923 gnd.n4710 gnd.n4709 585
R3924 gnd.n4709 gnd.n4708 585
R3925 gnd.n3503 gnd.n3502 585
R3926 gnd.n3511 gnd.n3503 585
R3927 gnd.n4675 gnd.n4674 585
R3928 gnd.n4676 gnd.n4675 585
R3929 gnd.n3523 gnd.n3522 585
R3930 gnd.n3538 gnd.n3522 585
R3931 gnd.n4670 gnd.n4669 585
R3932 gnd.n4669 gnd.n4668 585
R3933 gnd.n3526 gnd.n3525 585
R3934 gnd.n4658 gnd.n3526 585
R3935 gnd.n4624 gnd.n3555 585
R3936 gnd.n3555 gnd.n3547 585
R3937 gnd.n4626 gnd.n4625 585
R3938 gnd.n4627 gnd.n4626 585
R3939 gnd.n3556 gnd.n3554 585
R3940 gnd.n3554 gnd.n3551 585
R3941 gnd.n4619 gnd.n4618 585
R3942 gnd.n4618 gnd.n4617 585
R3943 gnd.n3559 gnd.n3558 585
R3944 gnd.n3565 gnd.n3559 585
R3945 gnd.n4597 gnd.n4596 585
R3946 gnd.n4598 gnd.n4597 585
R3947 gnd.n3574 gnd.n3573 585
R3948 gnd.n3580 gnd.n3573 585
R3949 gnd.n4592 gnd.n4591 585
R3950 gnd.n4591 gnd.n4590 585
R3951 gnd.n3577 gnd.n3576 585
R3952 gnd.n3584 gnd.n3577 585
R3953 gnd.n4535 gnd.n3599 585
R3954 gnd.n3599 gnd.n3589 585
R3955 gnd.n4537 gnd.n4536 585
R3956 gnd.n4538 gnd.n4537 585
R3957 gnd.n3600 gnd.n3598 585
R3958 gnd.n4512 gnd.n3598 585
R3959 gnd.n4530 gnd.n4529 585
R3960 gnd.n4529 gnd.n4528 585
R3961 gnd.n3603 gnd.n3602 585
R3962 gnd.n4502 gnd.n3603 585
R3963 gnd.n4465 gnd.n4464 585
R3964 gnd.n4465 gnd.n2911 585
R3965 gnd.n4467 gnd.n4461 585
R3966 gnd.n4467 gnd.n4466 585
R3967 gnd.n4469 gnd.n4468 585
R3968 gnd.n4468 gnd.n3681 585
R3969 gnd.n4470 gnd.n3693 585
R3970 gnd.n3693 gnd.n3680 585
R3971 gnd.n4472 gnd.n4471 585
R3972 gnd.n4473 gnd.n4472 585
R3973 gnd.n3694 gnd.n3692 585
R3974 gnd.n3692 gnd.n3689 585
R3975 gnd.n4455 gnd.n4454 585
R3976 gnd.n4454 gnd.n4453 585
R3977 gnd.n3697 gnd.n3696 585
R3978 gnd.n3706 gnd.n3697 585
R3979 gnd.n4430 gnd.n3718 585
R3980 gnd.n3718 gnd.n3705 585
R3981 gnd.n4432 gnd.n4431 585
R3982 gnd.n4433 gnd.n4432 585
R3983 gnd.n3719 gnd.n3717 585
R3984 gnd.n3717 gnd.n3714 585
R3985 gnd.n4425 gnd.n4424 585
R3986 gnd.n4424 gnd.n4423 585
R3987 gnd.n3722 gnd.n3721 585
R3988 gnd.n3730 gnd.n3722 585
R3989 gnd.n4400 gnd.n3743 585
R3990 gnd.n3743 gnd.n3729 585
R3991 gnd.n4402 gnd.n4401 585
R3992 gnd.n4403 gnd.n4402 585
R3993 gnd.n3744 gnd.n3742 585
R3994 gnd.n3742 gnd.n3739 585
R3995 gnd.n4395 gnd.n4394 585
R3996 gnd.n4394 gnd.n4393 585
R3997 gnd.n3747 gnd.n3746 585
R3998 gnd.n4375 gnd.n3747 585
R3999 gnd.n4372 gnd.n4371 585
R4000 gnd.n4373 gnd.n4372 585
R4001 gnd.n3749 gnd.n3748 585
R4002 gnd.n3748 gnd.n2601 585
R4003 gnd.n4367 gnd.n4366 585
R4004 gnd.n4366 gnd.n2587 585
R4005 gnd.n4365 gnd.n3751 585
R4006 gnd.n4365 gnd.n4364 585
R4007 gnd.n4363 gnd.n4362 585
R4008 gnd.n4363 gnd.n2690 585
R4009 gnd.n3753 gnd.n3752 585
R4010 gnd.n3752 gnd.n2676 585
R4011 gnd.n4358 gnd.n4357 585
R4012 gnd.n4357 gnd.n2574 585
R4013 gnd.n4356 gnd.n3755 585
R4014 gnd.n4356 gnd.n2571 585
R4015 gnd.n4355 gnd.n4354 585
R4016 gnd.n4355 gnd.n2564 585
R4017 gnd.n3757 gnd.n3756 585
R4018 gnd.n3756 gnd.n2561 585
R4019 gnd.n4350 gnd.n4349 585
R4020 gnd.n4349 gnd.n2554 585
R4021 gnd.n4348 gnd.n3759 585
R4022 gnd.n4348 gnd.n2551 585
R4023 gnd.n4347 gnd.n4346 585
R4024 gnd.n4347 gnd.n2543 585
R4025 gnd.n3761 gnd.n3760 585
R4026 gnd.n4302 gnd.n3760 585
R4027 gnd.n4342 gnd.n4341 585
R4028 gnd.n4341 gnd.n2534 585
R4029 gnd.n4340 gnd.n3763 585
R4030 gnd.n4340 gnd.n2531 585
R4031 gnd.n4339 gnd.n4338 585
R4032 gnd.n4339 gnd.n2523 585
R4033 gnd.n3765 gnd.n3764 585
R4034 gnd.n3764 gnd.n2520 585
R4035 gnd.n4334 gnd.n4333 585
R4036 gnd.n4333 gnd.n4332 585
R4037 gnd.n3768 gnd.n3767 585
R4038 gnd.n3768 gnd.n2511 585
R4039 gnd.n4279 gnd.n3786 585
R4040 gnd.n3786 gnd.n2503 585
R4041 gnd.n4281 gnd.n4280 585
R4042 gnd.n4282 gnd.n4281 585
R4043 gnd.n3787 gnd.n3785 585
R4044 gnd.n3785 gnd.n2494 585
R4045 gnd.n4233 gnd.n4232 585
R4046 gnd.n4233 gnd.n2491 585
R4047 gnd.n4235 gnd.n4234 585
R4048 gnd.n4234 gnd.n2486 585
R4049 gnd.n4237 gnd.n4236 585
R4050 gnd.n4237 gnd.n2483 585
R4051 gnd.n4240 gnd.n4239 585
R4052 gnd.n4241 gnd.n4240 585
R4053 gnd.n4238 gnd.n4231 585
R4054 gnd.n4231 gnd.n2474 585
R4055 gnd.n3798 gnd.n3797 585
R4056 gnd.n3797 gnd.n2469 585
R4057 gnd.n4266 gnd.n3799 585
R4058 gnd.n4266 gnd.n4265 585
R4059 gnd.n4268 gnd.n4267 585
R4060 gnd.n4267 gnd.n2460 585
R4061 gnd.n4270 gnd.n4269 585
R4062 gnd.n4270 gnd.n2457 585
R4063 gnd.n4271 gnd.n3795 585
R4064 gnd.n4271 gnd.n2451 585
R4065 gnd.n4273 gnd.n4272 585
R4066 gnd.n4272 gnd.n2448 585
R4067 gnd.n3796 gnd.n3794 585
R4068 gnd.n3796 gnd.n2441 585
R4069 gnd.n4192 gnd.n4191 585
R4070 gnd.n4191 gnd.n2438 585
R4071 gnd.n4193 gnd.n3820 585
R4072 gnd.n3820 gnd.n2430 585
R4073 gnd.n4195 gnd.n4194 585
R4074 gnd.n4196 gnd.n4195 585
R4075 gnd.n3821 gnd.n3819 585
R4076 gnd.n3819 gnd.n2421 585
R4077 gnd.n4185 gnd.n4184 585
R4078 gnd.n4184 gnd.n2418 585
R4079 gnd.n4183 gnd.n3823 585
R4080 gnd.n4183 gnd.n2410 585
R4081 gnd.n4182 gnd.n4181 585
R4082 gnd.n4182 gnd.n2407 585
R4083 gnd.n3825 gnd.n3824 585
R4084 gnd.n3824 gnd.n2400 585
R4085 gnd.n4177 gnd.n4176 585
R4086 gnd.n4176 gnd.n2397 585
R4087 gnd.n4175 gnd.n3827 585
R4088 gnd.n4175 gnd.n2389 585
R4089 gnd.n4174 gnd.n4173 585
R4090 gnd.n4174 gnd.n2386 585
R4091 gnd.n3829 gnd.n3828 585
R4092 gnd.n3828 gnd.n2377 585
R4093 gnd.n4169 gnd.n4168 585
R4094 gnd.n4168 gnd.n4167 585
R4095 gnd.n3833 gnd.n3832 585
R4096 gnd.n3833 gnd.n2366 585
R4097 gnd.n2362 gnd.n2361 585
R4098 gnd.n6297 gnd.n2362 585
R4099 gnd.n6300 gnd.n6299 585
R4100 gnd.n6299 gnd.n6298 585
R4101 gnd.n6301 gnd.n2356 585
R4102 gnd.n2356 gnd.n2355 585
R4103 gnd.n6303 gnd.n6302 585
R4104 gnd.n6304 gnd.n6303 585
R4105 gnd.n2354 gnd.n2353 585
R4106 gnd.n6305 gnd.n2354 585
R4107 gnd.n6308 gnd.n6307 585
R4108 gnd.n6307 gnd.n6306 585
R4109 gnd.n6309 gnd.n2348 585
R4110 gnd.n2348 gnd.n2347 585
R4111 gnd.n6311 gnd.n6310 585
R4112 gnd.n6312 gnd.n6311 585
R4113 gnd.n2346 gnd.n2345 585
R4114 gnd.n6313 gnd.n2346 585
R4115 gnd.n6316 gnd.n6315 585
R4116 gnd.n6315 gnd.n6314 585
R4117 gnd.n6317 gnd.n2341 585
R4118 gnd.n2341 gnd.n2340 585
R4119 gnd.n6319 gnd.n6318 585
R4120 gnd.n6320 gnd.n6319 585
R4121 gnd.n876 gnd.n875 585
R4122 gnd.n6321 gnd.n876 585
R4123 gnd.n6324 gnd.n6323 585
R4124 gnd.n6323 gnd.n6322 585
R4125 gnd.n5861 gnd.n5860 585
R4126 gnd.n5860 gnd.n5859 585
R4127 gnd.n5862 gnd.n2997 585
R4128 gnd.n5174 gnd.n2997 585
R4129 gnd.n5863 gnd.n2996 585
R4130 gnd.n5181 gnd.n2996 585
R4131 gnd.n5183 gnd.n2994 585
R4132 gnd.n5184 gnd.n5183 585
R4133 gnd.n5867 gnd.n2993 585
R4134 gnd.n3356 gnd.n2993 585
R4135 gnd.n5868 gnd.n2992 585
R4136 gnd.n3347 gnd.n2992 585
R4137 gnd.n5869 gnd.n2991 585
R4138 gnd.n5192 gnd.n2991 585
R4139 gnd.n5194 gnd.n2989 585
R4140 gnd.n5195 gnd.n5194 585
R4141 gnd.n5873 gnd.n2988 585
R4142 gnd.n3344 gnd.n2988 585
R4143 gnd.n5874 gnd.n2987 585
R4144 gnd.n3335 gnd.n2987 585
R4145 gnd.n5875 gnd.n2986 585
R4146 gnd.n5203 gnd.n2986 585
R4147 gnd.n5205 gnd.n2984 585
R4148 gnd.n5206 gnd.n5205 585
R4149 gnd.n5879 gnd.n2983 585
R4150 gnd.n3332 gnd.n2983 585
R4151 gnd.n5880 gnd.n2982 585
R4152 gnd.n3323 gnd.n2982 585
R4153 gnd.n5881 gnd.n2981 585
R4154 gnd.n5214 gnd.n2981 585
R4155 gnd.n5216 gnd.n2979 585
R4156 gnd.n5217 gnd.n5216 585
R4157 gnd.n5885 gnd.n2978 585
R4158 gnd.n3267 gnd.n2978 585
R4159 gnd.n5886 gnd.n2977 585
R4160 gnd.n3304 gnd.n2977 585
R4161 gnd.n5887 gnd.n2976 585
R4162 gnd.n5226 gnd.n2976 585
R4163 gnd.n4954 gnd.n2974 585
R4164 gnd.n4955 gnd.n4954 585
R4165 gnd.n5891 gnd.n2973 585
R4166 gnd.n3378 gnd.n2973 585
R4167 gnd.n5892 gnd.n2972 585
R4168 gnd.n3386 gnd.n2972 585
R4169 gnd.n5893 gnd.n2971 585
R4170 gnd.n3383 gnd.n2971 585
R4171 gnd.n4921 gnd.n2969 585
R4172 gnd.n4922 gnd.n4921 585
R4173 gnd.n5897 gnd.n2968 585
R4174 gnd.n4913 gnd.n2968 585
R4175 gnd.n5898 gnd.n2967 585
R4176 gnd.n4828 gnd.n2967 585
R4177 gnd.n5899 gnd.n2966 585
R4178 gnd.n4898 gnd.n2966 585
R4179 gnd.n4889 gnd.n2964 585
R4180 gnd.n4890 gnd.n4889 585
R4181 gnd.n5903 gnd.n2963 585
R4182 gnd.n3422 gnd.n2963 585
R4183 gnd.n5904 gnd.n2962 585
R4184 gnd.n4868 gnd.n2962 585
R4185 gnd.n5905 gnd.n2961 585
R4186 gnd.n3426 gnd.n2961 585
R4187 gnd.n4858 gnd.n2959 585
R4188 gnd.n4859 gnd.n4858 585
R4189 gnd.n5909 gnd.n2958 585
R4190 gnd.n3444 gnd.n2958 585
R4191 gnd.n5910 gnd.n2957 585
R4192 gnd.n4738 gnd.n2957 585
R4193 gnd.n5911 gnd.n2956 585
R4194 gnd.n3449 gnd.n2956 585
R4195 gnd.n4799 gnd.n2954 585
R4196 gnd.n4800 gnd.n4799 585
R4197 gnd.n5915 gnd.n2953 585
R4198 gnd.n4788 gnd.n2953 585
R4199 gnd.n5916 gnd.n2952 585
R4200 gnd.n3469 gnd.n2952 585
R4201 gnd.n5917 gnd.n2951 585
R4202 gnd.n3476 gnd.n2951 585
R4203 gnd.n4729 gnd.n2949 585
R4204 gnd.n4730 gnd.n4729 585
R4205 gnd.n5921 gnd.n2948 585
R4206 gnd.n4763 gnd.n2948 585
R4207 gnd.n5922 gnd.n2947 585
R4208 gnd.n4755 gnd.n2947 585
R4209 gnd.n5923 gnd.n2946 585
R4210 gnd.n4717 gnd.n2946 585
R4211 gnd.n4688 gnd.n2944 585
R4212 gnd.n4689 gnd.n4688 585
R4213 gnd.n5927 gnd.n2943 585
R4214 gnd.n3506 gnd.n2943 585
R4215 gnd.n5928 gnd.n2942 585
R4216 gnd.n4697 gnd.n2942 585
R4217 gnd.n5929 gnd.n2941 585
R4218 gnd.n4677 gnd.n2941 585
R4219 gnd.n4649 gnd.n2939 585
R4220 gnd.n4650 gnd.n4649 585
R4221 gnd.n5933 gnd.n2938 585
R4222 gnd.n3529 gnd.n2938 585
R4223 gnd.n5934 gnd.n2937 585
R4224 gnd.n4641 gnd.n2937 585
R4225 gnd.n5935 gnd.n2936 585
R4226 gnd.n3534 gnd.n2936 585
R4227 gnd.n4637 gnd.n2934 585
R4228 gnd.n4638 gnd.n4637 585
R4229 gnd.n5939 gnd.n2933 585
R4230 gnd.n4629 gnd.n2933 585
R4231 gnd.n5940 gnd.n2932 585
R4232 gnd.n4616 gnd.n2932 585
R4233 gnd.n5941 gnd.n2931 585
R4234 gnd.n3566 gnd.n2931 585
R4235 gnd.n4547 gnd.n2929 585
R4236 gnd.n4548 gnd.n4547 585
R4237 gnd.n5945 gnd.n2928 585
R4238 gnd.n3571 gnd.n2928 585
R4239 gnd.n5946 gnd.n2927 585
R4240 gnd.n4589 gnd.n2927 585
R4241 gnd.n5947 gnd.n2926 585
R4242 gnd.n4581 gnd.n2926 585
R4243 gnd.n4567 gnd.n2924 585
R4244 gnd.n4568 gnd.n4567 585
R4245 gnd.n5951 gnd.n2923 585
R4246 gnd.n4518 gnd.n2923 585
R4247 gnd.n5952 gnd.n2922 585
R4248 gnd.n4539 gnd.n2922 585
R4249 gnd.n5953 gnd.n2921 585
R4250 gnd.n3606 gnd.n2921 585
R4251 gnd.n2918 gnd.n2916 585
R4252 gnd.n3604 gnd.n2916 585
R4253 gnd.n5958 gnd.n5957 585
R4254 gnd.n5959 gnd.n5958 585
R4255 gnd.n2917 gnd.n2915 585
R4256 gnd.n4495 gnd.n2915 585
R4257 gnd.n3685 gnd.n3683 585
R4258 gnd.n3683 gnd.n2885 585
R4259 gnd.n4482 gnd.n4481 585
R4260 gnd.n4483 gnd.n4482 585
R4261 gnd.n3684 gnd.n3682 585
R4262 gnd.n3691 gnd.n3682 585
R4263 gnd.n4476 gnd.n4475 585
R4264 gnd.n4475 gnd.n4474 585
R4265 gnd.n3688 gnd.n3687 585
R4266 gnd.n4452 gnd.n3688 585
R4267 gnd.n3710 gnd.n3708 585
R4268 gnd.n3708 gnd.n3698 585
R4269 gnd.n4442 gnd.n4441 585
R4270 gnd.n4443 gnd.n4442 585
R4271 gnd.n3709 gnd.n3707 585
R4272 gnd.n3716 gnd.n3707 585
R4273 gnd.n4436 gnd.n4435 585
R4274 gnd.n4435 gnd.n4434 585
R4275 gnd.n3713 gnd.n3712 585
R4276 gnd.n4422 gnd.n3713 585
R4277 gnd.n3735 gnd.n3733 585
R4278 gnd.n3733 gnd.n3732 585
R4279 gnd.n4412 gnd.n4411 585
R4280 gnd.n4413 gnd.n4412 585
R4281 gnd.n3734 gnd.n3731 585
R4282 gnd.n3741 gnd.n3731 585
R4283 gnd.n4406 gnd.n4405 585
R4284 gnd.n4405 gnd.n4404 585
R4285 gnd.n3738 gnd.n3737 585
R4286 gnd.n4392 gnd.n3738 585
R4287 gnd.n4380 gnd.n4379 585
R4288 gnd.n4381 gnd.n4380 585
R4289 gnd.n4376 gnd.n2604 585
R4290 gnd.n4374 gnd.n2604 585
R4291 gnd.n6147 gnd.n6146 585
R4292 gnd.n6145 gnd.n2603 585
R4293 gnd.n2606 gnd.n2602 585
R4294 gnd.n6149 gnd.n2602 585
R4295 gnd.n6141 gnd.n2608 585
R4296 gnd.n6140 gnd.n2609 585
R4297 gnd.n6139 gnd.n2610 585
R4298 gnd.n2613 gnd.n2611 585
R4299 gnd.n6134 gnd.n2614 585
R4300 gnd.n6133 gnd.n2615 585
R4301 gnd.n6132 gnd.n2616 585
R4302 gnd.n2625 gnd.n2617 585
R4303 gnd.n6125 gnd.n2626 585
R4304 gnd.n6124 gnd.n2627 585
R4305 gnd.n2629 gnd.n2628 585
R4306 gnd.n6117 gnd.n2635 585
R4307 gnd.n6116 gnd.n2636 585
R4308 gnd.n2643 gnd.n2637 585
R4309 gnd.n6109 gnd.n2644 585
R4310 gnd.n6108 gnd.n2645 585
R4311 gnd.n2647 gnd.n2646 585
R4312 gnd.n6101 gnd.n2653 585
R4313 gnd.n6100 gnd.n2654 585
R4314 gnd.n2661 gnd.n2655 585
R4315 gnd.n6093 gnd.n2662 585
R4316 gnd.n6092 gnd.n2663 585
R4317 gnd.n2668 gnd.n2667 585
R4318 gnd.n2599 gnd.n2584 585
R4319 gnd.n6153 gnd.n2585 585
R4320 gnd.n6152 gnd.n6151 585
R4321 gnd.n3360 gnd.n3001 585
R4322 gnd.n5859 gnd.n3001 585
R4323 gnd.n5173 gnd.n5172 585
R4324 gnd.n5174 gnd.n5173 585
R4325 gnd.n3359 gnd.n3358 585
R4326 gnd.n5181 gnd.n3358 585
R4327 gnd.n4989 gnd.n3357 585
R4328 gnd.n5184 gnd.n3357 585
R4329 gnd.n4988 gnd.n4987 585
R4330 gnd.n4987 gnd.n3356 585
R4331 gnd.n4986 gnd.n4985 585
R4332 gnd.n4986 gnd.n3347 585
R4333 gnd.n3362 gnd.n3346 585
R4334 gnd.n5192 gnd.n3346 585
R4335 gnd.n4981 gnd.n3345 585
R4336 gnd.n5195 gnd.n3345 585
R4337 gnd.n4980 gnd.n4979 585
R4338 gnd.n4979 gnd.n3344 585
R4339 gnd.n4978 gnd.n4977 585
R4340 gnd.n4978 gnd.n3335 585
R4341 gnd.n3364 gnd.n3334 585
R4342 gnd.n5203 gnd.n3334 585
R4343 gnd.n4973 gnd.n3333 585
R4344 gnd.n5206 gnd.n3333 585
R4345 gnd.n4972 gnd.n4971 585
R4346 gnd.n4971 gnd.n3332 585
R4347 gnd.n4970 gnd.n4969 585
R4348 gnd.n4970 gnd.n3323 585
R4349 gnd.n3366 gnd.n3322 585
R4350 gnd.n5214 gnd.n3322 585
R4351 gnd.n4965 gnd.n3321 585
R4352 gnd.n5217 gnd.n3321 585
R4353 gnd.n4964 gnd.n4963 585
R4354 gnd.n4963 gnd.n3267 585
R4355 gnd.n4962 gnd.n4961 585
R4356 gnd.n4962 gnd.n3304 585
R4357 gnd.n3368 gnd.n3312 585
R4358 gnd.n5226 gnd.n3312 585
R4359 gnd.n4957 gnd.n4956 585
R4360 gnd.n4956 gnd.n4955 585
R4361 gnd.n3371 gnd.n3370 585
R4362 gnd.n3378 gnd.n3371 585
R4363 gnd.n4906 gnd.n4905 585
R4364 gnd.n4905 gnd.n3386 585
R4365 gnd.n4907 gnd.n4904 585
R4366 gnd.n4904 gnd.n3383 585
R4367 gnd.n3403 gnd.n3394 585
R4368 gnd.n4922 gnd.n3394 585
R4369 gnd.n4912 gnd.n4911 585
R4370 gnd.n4913 gnd.n4912 585
R4371 gnd.n3402 gnd.n3401 585
R4372 gnd.n4828 gnd.n3401 585
R4373 gnd.n4900 gnd.n4899 585
R4374 gnd.n4899 gnd.n4898 585
R4375 gnd.n3406 gnd.n3405 585
R4376 gnd.n4890 gnd.n3406 585
R4377 gnd.n3432 gnd.n3430 585
R4378 gnd.n3430 gnd.n3422 585
R4379 gnd.n4867 gnd.n4866 585
R4380 gnd.n4868 gnd.n4867 585
R4381 gnd.n3431 gnd.n3429 585
R4382 gnd.n3429 gnd.n3426 585
R4383 gnd.n4861 gnd.n4860 585
R4384 gnd.n4860 gnd.n4859 585
R4385 gnd.n3435 gnd.n3434 585
R4386 gnd.n3444 gnd.n3435 585
R4387 gnd.n4741 gnd.n4739 585
R4388 gnd.n4739 gnd.n4738 585
R4389 gnd.n4742 gnd.n4736 585
R4390 gnd.n4736 gnd.n3449 585
R4391 gnd.n4743 gnd.n3457 585
R4392 gnd.n4800 gnd.n3457 585
R4393 gnd.n4734 gnd.n3464 585
R4394 gnd.n4788 gnd.n3464 585
R4395 gnd.n4747 gnd.n4733 585
R4396 gnd.n4733 gnd.n3469 585
R4397 gnd.n4748 gnd.n4732 585
R4398 gnd.n4732 gnd.n3476 585
R4399 gnd.n4749 gnd.n4731 585
R4400 gnd.n4731 gnd.n4730 585
R4401 gnd.n3493 gnd.n3483 585
R4402 gnd.n4763 gnd.n3483 585
R4403 gnd.n4754 gnd.n4753 585
R4404 gnd.n4755 gnd.n4754 585
R4405 gnd.n3492 gnd.n3491 585
R4406 gnd.n4717 gnd.n3491 585
R4407 gnd.n4691 gnd.n4690 585
R4408 gnd.n4690 gnd.n4689 585
R4409 gnd.n3516 gnd.n3514 585
R4410 gnd.n3514 gnd.n3506 585
R4411 gnd.n4696 gnd.n4695 585
R4412 gnd.n4697 gnd.n4696 585
R4413 gnd.n3515 gnd.n3513 585
R4414 gnd.n4677 gnd.n3513 585
R4415 gnd.n4648 gnd.n4647 585
R4416 gnd.n4650 gnd.n4648 585
R4417 gnd.n3540 gnd.n3539 585
R4418 gnd.n3539 gnd.n3529 585
R4419 gnd.n4643 gnd.n4642 585
R4420 gnd.n4642 gnd.n4641 585
R4421 gnd.n4640 gnd.n3542 585
R4422 gnd.n4640 gnd.n3534 585
R4423 gnd.n4639 gnd.n3544 585
R4424 gnd.n4639 gnd.n4638 585
R4425 gnd.n4554 gnd.n3543 585
R4426 gnd.n4629 gnd.n3543 585
R4427 gnd.n4555 gnd.n3561 585
R4428 gnd.n4616 gnd.n3561 585
R4429 gnd.n4551 gnd.n4550 585
R4430 gnd.n4550 gnd.n3566 585
R4431 gnd.n4559 gnd.n4549 585
R4432 gnd.n4549 gnd.n4548 585
R4433 gnd.n4560 gnd.n4545 585
R4434 gnd.n4545 gnd.n3571 585
R4435 gnd.n4561 gnd.n3578 585
R4436 gnd.n4589 gnd.n3578 585
R4437 gnd.n3592 gnd.n3586 585
R4438 gnd.n4581 gnd.n3586 585
R4439 gnd.n4566 gnd.n4565 585
R4440 gnd.n4568 gnd.n4566 585
R4441 gnd.n3591 gnd.n3590 585
R4442 gnd.n4518 gnd.n3590 585
R4443 gnd.n4541 gnd.n4540 585
R4444 gnd.n4540 gnd.n4539 585
R4445 gnd.n3595 gnd.n3594 585
R4446 gnd.n3606 gnd.n3595 585
R4447 gnd.n4489 gnd.n4488 585
R4448 gnd.n4488 gnd.n3604 585
R4449 gnd.n3676 gnd.n2913 585
R4450 gnd.n5959 gnd.n2913 585
R4451 gnd.n4494 gnd.n4493 585
R4452 gnd.n4495 gnd.n4494 585
R4453 gnd.n3675 gnd.n3674 585
R4454 gnd.n3674 gnd.n2885 585
R4455 gnd.n4485 gnd.n4484 585
R4456 gnd.n4484 gnd.n4483 585
R4457 gnd.n3679 gnd.n3678 585
R4458 gnd.n3691 gnd.n3679 585
R4459 gnd.n3701 gnd.n3690 585
R4460 gnd.n4474 gnd.n3690 585
R4461 gnd.n4451 gnd.n4450 585
R4462 gnd.n4452 gnd.n4451 585
R4463 gnd.n3700 gnd.n3699 585
R4464 gnd.n3699 gnd.n3698 585
R4465 gnd.n4445 gnd.n4444 585
R4466 gnd.n4444 gnd.n4443 585
R4467 gnd.n3704 gnd.n3703 585
R4468 gnd.n3716 gnd.n3704 585
R4469 gnd.n3725 gnd.n3715 585
R4470 gnd.n4434 gnd.n3715 585
R4471 gnd.n4421 gnd.n4420 585
R4472 gnd.n4422 gnd.n4421 585
R4473 gnd.n3724 gnd.n3723 585
R4474 gnd.n3732 gnd.n3723 585
R4475 gnd.n4415 gnd.n4414 585
R4476 gnd.n4414 gnd.n4413 585
R4477 gnd.n3728 gnd.n3727 585
R4478 gnd.n3741 gnd.n3728 585
R4479 gnd.n4384 gnd.n3740 585
R4480 gnd.n4404 gnd.n3740 585
R4481 gnd.n4391 gnd.n4390 585
R4482 gnd.n4392 gnd.n4391 585
R4483 gnd.n4383 gnd.n4382 585
R4484 gnd.n4382 gnd.n4381 585
R4485 gnd.n4385 gnd.n2586 585
R4486 gnd.n4374 gnd.n2586 585
R4487 gnd.n5147 gnd.n5001 585
R4488 gnd.n5001 gnd.n3011 585
R4489 gnd.n5148 gnd.n5145 585
R4490 gnd.n5143 gnd.n5019 585
R4491 gnd.n5142 gnd.n5141 585
R4492 gnd.n5126 gnd.n5021 585
R4493 gnd.n5128 gnd.n5127 585
R4494 gnd.n5124 gnd.n5028 585
R4495 gnd.n5123 gnd.n5122 585
R4496 gnd.n5107 gnd.n5030 585
R4497 gnd.n5109 gnd.n5108 585
R4498 gnd.n5105 gnd.n5037 585
R4499 gnd.n5104 gnd.n5103 585
R4500 gnd.n5088 gnd.n5039 585
R4501 gnd.n5090 gnd.n5089 585
R4502 gnd.n5086 gnd.n5046 585
R4503 gnd.n5085 gnd.n5084 585
R4504 gnd.n5073 gnd.n5048 585
R4505 gnd.n5075 gnd.n5074 585
R4506 gnd.n5071 gnd.n5049 585
R4507 gnd.n5070 gnd.n5069 585
R4508 gnd.n5062 gnd.n5051 585
R4509 gnd.n5064 gnd.n5063 585
R4510 gnd.n5060 gnd.n5053 585
R4511 gnd.n5059 gnd.n5058 585
R4512 gnd.n5055 gnd.n2999 585
R4513 gnd.n5168 gnd.n5167 585
R4514 gnd.n5165 gnd.n4999 585
R4515 gnd.n5164 gnd.n5000 585
R4516 gnd.n5162 gnd.n5161 585
R4517 gnd.n6500 gnd.n705 540.215
R4518 gnd.n5316 gnd.n3307 463.671
R4519 gnd.n5319 gnd.n5318 463.671
R4520 gnd.n4497 gnd.n3673 463.671
R4521 gnd.n6028 gnd.n2888 463.671
R4522 gnd.n3609 gnd.t206 443.966
R4523 gnd.n3300 gnd.t227 443.966
R4524 gnd.n5965 gnd.t257 443.966
R4525 gnd.n5250 gnd.t279 443.966
R4526 gnd.n2664 gnd.t237 371.625
R4527 gnd.n5012 gnd.t263 371.625
R4528 gnd.n2671 gnd.t285 371.625
R4529 gnd.n5456 gnd.t260 371.625
R4530 gnd.n5508 gnd.t248 371.625
R4531 gnd.n3231 gnd.t193 371.625
R4532 gnd.n7348 gnd.t174 371.625
R4533 gnd.n7327 gnd.t190 371.625
R4534 gnd.n7434 gnd.t254 371.625
R4535 gnd.n180 gnd.t276 371.625
R4536 gnd.n3955 gnd.t221 371.625
R4537 gnd.n4066 gnd.t203 371.625
R4538 gnd.n3911 gnd.t231 371.625
R4539 gnd.n3871 gnd.t186 371.625
R4540 gnd.n2741 gnd.t269 371.625
R4541 gnd.n2782 gnd.t210 371.625
R4542 gnd.n2761 gnd.t234 371.625
R4543 gnd.n5002 gnd.t217 371.625
R4544 gnd.n7232 gnd.n268 368.44
R4545 gnd.n1356 gnd.t244 323.425
R4546 gnd.n916 gnd.t272 323.425
R4547 gnd.n7022 gnd.n7021 301.784
R4548 gnd.n7023 gnd.n7022 301.784
R4549 gnd.n7023 gnd.n388 301.784
R4550 gnd.n7031 gnd.n388 301.784
R4551 gnd.n7032 gnd.n7031 301.784
R4552 gnd.n7033 gnd.n7032 301.784
R4553 gnd.n7033 gnd.n382 301.784
R4554 gnd.n7041 gnd.n382 301.784
R4555 gnd.n7042 gnd.n7041 301.784
R4556 gnd.n7043 gnd.n7042 301.784
R4557 gnd.n7043 gnd.n376 301.784
R4558 gnd.n7051 gnd.n376 301.784
R4559 gnd.n7052 gnd.n7051 301.784
R4560 gnd.n7053 gnd.n7052 301.784
R4561 gnd.n7053 gnd.n370 301.784
R4562 gnd.n7061 gnd.n370 301.784
R4563 gnd.n7062 gnd.n7061 301.784
R4564 gnd.n7063 gnd.n7062 301.784
R4565 gnd.n7063 gnd.n364 301.784
R4566 gnd.n7071 gnd.n364 301.784
R4567 gnd.n7072 gnd.n7071 301.784
R4568 gnd.n7073 gnd.n7072 301.784
R4569 gnd.n7073 gnd.n358 301.784
R4570 gnd.n7081 gnd.n358 301.784
R4571 gnd.n7082 gnd.n7081 301.784
R4572 gnd.n7083 gnd.n7082 301.784
R4573 gnd.n7083 gnd.n352 301.784
R4574 gnd.n7091 gnd.n352 301.784
R4575 gnd.n7092 gnd.n7091 301.784
R4576 gnd.n7093 gnd.n7092 301.784
R4577 gnd.n7093 gnd.n346 301.784
R4578 gnd.n7101 gnd.n346 301.784
R4579 gnd.n7102 gnd.n7101 301.784
R4580 gnd.n7103 gnd.n7102 301.784
R4581 gnd.n7103 gnd.n340 301.784
R4582 gnd.n7111 gnd.n340 301.784
R4583 gnd.n7112 gnd.n7111 301.784
R4584 gnd.n7113 gnd.n7112 301.784
R4585 gnd.n7113 gnd.n334 301.784
R4586 gnd.n7121 gnd.n334 301.784
R4587 gnd.n7122 gnd.n7121 301.784
R4588 gnd.n7123 gnd.n7122 301.784
R4589 gnd.n7123 gnd.n328 301.784
R4590 gnd.n7131 gnd.n328 301.784
R4591 gnd.n7132 gnd.n7131 301.784
R4592 gnd.n7133 gnd.n7132 301.784
R4593 gnd.n7133 gnd.n322 301.784
R4594 gnd.n7141 gnd.n322 301.784
R4595 gnd.n7142 gnd.n7141 301.784
R4596 gnd.n7143 gnd.n7142 301.784
R4597 gnd.n7143 gnd.n316 301.784
R4598 gnd.n7151 gnd.n316 301.784
R4599 gnd.n7152 gnd.n7151 301.784
R4600 gnd.n7153 gnd.n7152 301.784
R4601 gnd.n7153 gnd.n310 301.784
R4602 gnd.n7161 gnd.n310 301.784
R4603 gnd.n7162 gnd.n7161 301.784
R4604 gnd.n7163 gnd.n7162 301.784
R4605 gnd.n7163 gnd.n304 301.784
R4606 gnd.n7171 gnd.n304 301.784
R4607 gnd.n7172 gnd.n7171 301.784
R4608 gnd.n7173 gnd.n7172 301.784
R4609 gnd.n7173 gnd.n298 301.784
R4610 gnd.n7181 gnd.n298 301.784
R4611 gnd.n7182 gnd.n7181 301.784
R4612 gnd.n7183 gnd.n7182 301.784
R4613 gnd.n7183 gnd.n292 301.784
R4614 gnd.n7191 gnd.n292 301.784
R4615 gnd.n7192 gnd.n7191 301.784
R4616 gnd.n7193 gnd.n7192 301.784
R4617 gnd.n7193 gnd.n286 301.784
R4618 gnd.n7201 gnd.n286 301.784
R4619 gnd.n7202 gnd.n7201 301.784
R4620 gnd.n7203 gnd.n7202 301.784
R4621 gnd.n7203 gnd.n280 301.784
R4622 gnd.n7211 gnd.n280 301.784
R4623 gnd.n7212 gnd.n7211 301.784
R4624 gnd.n7213 gnd.n7212 301.784
R4625 gnd.n7213 gnd.n274 301.784
R4626 gnd.n7221 gnd.n274 301.784
R4627 gnd.n7222 gnd.n7221 301.784
R4628 gnd.n7223 gnd.n7222 301.784
R4629 gnd.n7223 gnd.n268 301.784
R4630 gnd.n2206 gnd.n2180 289.615
R4631 gnd.n2174 gnd.n2148 289.615
R4632 gnd.n2142 gnd.n2116 289.615
R4633 gnd.n2111 gnd.n2085 289.615
R4634 gnd.n2079 gnd.n2053 289.615
R4635 gnd.n2047 gnd.n2021 289.615
R4636 gnd.n2015 gnd.n1989 289.615
R4637 gnd.n1984 gnd.n1958 289.615
R4638 gnd.n1430 gnd.t182 279.217
R4639 gnd.n942 gnd.t178 279.217
R4640 gnd.n2895 gnd.t216 260.649
R4641 gnd.n5242 gnd.t202 260.649
R4642 gnd.n6030 gnd.n6029 256.663
R4643 gnd.n6030 gnd.n2854 256.663
R4644 gnd.n6030 gnd.n2855 256.663
R4645 gnd.n6030 gnd.n2856 256.663
R4646 gnd.n6030 gnd.n2857 256.663
R4647 gnd.n6030 gnd.n2858 256.663
R4648 gnd.n6030 gnd.n2859 256.663
R4649 gnd.n6030 gnd.n2860 256.663
R4650 gnd.n6030 gnd.n2861 256.663
R4651 gnd.n6030 gnd.n2862 256.663
R4652 gnd.n6030 gnd.n2863 256.663
R4653 gnd.n6030 gnd.n2864 256.663
R4654 gnd.n6030 gnd.n2865 256.663
R4655 gnd.n6030 gnd.n2866 256.663
R4656 gnd.n6030 gnd.n2867 256.663
R4657 gnd.n6030 gnd.n2868 256.663
R4658 gnd.n6033 gnd.n2852 256.663
R4659 gnd.n6031 gnd.n6030 256.663
R4660 gnd.n6030 gnd.n2869 256.663
R4661 gnd.n6030 gnd.n2870 256.663
R4662 gnd.n6030 gnd.n2871 256.663
R4663 gnd.n6030 gnd.n2872 256.663
R4664 gnd.n6030 gnd.n2873 256.663
R4665 gnd.n6030 gnd.n2874 256.663
R4666 gnd.n6030 gnd.n2875 256.663
R4667 gnd.n6030 gnd.n2876 256.663
R4668 gnd.n6030 gnd.n2877 256.663
R4669 gnd.n6030 gnd.n2878 256.663
R4670 gnd.n6030 gnd.n2879 256.663
R4671 gnd.n6030 gnd.n2880 256.663
R4672 gnd.n6030 gnd.n2881 256.663
R4673 gnd.n6030 gnd.n2882 256.663
R4674 gnd.n6030 gnd.n2883 256.663
R4675 gnd.n6030 gnd.n2884 256.663
R4676 gnd.n5384 gnd.n3284 256.663
R4677 gnd.n5384 gnd.n3285 256.663
R4678 gnd.n5384 gnd.n3286 256.663
R4679 gnd.n5384 gnd.n3287 256.663
R4680 gnd.n5384 gnd.n3288 256.663
R4681 gnd.n5384 gnd.n3289 256.663
R4682 gnd.n5384 gnd.n3290 256.663
R4683 gnd.n5384 gnd.n3291 256.663
R4684 gnd.n5384 gnd.n3292 256.663
R4685 gnd.n5384 gnd.n3293 256.663
R4686 gnd.n5384 gnd.n3294 256.663
R4687 gnd.n5384 gnd.n3295 256.663
R4688 gnd.n5384 gnd.n3296 256.663
R4689 gnd.n5384 gnd.n3297 256.663
R4690 gnd.n5384 gnd.n3298 256.663
R4691 gnd.n5384 gnd.n5381 256.663
R4692 gnd.n5387 gnd.n3265 256.663
R4693 gnd.n5385 gnd.n5384 256.663
R4694 gnd.n5384 gnd.n3283 256.663
R4695 gnd.n5384 gnd.n3282 256.663
R4696 gnd.n5384 gnd.n3281 256.663
R4697 gnd.n5384 gnd.n3280 256.663
R4698 gnd.n5384 gnd.n3279 256.663
R4699 gnd.n5384 gnd.n3278 256.663
R4700 gnd.n5384 gnd.n3277 256.663
R4701 gnd.n5384 gnd.n3276 256.663
R4702 gnd.n5384 gnd.n3275 256.663
R4703 gnd.n5384 gnd.n3274 256.663
R4704 gnd.n5384 gnd.n3273 256.663
R4705 gnd.n5384 gnd.n3272 256.663
R4706 gnd.n5384 gnd.n3271 256.663
R4707 gnd.n5384 gnd.n3270 256.663
R4708 gnd.n5384 gnd.n3269 256.663
R4709 gnd.n5384 gnd.n3268 256.663
R4710 gnd.n3906 gnd.n2363 242.672
R4711 gnd.n3843 gnd.n2363 242.672
R4712 gnd.n3899 gnd.n2363 242.672
R4713 gnd.n3893 gnd.n2363 242.672
R4714 gnd.n3891 gnd.n2363 242.672
R4715 gnd.n3885 gnd.n2363 242.672
R4716 gnd.n3883 gnd.n2363 242.672
R4717 gnd.n3877 gnd.n2363 242.672
R4718 gnd.n3875 gnd.n2363 242.672
R4719 gnd.n6085 gnd.n6084 242.672
R4720 gnd.n6084 gnd.n2689 242.672
R4721 gnd.n6084 gnd.n2687 242.672
R4722 gnd.n6084 gnd.n2686 242.672
R4723 gnd.n6084 gnd.n2684 242.672
R4724 gnd.n6084 gnd.n2682 242.672
R4725 gnd.n6084 gnd.n2681 242.672
R4726 gnd.n6084 gnd.n2679 242.672
R4727 gnd.n6084 gnd.n2677 242.672
R4728 gnd.n1484 gnd.n1483 242.672
R4729 gnd.n1484 gnd.n1394 242.672
R4730 gnd.n1484 gnd.n1395 242.672
R4731 gnd.n1484 gnd.n1396 242.672
R4732 gnd.n1484 gnd.n1397 242.672
R4733 gnd.n1484 gnd.n1398 242.672
R4734 gnd.n1484 gnd.n1399 242.672
R4735 gnd.n1484 gnd.n1400 242.672
R4736 gnd.n1484 gnd.n1401 242.672
R4737 gnd.n1484 gnd.n1402 242.672
R4738 gnd.n1484 gnd.n1403 242.672
R4739 gnd.n1484 gnd.n1404 242.672
R4740 gnd.n1485 gnd.n1484 242.672
R4741 gnd.n2338 gnd.n891 242.672
R4742 gnd.n2338 gnd.n890 242.672
R4743 gnd.n2338 gnd.n889 242.672
R4744 gnd.n2338 gnd.n888 242.672
R4745 gnd.n2338 gnd.n887 242.672
R4746 gnd.n2338 gnd.n886 242.672
R4747 gnd.n2338 gnd.n885 242.672
R4748 gnd.n2338 gnd.n884 242.672
R4749 gnd.n2338 gnd.n883 242.672
R4750 gnd.n2338 gnd.n882 242.672
R4751 gnd.n2338 gnd.n881 242.672
R4752 gnd.n2338 gnd.n880 242.672
R4753 gnd.n2338 gnd.n879 242.672
R4754 gnd.n5078 gnd.n3012 242.672
R4755 gnd.n5095 gnd.n3012 242.672
R4756 gnd.n5097 gnd.n3012 242.672
R4757 gnd.n5114 gnd.n3012 242.672
R4758 gnd.n5116 gnd.n3012 242.672
R4759 gnd.n5133 gnd.n3012 242.672
R4760 gnd.n5135 gnd.n3012 242.672
R4761 gnd.n5153 gnd.n3012 242.672
R4762 gnd.n5155 gnd.n3012 242.672
R4763 gnd.n7470 gnd.n7469 242.672
R4764 gnd.n7469 gnd.n242 242.672
R4765 gnd.n7469 gnd.n191 242.672
R4766 gnd.n7469 gnd.n190 242.672
R4767 gnd.n7469 gnd.n189 242.672
R4768 gnd.n7469 gnd.n188 242.672
R4769 gnd.n7469 gnd.n187 242.672
R4770 gnd.n7469 gnd.n186 242.672
R4771 gnd.n7469 gnd.n185 242.672
R4772 gnd.n1568 gnd.n1567 242.672
R4773 gnd.n1567 gnd.n1306 242.672
R4774 gnd.n1567 gnd.n1307 242.672
R4775 gnd.n1567 gnd.n1308 242.672
R4776 gnd.n1567 gnd.n1309 242.672
R4777 gnd.n1567 gnd.n1310 242.672
R4778 gnd.n1567 gnd.n1311 242.672
R4779 gnd.n1567 gnd.n1312 242.672
R4780 gnd.n2338 gnd.n892 242.672
R4781 gnd.n2338 gnd.n893 242.672
R4782 gnd.n2338 gnd.n894 242.672
R4783 gnd.n2338 gnd.n895 242.672
R4784 gnd.n2338 gnd.n896 242.672
R4785 gnd.n2338 gnd.n897 242.672
R4786 gnd.n2338 gnd.n898 242.672
R4787 gnd.n2338 gnd.n899 242.672
R4788 gnd.n3974 gnd.n2363 242.672
R4789 gnd.n3982 gnd.n2363 242.672
R4790 gnd.n3984 gnd.n2363 242.672
R4791 gnd.n3992 gnd.n2363 242.672
R4792 gnd.n3994 gnd.n2363 242.672
R4793 gnd.n4002 gnd.n2363 242.672
R4794 gnd.n4004 gnd.n2363 242.672
R4795 gnd.n4012 gnd.n2363 242.672
R4796 gnd.n4014 gnd.n2363 242.672
R4797 gnd.n4022 gnd.n2363 242.672
R4798 gnd.n4024 gnd.n2363 242.672
R4799 gnd.n4032 gnd.n2363 242.672
R4800 gnd.n4034 gnd.n2363 242.672
R4801 gnd.n4042 gnd.n2363 242.672
R4802 gnd.n4044 gnd.n2363 242.672
R4803 gnd.n4052 gnd.n2363 242.672
R4804 gnd.n4054 gnd.n2363 242.672
R4805 gnd.n4062 gnd.n2363 242.672
R4806 gnd.n4064 gnd.n2363 242.672
R4807 gnd.n4074 gnd.n2363 242.672
R4808 gnd.n4076 gnd.n2363 242.672
R4809 gnd.n4084 gnd.n2363 242.672
R4810 gnd.n4086 gnd.n2363 242.672
R4811 gnd.n4094 gnd.n2363 242.672
R4812 gnd.n4096 gnd.n2363 242.672
R4813 gnd.n4104 gnd.n2363 242.672
R4814 gnd.n4106 gnd.n2363 242.672
R4815 gnd.n4115 gnd.n2363 242.672
R4816 gnd.n4118 gnd.n2363 242.672
R4817 gnd.n6084 gnd.n2691 242.672
R4818 gnd.n6084 gnd.n2692 242.672
R4819 gnd.n6084 gnd.n2693 242.672
R4820 gnd.n6084 gnd.n2694 242.672
R4821 gnd.n6084 gnd.n2695 242.672
R4822 gnd.n6084 gnd.n2696 242.672
R4823 gnd.n6084 gnd.n2697 242.672
R4824 gnd.n6084 gnd.n2698 242.672
R4825 gnd.n6084 gnd.n2699 242.672
R4826 gnd.n6084 gnd.n2700 242.672
R4827 gnd.n6084 gnd.n2701 242.672
R4828 gnd.n6084 gnd.n2702 242.672
R4829 gnd.n6084 gnd.n2703 242.672
R4830 gnd.n6084 gnd.n2704 242.672
R4831 gnd.n6084 gnd.n2705 242.672
R4832 gnd.n6084 gnd.n2706 242.672
R4833 gnd.n6034 gnd.n2752 242.672
R4834 gnd.n6084 gnd.n2707 242.672
R4835 gnd.n6084 gnd.n2708 242.672
R4836 gnd.n6084 gnd.n2709 242.672
R4837 gnd.n6084 gnd.n2710 242.672
R4838 gnd.n6084 gnd.n2711 242.672
R4839 gnd.n6084 gnd.n2712 242.672
R4840 gnd.n6084 gnd.n2713 242.672
R4841 gnd.n6084 gnd.n2714 242.672
R4842 gnd.n6084 gnd.n2715 242.672
R4843 gnd.n6084 gnd.n2716 242.672
R4844 gnd.n6084 gnd.n2717 242.672
R4845 gnd.n6084 gnd.n2718 242.672
R4846 gnd.n6084 gnd.n6083 242.672
R4847 gnd.n5417 gnd.n3012 242.672
R4848 gnd.n5420 gnd.n3012 242.672
R4849 gnd.n5428 gnd.n3012 242.672
R4850 gnd.n5430 gnd.n3012 242.672
R4851 gnd.n5438 gnd.n3012 242.672
R4852 gnd.n5440 gnd.n3012 242.672
R4853 gnd.n5448 gnd.n3012 242.672
R4854 gnd.n5450 gnd.n3012 242.672
R4855 gnd.n5461 gnd.n3012 242.672
R4856 gnd.n5463 gnd.n3012 242.672
R4857 gnd.n5471 gnd.n3012 242.672
R4858 gnd.n5473 gnd.n3012 242.672
R4859 gnd.n5482 gnd.n3012 242.672
R4860 gnd.n5483 gnd.n5388 242.672
R4861 gnd.n5484 gnd.n3012 242.672
R4862 gnd.n5486 gnd.n3012 242.672
R4863 gnd.n5494 gnd.n3012 242.672
R4864 gnd.n5496 gnd.n3012 242.672
R4865 gnd.n5504 gnd.n3012 242.672
R4866 gnd.n5506 gnd.n3012 242.672
R4867 gnd.n5516 gnd.n3012 242.672
R4868 gnd.n5518 gnd.n3012 242.672
R4869 gnd.n5526 gnd.n3012 242.672
R4870 gnd.n5528 gnd.n3012 242.672
R4871 gnd.n5536 gnd.n3012 242.672
R4872 gnd.n5538 gnd.n3012 242.672
R4873 gnd.n5546 gnd.n3012 242.672
R4874 gnd.n5548 gnd.n3012 242.672
R4875 gnd.n5557 gnd.n3012 242.672
R4876 gnd.n5560 gnd.n3012 242.672
R4877 gnd.n7469 gnd.n7257 242.672
R4878 gnd.n7469 gnd.n7258 242.672
R4879 gnd.n7469 gnd.n7259 242.672
R4880 gnd.n7469 gnd.n7260 242.672
R4881 gnd.n7469 gnd.n7261 242.672
R4882 gnd.n7469 gnd.n7262 242.672
R4883 gnd.n7469 gnd.n7263 242.672
R4884 gnd.n7469 gnd.n7264 242.672
R4885 gnd.n7469 gnd.n7265 242.672
R4886 gnd.n7469 gnd.n7266 242.672
R4887 gnd.n7469 gnd.n7267 242.672
R4888 gnd.n7469 gnd.n7268 242.672
R4889 gnd.n7469 gnd.n7269 242.672
R4890 gnd.n7469 gnd.n7270 242.672
R4891 gnd.n7469 gnd.n7271 242.672
R4892 gnd.n7469 gnd.n7272 242.672
R4893 gnd.n7469 gnd.n7273 242.672
R4894 gnd.n7469 gnd.n7274 242.672
R4895 gnd.n7469 gnd.n7275 242.672
R4896 gnd.n7469 gnd.n7276 242.672
R4897 gnd.n7469 gnd.n7277 242.672
R4898 gnd.n7469 gnd.n7278 242.672
R4899 gnd.n7469 gnd.n7279 242.672
R4900 gnd.n7469 gnd.n7280 242.672
R4901 gnd.n7469 gnd.n7281 242.672
R4902 gnd.n7469 gnd.n7282 242.672
R4903 gnd.n7469 gnd.n7283 242.672
R4904 gnd.n7469 gnd.n7284 242.672
R4905 gnd.n7469 gnd.n7468 242.672
R4906 gnd.n6149 gnd.n6148 242.672
R4907 gnd.n6149 gnd.n2588 242.672
R4908 gnd.n6149 gnd.n2589 242.672
R4909 gnd.n6149 gnd.n2590 242.672
R4910 gnd.n6149 gnd.n2591 242.672
R4911 gnd.n6149 gnd.n2592 242.672
R4912 gnd.n6149 gnd.n2593 242.672
R4913 gnd.n6149 gnd.n2594 242.672
R4914 gnd.n6149 gnd.n2595 242.672
R4915 gnd.n6149 gnd.n2596 242.672
R4916 gnd.n6149 gnd.n2597 242.672
R4917 gnd.n6149 gnd.n2598 242.672
R4918 gnd.n6149 gnd.n2600 242.672
R4919 gnd.n6150 gnd.n6149 242.672
R4920 gnd.n5144 gnd.n3011 242.672
R4921 gnd.n5020 gnd.n3011 242.672
R4922 gnd.n5125 gnd.n3011 242.672
R4923 gnd.n5029 gnd.n3011 242.672
R4924 gnd.n5106 gnd.n3011 242.672
R4925 gnd.n5038 gnd.n3011 242.672
R4926 gnd.n5087 gnd.n3011 242.672
R4927 gnd.n5047 gnd.n3011 242.672
R4928 gnd.n5072 gnd.n3011 242.672
R4929 gnd.n5050 gnd.n3011 242.672
R4930 gnd.n5061 gnd.n3011 242.672
R4931 gnd.n5054 gnd.n3011 242.672
R4932 gnd.n5166 gnd.n3011 242.672
R4933 gnd.n5163 gnd.n3011 242.672
R4934 gnd.n7285 gnd.n167 240.244
R4935 gnd.n7467 gnd.n7286 240.244
R4936 gnd.n7463 gnd.n7462 240.244
R4937 gnd.n7459 gnd.n7458 240.244
R4938 gnd.n7455 gnd.n7454 240.244
R4939 gnd.n7451 gnd.n7450 240.244
R4940 gnd.n7447 gnd.n7446 240.244
R4941 gnd.n7443 gnd.n7442 240.244
R4942 gnd.n7439 gnd.n7438 240.244
R4943 gnd.n7432 gnd.n7431 240.244
R4944 gnd.n7428 gnd.n7427 240.244
R4945 gnd.n7424 gnd.n7423 240.244
R4946 gnd.n7420 gnd.n7419 240.244
R4947 gnd.n7416 gnd.n7415 240.244
R4948 gnd.n7412 gnd.n7411 240.244
R4949 gnd.n7408 gnd.n7407 240.244
R4950 gnd.n7404 gnd.n7403 240.244
R4951 gnd.n7400 gnd.n7399 240.244
R4952 gnd.n7396 gnd.n7395 240.244
R4953 gnd.n7389 gnd.n7388 240.244
R4954 gnd.n7386 gnd.n7385 240.244
R4955 gnd.n7382 gnd.n7381 240.244
R4956 gnd.n7378 gnd.n7377 240.244
R4957 gnd.n7374 gnd.n7373 240.244
R4958 gnd.n7370 gnd.n7369 240.244
R4959 gnd.n7366 gnd.n7365 240.244
R4960 gnd.n7362 gnd.n7361 240.244
R4961 gnd.n7358 gnd.n7357 240.244
R4962 gnd.n7354 gnd.n7353 240.244
R4963 gnd.n3228 gnd.n3021 240.244
R4964 gnd.n3228 gnd.n3033 240.244
R4965 gnd.n5571 gnd.n3033 240.244
R4966 gnd.n5571 gnd.n3045 240.244
R4967 gnd.n5581 gnd.n3045 240.244
R4968 gnd.n5581 gnd.n3056 240.244
R4969 gnd.n3217 gnd.n3056 240.244
R4970 gnd.n3217 gnd.n3065 240.244
R4971 gnd.n5588 gnd.n3065 240.244
R4972 gnd.n5588 gnd.n3076 240.244
R4973 gnd.n5646 gnd.n3076 240.244
R4974 gnd.n5646 gnd.n3085 240.244
R4975 gnd.n5651 gnd.n3085 240.244
R4976 gnd.n5651 gnd.n3096 240.244
R4977 gnd.n5671 gnd.n3096 240.244
R4978 gnd.n5671 gnd.n3105 240.244
R4979 gnd.n3111 gnd.n3105 240.244
R4980 gnd.n5676 gnd.n3111 240.244
R4981 gnd.n5676 gnd.n5675 240.244
R4982 gnd.n5675 gnd.n3121 240.244
R4983 gnd.n3128 gnd.n3121 240.244
R4984 gnd.n5688 gnd.n3128 240.244
R4985 gnd.n5688 gnd.n70 240.244
R4986 gnd.n3137 gnd.n70 240.244
R4987 gnd.n5698 gnd.n3137 240.244
R4988 gnd.n5698 gnd.n87 240.244
R4989 gnd.n5702 gnd.n87 240.244
R4990 gnd.n5702 gnd.n99 240.244
R4991 gnd.n5713 gnd.n99 240.244
R4992 gnd.n5713 gnd.n109 240.244
R4993 gnd.n3191 gnd.n109 240.244
R4994 gnd.n3191 gnd.n118 240.244
R4995 gnd.n5748 gnd.n118 240.244
R4996 gnd.n5748 gnd.n129 240.244
R4997 gnd.n5744 gnd.n129 240.244
R4998 gnd.n5744 gnd.n139 240.244
R4999 gnd.n5736 gnd.n139 240.244
R5000 gnd.n5736 gnd.n150 240.244
R5001 gnd.n5732 gnd.n150 240.244
R5002 gnd.n5732 gnd.n160 240.244
R5003 gnd.n7479 gnd.n160 240.244
R5004 gnd.n7479 gnd.n169 240.244
R5005 gnd.n5419 gnd.n5418 240.244
R5006 gnd.n5421 gnd.n5419 240.244
R5007 gnd.n5427 gnd.n5409 240.244
R5008 gnd.n5431 gnd.n5429 240.244
R5009 gnd.n5437 gnd.n5405 240.244
R5010 gnd.n5441 gnd.n5439 240.244
R5011 gnd.n5447 gnd.n5401 240.244
R5012 gnd.n5451 gnd.n5449 240.244
R5013 gnd.n5460 gnd.n5397 240.244
R5014 gnd.n5464 gnd.n5462 240.244
R5015 gnd.n5470 gnd.n5393 240.244
R5016 gnd.n5474 gnd.n5472 240.244
R5017 gnd.n5481 gnd.n5389 240.244
R5018 gnd.n5487 gnd.n5485 240.244
R5019 gnd.n5493 gnd.n3259 240.244
R5020 gnd.n5497 gnd.n5495 240.244
R5021 gnd.n5503 gnd.n3255 240.244
R5022 gnd.n5507 gnd.n5505 240.244
R5023 gnd.n5515 gnd.n3251 240.244
R5024 gnd.n5519 gnd.n5517 240.244
R5025 gnd.n5525 gnd.n3247 240.244
R5026 gnd.n5529 gnd.n5527 240.244
R5027 gnd.n5535 gnd.n3243 240.244
R5028 gnd.n5539 gnd.n5537 240.244
R5029 gnd.n5545 gnd.n3239 240.244
R5030 gnd.n5549 gnd.n5547 240.244
R5031 gnd.n5556 gnd.n3235 240.244
R5032 gnd.n5559 gnd.n5558 240.244
R5033 gnd.n5842 gnd.n3026 240.244
R5034 gnd.n5838 gnd.n3026 240.244
R5035 gnd.n5838 gnd.n3031 240.244
R5036 gnd.n5830 gnd.n3031 240.244
R5037 gnd.n5830 gnd.n3048 240.244
R5038 gnd.n5826 gnd.n3048 240.244
R5039 gnd.n5826 gnd.n3054 240.244
R5040 gnd.n5818 gnd.n3054 240.244
R5041 gnd.n5818 gnd.n3068 240.244
R5042 gnd.n5814 gnd.n3068 240.244
R5043 gnd.n5814 gnd.n3074 240.244
R5044 gnd.n5806 gnd.n3074 240.244
R5045 gnd.n5806 gnd.n3088 240.244
R5046 gnd.n5802 gnd.n3088 240.244
R5047 gnd.n5802 gnd.n3094 240.244
R5048 gnd.n5794 gnd.n3094 240.244
R5049 gnd.n5794 gnd.n5792 240.244
R5050 gnd.n5792 gnd.n3108 240.244
R5051 gnd.n3125 gnd.n3108 240.244
R5052 gnd.n5781 gnd.n3125 240.244
R5053 gnd.n5781 gnd.n5778 240.244
R5054 gnd.n5778 gnd.n73 240.244
R5055 gnd.n7540 gnd.n73 240.244
R5056 gnd.n7540 gnd.n74 240.244
R5057 gnd.n84 gnd.n74 240.244
R5058 gnd.n7534 gnd.n84 240.244
R5059 gnd.n7534 gnd.n85 240.244
R5060 gnd.n7526 gnd.n85 240.244
R5061 gnd.n7526 gnd.n102 240.244
R5062 gnd.n7522 gnd.n102 240.244
R5063 gnd.n7522 gnd.n107 240.244
R5064 gnd.n7514 gnd.n107 240.244
R5065 gnd.n7514 gnd.n121 240.244
R5066 gnd.n7510 gnd.n121 240.244
R5067 gnd.n7510 gnd.n127 240.244
R5068 gnd.n7502 gnd.n127 240.244
R5069 gnd.n7502 gnd.n142 240.244
R5070 gnd.n7498 gnd.n142 240.244
R5071 gnd.n7498 gnd.n148 240.244
R5072 gnd.n7490 gnd.n148 240.244
R5073 gnd.n7490 gnd.n162 240.244
R5074 gnd.n7486 gnd.n162 240.244
R5075 gnd.n2719 gnd.n2570 240.244
R5076 gnd.n6082 gnd.n2720 240.244
R5077 gnd.n6078 gnd.n6077 240.244
R5078 gnd.n6074 gnd.n6073 240.244
R5079 gnd.n6070 gnd.n6069 240.244
R5080 gnd.n6066 gnd.n6065 240.244
R5081 gnd.n6062 gnd.n6061 240.244
R5082 gnd.n6058 gnd.n6057 240.244
R5083 gnd.n6054 gnd.n6053 240.244
R5084 gnd.n6049 gnd.n6048 240.244
R5085 gnd.n6045 gnd.n6044 240.244
R5086 gnd.n6041 gnd.n6040 240.244
R5087 gnd.n6037 gnd.n6036 240.244
R5088 gnd.n2845 gnd.n2844 240.244
R5089 gnd.n2842 gnd.n2841 240.244
R5090 gnd.n2838 gnd.n2837 240.244
R5091 gnd.n2834 gnd.n2833 240.244
R5092 gnd.n2830 gnd.n2829 240.244
R5093 gnd.n2823 gnd.n2822 240.244
R5094 gnd.n2820 gnd.n2819 240.244
R5095 gnd.n2816 gnd.n2815 240.244
R5096 gnd.n2812 gnd.n2811 240.244
R5097 gnd.n2808 gnd.n2807 240.244
R5098 gnd.n2804 gnd.n2803 240.244
R5099 gnd.n2800 gnd.n2799 240.244
R5100 gnd.n2796 gnd.n2795 240.244
R5101 gnd.n2792 gnd.n2791 240.244
R5102 gnd.n2788 gnd.n2787 240.244
R5103 gnd.n3834 gnd.n2364 240.244
R5104 gnd.n3834 gnd.n2375 240.244
R5105 gnd.n4159 gnd.n2375 240.244
R5106 gnd.n4159 gnd.n2387 240.244
R5107 gnd.n4155 gnd.n2387 240.244
R5108 gnd.n4155 gnd.n2398 240.244
R5109 gnd.n4147 gnd.n2398 240.244
R5110 gnd.n4147 gnd.n2408 240.244
R5111 gnd.n4143 gnd.n2408 240.244
R5112 gnd.n4143 gnd.n2419 240.244
R5113 gnd.n3818 gnd.n2419 240.244
R5114 gnd.n3818 gnd.n2428 240.244
R5115 gnd.n4206 gnd.n2428 240.244
R5116 gnd.n4206 gnd.n2439 240.244
R5117 gnd.n4210 gnd.n2439 240.244
R5118 gnd.n4210 gnd.n2449 240.244
R5119 gnd.n4221 gnd.n2449 240.244
R5120 gnd.n4221 gnd.n2458 240.244
R5121 gnd.n3800 gnd.n2458 240.244
R5122 gnd.n3800 gnd.n2467 240.244
R5123 gnd.n4228 gnd.n2467 240.244
R5124 gnd.n4228 gnd.n2475 240.244
R5125 gnd.n4243 gnd.n2475 240.244
R5126 gnd.n4243 gnd.n2484 240.244
R5127 gnd.n4250 gnd.n2484 240.244
R5128 gnd.n4250 gnd.n2492 240.244
R5129 gnd.n3784 gnd.n2492 240.244
R5130 gnd.n3784 gnd.n2501 240.244
R5131 gnd.n4292 gnd.n2501 240.244
R5132 gnd.n4292 gnd.n2512 240.244
R5133 gnd.n3769 gnd.n2512 240.244
R5134 gnd.n3769 gnd.n2521 240.244
R5135 gnd.n4299 gnd.n2521 240.244
R5136 gnd.n4299 gnd.n2532 240.244
R5137 gnd.n4304 gnd.n2532 240.244
R5138 gnd.n4304 gnd.n2541 240.244
R5139 gnd.n4309 gnd.n2541 240.244
R5140 gnd.n4309 gnd.n2552 240.244
R5141 gnd.n4313 gnd.n2552 240.244
R5142 gnd.n4313 gnd.n2562 240.244
R5143 gnd.n6161 gnd.n2562 240.244
R5144 gnd.n6161 gnd.n2572 240.244
R5145 gnd.n3975 gnd.n3970 240.244
R5146 gnd.n3981 gnd.n3970 240.244
R5147 gnd.n3985 gnd.n3983 240.244
R5148 gnd.n3991 gnd.n3966 240.244
R5149 gnd.n3995 gnd.n3993 240.244
R5150 gnd.n4001 gnd.n3962 240.244
R5151 gnd.n4005 gnd.n4003 240.244
R5152 gnd.n4011 gnd.n3958 240.244
R5153 gnd.n4015 gnd.n4013 240.244
R5154 gnd.n4021 gnd.n3951 240.244
R5155 gnd.n4025 gnd.n4023 240.244
R5156 gnd.n4031 gnd.n3947 240.244
R5157 gnd.n4035 gnd.n4033 240.244
R5158 gnd.n4041 gnd.n3943 240.244
R5159 gnd.n4045 gnd.n4043 240.244
R5160 gnd.n4051 gnd.n3939 240.244
R5161 gnd.n4055 gnd.n4053 240.244
R5162 gnd.n4061 gnd.n3935 240.244
R5163 gnd.n4065 gnd.n4063 240.244
R5164 gnd.n4073 gnd.n3931 240.244
R5165 gnd.n4077 gnd.n4075 240.244
R5166 gnd.n4083 gnd.n3927 240.244
R5167 gnd.n4087 gnd.n4085 240.244
R5168 gnd.n4093 gnd.n3923 240.244
R5169 gnd.n4097 gnd.n4095 240.244
R5170 gnd.n4103 gnd.n3919 240.244
R5171 gnd.n4107 gnd.n4105 240.244
R5172 gnd.n4114 gnd.n3915 240.244
R5173 gnd.n4117 gnd.n4116 240.244
R5174 gnd.n6295 gnd.n2369 240.244
R5175 gnd.n6291 gnd.n2369 240.244
R5176 gnd.n6291 gnd.n2374 240.244
R5177 gnd.n6283 gnd.n2374 240.244
R5178 gnd.n6283 gnd.n2390 240.244
R5179 gnd.n6279 gnd.n2390 240.244
R5180 gnd.n6279 gnd.n2396 240.244
R5181 gnd.n6271 gnd.n2396 240.244
R5182 gnd.n6271 gnd.n2411 240.244
R5183 gnd.n6267 gnd.n2411 240.244
R5184 gnd.n6267 gnd.n2417 240.244
R5185 gnd.n6259 gnd.n2417 240.244
R5186 gnd.n6259 gnd.n2431 240.244
R5187 gnd.n6255 gnd.n2431 240.244
R5188 gnd.n6255 gnd.n2437 240.244
R5189 gnd.n6247 gnd.n2437 240.244
R5190 gnd.n6247 gnd.n2452 240.244
R5191 gnd.n6242 gnd.n2452 240.244
R5192 gnd.n6242 gnd.n2456 240.244
R5193 gnd.n6234 gnd.n2456 240.244
R5194 gnd.n6234 gnd.n2470 240.244
R5195 gnd.n6229 gnd.n2470 240.244
R5196 gnd.n6229 gnd.n2473 240.244
R5197 gnd.n6221 gnd.n2473 240.244
R5198 gnd.n6221 gnd.n2487 240.244
R5199 gnd.n6216 gnd.n2487 240.244
R5200 gnd.n6216 gnd.n2490 240.244
R5201 gnd.n6208 gnd.n2490 240.244
R5202 gnd.n6208 gnd.n2504 240.244
R5203 gnd.n6204 gnd.n2504 240.244
R5204 gnd.n6204 gnd.n2510 240.244
R5205 gnd.n6196 gnd.n2510 240.244
R5206 gnd.n6196 gnd.n2524 240.244
R5207 gnd.n6192 gnd.n2524 240.244
R5208 gnd.n6192 gnd.n2530 240.244
R5209 gnd.n6184 gnd.n2530 240.244
R5210 gnd.n6184 gnd.n2544 240.244
R5211 gnd.n6180 gnd.n2544 240.244
R5212 gnd.n6180 gnd.n2550 240.244
R5213 gnd.n6172 gnd.n2550 240.244
R5214 gnd.n6172 gnd.n2565 240.244
R5215 gnd.n6168 gnd.n2565 240.244
R5216 gnd.n2337 gnd.n901 240.244
R5217 gnd.n2330 gnd.n2329 240.244
R5218 gnd.n2327 gnd.n2326 240.244
R5219 gnd.n2323 gnd.n2322 240.244
R5220 gnd.n2319 gnd.n2318 240.244
R5221 gnd.n2315 gnd.n2314 240.244
R5222 gnd.n2311 gnd.n2310 240.244
R5223 gnd.n2307 gnd.n2306 240.244
R5224 gnd.n1579 gnd.n1291 240.244
R5225 gnd.n1589 gnd.n1291 240.244
R5226 gnd.n1589 gnd.n1282 240.244
R5227 gnd.n1282 gnd.n1271 240.244
R5228 gnd.n1610 gnd.n1271 240.244
R5229 gnd.n1610 gnd.n1265 240.244
R5230 gnd.n1620 gnd.n1265 240.244
R5231 gnd.n1620 gnd.n1254 240.244
R5232 gnd.n1254 gnd.n1246 240.244
R5233 gnd.n1638 gnd.n1246 240.244
R5234 gnd.n1639 gnd.n1638 240.244
R5235 gnd.n1639 gnd.n1231 240.244
R5236 gnd.n1641 gnd.n1231 240.244
R5237 gnd.n1641 gnd.n1217 240.244
R5238 gnd.n1683 gnd.n1217 240.244
R5239 gnd.n1684 gnd.n1683 240.244
R5240 gnd.n1687 gnd.n1684 240.244
R5241 gnd.n1687 gnd.n1172 240.244
R5242 gnd.n1212 gnd.n1172 240.244
R5243 gnd.n1212 gnd.n1182 240.244
R5244 gnd.n1697 gnd.n1182 240.244
R5245 gnd.n1697 gnd.n1203 240.244
R5246 gnd.n1707 gnd.n1203 240.244
R5247 gnd.n1707 gnd.n1101 240.244
R5248 gnd.n1752 gnd.n1101 240.244
R5249 gnd.n1752 gnd.n1087 240.244
R5250 gnd.n1774 gnd.n1087 240.244
R5251 gnd.n1775 gnd.n1774 240.244
R5252 gnd.n1775 gnd.n1074 240.244
R5253 gnd.n1074 gnd.n1063 240.244
R5254 gnd.n1806 gnd.n1063 240.244
R5255 gnd.n1807 gnd.n1806 240.244
R5256 gnd.n1808 gnd.n1807 240.244
R5257 gnd.n1808 gnd.n1048 240.244
R5258 gnd.n1839 gnd.n1048 240.244
R5259 gnd.n1839 gnd.n1034 240.244
R5260 gnd.n1861 gnd.n1034 240.244
R5261 gnd.n1862 gnd.n1861 240.244
R5262 gnd.n1862 gnd.n1021 240.244
R5263 gnd.n1021 gnd.n1010 240.244
R5264 gnd.n1893 gnd.n1010 240.244
R5265 gnd.n1894 gnd.n1893 240.244
R5266 gnd.n1895 gnd.n1894 240.244
R5267 gnd.n1895 gnd.n994 240.244
R5268 gnd.n994 gnd.n993 240.244
R5269 gnd.n993 gnd.n980 240.244
R5270 gnd.n1950 gnd.n980 240.244
R5271 gnd.n1951 gnd.n1950 240.244
R5272 gnd.n1951 gnd.n967 240.244
R5273 gnd.n967 gnd.n957 240.244
R5274 gnd.n2238 gnd.n957 240.244
R5275 gnd.n2241 gnd.n2238 240.244
R5276 gnd.n2241 gnd.n2240 240.244
R5277 gnd.n1569 gnd.n1304 240.244
R5278 gnd.n1325 gnd.n1304 240.244
R5279 gnd.n1328 gnd.n1327 240.244
R5280 gnd.n1335 gnd.n1334 240.244
R5281 gnd.n1338 gnd.n1337 240.244
R5282 gnd.n1345 gnd.n1344 240.244
R5283 gnd.n1348 gnd.n1347 240.244
R5284 gnd.n1355 gnd.n1354 240.244
R5285 gnd.n1577 gnd.n1301 240.244
R5286 gnd.n1301 gnd.n1280 240.244
R5287 gnd.n1600 gnd.n1280 240.244
R5288 gnd.n1600 gnd.n1274 240.244
R5289 gnd.n1608 gnd.n1274 240.244
R5290 gnd.n1608 gnd.n1276 240.244
R5291 gnd.n1276 gnd.n1252 240.244
R5292 gnd.n1630 gnd.n1252 240.244
R5293 gnd.n1630 gnd.n1248 240.244
R5294 gnd.n1636 gnd.n1248 240.244
R5295 gnd.n1636 gnd.n1230 240.244
R5296 gnd.n1661 gnd.n1230 240.244
R5297 gnd.n1661 gnd.n1225 240.244
R5298 gnd.n1673 gnd.n1225 240.244
R5299 gnd.n1673 gnd.n1226 240.244
R5300 gnd.n1669 gnd.n1226 240.244
R5301 gnd.n1669 gnd.n1174 240.244
R5302 gnd.n1721 gnd.n1174 240.244
R5303 gnd.n1721 gnd.n1175 240.244
R5304 gnd.n1717 gnd.n1175 240.244
R5305 gnd.n1717 gnd.n1181 240.244
R5306 gnd.n1201 gnd.n1181 240.244
R5307 gnd.n1201 gnd.n1099 240.244
R5308 gnd.n1756 gnd.n1099 240.244
R5309 gnd.n1756 gnd.n1094 240.244
R5310 gnd.n1764 gnd.n1094 240.244
R5311 gnd.n1764 gnd.n1095 240.244
R5312 gnd.n1095 gnd.n1072 240.244
R5313 gnd.n1796 gnd.n1072 240.244
R5314 gnd.n1796 gnd.n1067 240.244
R5315 gnd.n1804 gnd.n1067 240.244
R5316 gnd.n1804 gnd.n1068 240.244
R5317 gnd.n1068 gnd.n1046 240.244
R5318 gnd.n1843 gnd.n1046 240.244
R5319 gnd.n1843 gnd.n1041 240.244
R5320 gnd.n1851 gnd.n1041 240.244
R5321 gnd.n1851 gnd.n1042 240.244
R5322 gnd.n1042 gnd.n1019 240.244
R5323 gnd.n1883 gnd.n1019 240.244
R5324 gnd.n1883 gnd.n1014 240.244
R5325 gnd.n1891 gnd.n1014 240.244
R5326 gnd.n1891 gnd.n1015 240.244
R5327 gnd.n1015 gnd.n992 240.244
R5328 gnd.n1932 gnd.n992 240.244
R5329 gnd.n1932 gnd.n987 240.244
R5330 gnd.n1940 gnd.n987 240.244
R5331 gnd.n1940 gnd.n988 240.244
R5332 gnd.n988 gnd.n965 240.244
R5333 gnd.n2226 gnd.n965 240.244
R5334 gnd.n2226 gnd.n960 240.244
R5335 gnd.n2236 gnd.n960 240.244
R5336 gnd.n2236 gnd.n961 240.244
R5337 gnd.n961 gnd.n900 240.244
R5338 gnd.n203 gnd.n172 240.244
R5339 gnd.n206 gnd.n205 240.244
R5340 gnd.n213 gnd.n212 240.244
R5341 gnd.n216 gnd.n215 240.244
R5342 gnd.n223 gnd.n222 240.244
R5343 gnd.n226 gnd.n225 240.244
R5344 gnd.n233 gnd.n232 240.244
R5345 gnd.n235 gnd.n192 240.244
R5346 gnd.n241 gnd.n183 240.244
R5347 gnd.n4994 gnd.n3022 240.244
R5348 gnd.n4994 gnd.n3034 240.244
R5349 gnd.n5573 gnd.n3034 240.244
R5350 gnd.n5573 gnd.n3046 240.244
R5351 gnd.n5579 gnd.n3046 240.244
R5352 gnd.n5579 gnd.n3057 240.244
R5353 gnd.n5599 gnd.n3057 240.244
R5354 gnd.n5599 gnd.n3066 240.244
R5355 gnd.n5590 gnd.n3066 240.244
R5356 gnd.n5590 gnd.n3077 240.244
R5357 gnd.n3211 gnd.n3077 240.244
R5358 gnd.n3211 gnd.n3086 240.244
R5359 gnd.n5653 gnd.n3086 240.244
R5360 gnd.n5653 gnd.n3097 240.244
R5361 gnd.n5669 gnd.n3097 240.244
R5362 gnd.n5669 gnd.n3106 240.244
R5363 gnd.n3112 gnd.n3106 240.244
R5364 gnd.n5658 gnd.n3112 240.244
R5365 gnd.n5659 gnd.n5658 240.244
R5366 gnd.n5659 gnd.n3122 240.244
R5367 gnd.n3129 gnd.n3122 240.244
R5368 gnd.n3129 gnd.n66 240.244
R5369 gnd.n7542 gnd.n66 240.244
R5370 gnd.n7542 gnd.n68 240.244
R5371 gnd.n5696 gnd.n68 240.244
R5372 gnd.n5696 gnd.n88 240.244
R5373 gnd.n5704 gnd.n88 240.244
R5374 gnd.n5704 gnd.n100 240.244
R5375 gnd.n5711 gnd.n100 240.244
R5376 gnd.n5711 gnd.n110 240.244
R5377 gnd.n5754 gnd.n110 240.244
R5378 gnd.n5754 gnd.n119 240.244
R5379 gnd.n5750 gnd.n119 240.244
R5380 gnd.n5750 gnd.n130 240.244
R5381 gnd.n5742 gnd.n130 240.244
R5382 gnd.n5742 gnd.n140 240.244
R5383 gnd.n5738 gnd.n140 240.244
R5384 gnd.n5738 gnd.n151 240.244
R5385 gnd.n5730 gnd.n151 240.244
R5386 gnd.n5730 gnd.n161 240.244
R5387 gnd.n7477 gnd.n161 240.244
R5388 gnd.n7477 gnd.n170 240.244
R5389 gnd.n5094 gnd.n5042 240.244
R5390 gnd.n5098 gnd.n5096 240.244
R5391 gnd.n5113 gnd.n5033 240.244
R5392 gnd.n5117 gnd.n5115 240.244
R5393 gnd.n5132 gnd.n5024 240.244
R5394 gnd.n5136 gnd.n5134 240.244
R5395 gnd.n5152 gnd.n5015 240.244
R5396 gnd.n5156 gnd.n5154 240.244
R5397 gnd.n5011 gnd.n5010 240.244
R5398 gnd.n3036 gnd.n3024 240.244
R5399 gnd.n5836 gnd.n3036 240.244
R5400 gnd.n5836 gnd.n3037 240.244
R5401 gnd.n5832 gnd.n3037 240.244
R5402 gnd.n5832 gnd.n3043 240.244
R5403 gnd.n5824 gnd.n3043 240.244
R5404 gnd.n5824 gnd.n3058 240.244
R5405 gnd.n5820 gnd.n3058 240.244
R5406 gnd.n5820 gnd.n3063 240.244
R5407 gnd.n5812 gnd.n3063 240.244
R5408 gnd.n5812 gnd.n3079 240.244
R5409 gnd.n5808 gnd.n3079 240.244
R5410 gnd.n5808 gnd.n3084 240.244
R5411 gnd.n5800 gnd.n3084 240.244
R5412 gnd.n5800 gnd.n3098 240.244
R5413 gnd.n5796 gnd.n3098 240.244
R5414 gnd.n5796 gnd.n3103 240.244
R5415 gnd.n5680 gnd.n3103 240.244
R5416 gnd.n5681 gnd.n5680 240.244
R5417 gnd.n5681 gnd.n3124 240.244
R5418 gnd.n5776 gnd.n3124 240.244
R5419 gnd.n5776 gnd.n3131 240.244
R5420 gnd.n3131 gnd.n72 240.244
R5421 gnd.n5771 gnd.n72 240.244
R5422 gnd.n5771 gnd.n90 240.244
R5423 gnd.n7532 gnd.n90 240.244
R5424 gnd.n7532 gnd.n91 240.244
R5425 gnd.n7528 gnd.n91 240.244
R5426 gnd.n7528 gnd.n97 240.244
R5427 gnd.n7520 gnd.n97 240.244
R5428 gnd.n7520 gnd.n111 240.244
R5429 gnd.n7516 gnd.n111 240.244
R5430 gnd.n7516 gnd.n116 240.244
R5431 gnd.n7508 gnd.n116 240.244
R5432 gnd.n7508 gnd.n132 240.244
R5433 gnd.n7504 gnd.n132 240.244
R5434 gnd.n7504 gnd.n137 240.244
R5435 gnd.n7496 gnd.n137 240.244
R5436 gnd.n7496 gnd.n153 240.244
R5437 gnd.n7492 gnd.n153 240.244
R5438 gnd.n7492 gnd.n158 240.244
R5439 gnd.n7484 gnd.n158 240.244
R5440 gnd.n920 gnd.n878 240.244
R5441 gnd.n2297 gnd.n2296 240.244
R5442 gnd.n2293 gnd.n2292 240.244
R5443 gnd.n2289 gnd.n2288 240.244
R5444 gnd.n2285 gnd.n2284 240.244
R5445 gnd.n2281 gnd.n2280 240.244
R5446 gnd.n2277 gnd.n2276 240.244
R5447 gnd.n2273 gnd.n2272 240.244
R5448 gnd.n2269 gnd.n2268 240.244
R5449 gnd.n2265 gnd.n2264 240.244
R5450 gnd.n2261 gnd.n2260 240.244
R5451 gnd.n2257 gnd.n2256 240.244
R5452 gnd.n2253 gnd.n2252 240.244
R5453 gnd.n1492 gnd.n1389 240.244
R5454 gnd.n1492 gnd.n1382 240.244
R5455 gnd.n1503 gnd.n1382 240.244
R5456 gnd.n1503 gnd.n1378 240.244
R5457 gnd.n1509 gnd.n1378 240.244
R5458 gnd.n1509 gnd.n1370 240.244
R5459 gnd.n1519 gnd.n1370 240.244
R5460 gnd.n1519 gnd.n1365 240.244
R5461 gnd.n1555 gnd.n1365 240.244
R5462 gnd.n1555 gnd.n1366 240.244
R5463 gnd.n1366 gnd.n1313 240.244
R5464 gnd.n1550 gnd.n1313 240.244
R5465 gnd.n1550 gnd.n1549 240.244
R5466 gnd.n1549 gnd.n1292 240.244
R5467 gnd.n1545 gnd.n1292 240.244
R5468 gnd.n1545 gnd.n1283 240.244
R5469 gnd.n1542 gnd.n1283 240.244
R5470 gnd.n1542 gnd.n1541 240.244
R5471 gnd.n1541 gnd.n1266 240.244
R5472 gnd.n1537 gnd.n1266 240.244
R5473 gnd.n1537 gnd.n1255 240.244
R5474 gnd.n1255 gnd.n1236 240.244
R5475 gnd.n1650 gnd.n1236 240.244
R5476 gnd.n1650 gnd.n1232 240.244
R5477 gnd.n1658 gnd.n1232 240.244
R5478 gnd.n1658 gnd.n1223 240.244
R5479 gnd.n1223 gnd.n1159 240.244
R5480 gnd.n1730 gnd.n1159 240.244
R5481 gnd.n1730 gnd.n1160 240.244
R5482 gnd.n1171 gnd.n1160 240.244
R5483 gnd.n1206 gnd.n1171 240.244
R5484 gnd.n1209 gnd.n1206 240.244
R5485 gnd.n1209 gnd.n1183 240.244
R5486 gnd.n1196 gnd.n1183 240.244
R5487 gnd.n1196 gnd.n1193 240.244
R5488 gnd.n1193 gnd.n1102 240.244
R5489 gnd.n1751 gnd.n1102 240.244
R5490 gnd.n1751 gnd.n1092 240.244
R5491 gnd.n1747 gnd.n1092 240.244
R5492 gnd.n1747 gnd.n1086 240.244
R5493 gnd.n1744 gnd.n1086 240.244
R5494 gnd.n1744 gnd.n1075 240.244
R5495 gnd.n1741 gnd.n1075 240.244
R5496 gnd.n1741 gnd.n1053 240.244
R5497 gnd.n1817 gnd.n1053 240.244
R5498 gnd.n1817 gnd.n1049 240.244
R5499 gnd.n1838 gnd.n1049 240.244
R5500 gnd.n1838 gnd.n1039 240.244
R5501 gnd.n1834 gnd.n1039 240.244
R5502 gnd.n1834 gnd.n1033 240.244
R5503 gnd.n1831 gnd.n1033 240.244
R5504 gnd.n1831 gnd.n1022 240.244
R5505 gnd.n1828 gnd.n1022 240.244
R5506 gnd.n1828 gnd.n999 240.244
R5507 gnd.n1904 gnd.n999 240.244
R5508 gnd.n1904 gnd.n995 240.244
R5509 gnd.n1929 gnd.n995 240.244
R5510 gnd.n1929 gnd.n986 240.244
R5511 gnd.n1925 gnd.n986 240.244
R5512 gnd.n1925 gnd.n979 240.244
R5513 gnd.n1921 gnd.n979 240.244
R5514 gnd.n1921 gnd.n968 240.244
R5515 gnd.n1918 gnd.n968 240.244
R5516 gnd.n1918 gnd.n949 240.244
R5517 gnd.n2248 gnd.n949 240.244
R5518 gnd.n1406 gnd.n1405 240.244
R5519 gnd.n1477 gnd.n1405 240.244
R5520 gnd.n1475 gnd.n1474 240.244
R5521 gnd.n1471 gnd.n1470 240.244
R5522 gnd.n1467 gnd.n1466 240.244
R5523 gnd.n1463 gnd.n1462 240.244
R5524 gnd.n1459 gnd.n1458 240.244
R5525 gnd.n1455 gnd.n1454 240.244
R5526 gnd.n1451 gnd.n1450 240.244
R5527 gnd.n1447 gnd.n1446 240.244
R5528 gnd.n1443 gnd.n1442 240.244
R5529 gnd.n1439 gnd.n1438 240.244
R5530 gnd.n1435 gnd.n1393 240.244
R5531 gnd.n1495 gnd.n1387 240.244
R5532 gnd.n1495 gnd.n1383 240.244
R5533 gnd.n1501 gnd.n1383 240.244
R5534 gnd.n1501 gnd.n1376 240.244
R5535 gnd.n1511 gnd.n1376 240.244
R5536 gnd.n1511 gnd.n1372 240.244
R5537 gnd.n1517 gnd.n1372 240.244
R5538 gnd.n1517 gnd.n1363 240.244
R5539 gnd.n1557 gnd.n1363 240.244
R5540 gnd.n1557 gnd.n1314 240.244
R5541 gnd.n1565 gnd.n1314 240.244
R5542 gnd.n1565 gnd.n1315 240.244
R5543 gnd.n1315 gnd.n1293 240.244
R5544 gnd.n1586 gnd.n1293 240.244
R5545 gnd.n1586 gnd.n1285 240.244
R5546 gnd.n1597 gnd.n1285 240.244
R5547 gnd.n1597 gnd.n1286 240.244
R5548 gnd.n1286 gnd.n1267 240.244
R5549 gnd.n1617 gnd.n1267 240.244
R5550 gnd.n1617 gnd.n1257 240.244
R5551 gnd.n1627 gnd.n1257 240.244
R5552 gnd.n1627 gnd.n1238 240.244
R5553 gnd.n1648 gnd.n1238 240.244
R5554 gnd.n1648 gnd.n1240 240.244
R5555 gnd.n1240 gnd.n1221 240.244
R5556 gnd.n1676 gnd.n1221 240.244
R5557 gnd.n1676 gnd.n1163 240.244
R5558 gnd.n1728 gnd.n1163 240.244
R5559 gnd.n1728 gnd.n1164 240.244
R5560 gnd.n1724 gnd.n1164 240.244
R5561 gnd.n1724 gnd.n1170 240.244
R5562 gnd.n1185 gnd.n1170 240.244
R5563 gnd.n1714 gnd.n1185 240.244
R5564 gnd.n1714 gnd.n1186 240.244
R5565 gnd.n1710 gnd.n1186 240.244
R5566 gnd.n1710 gnd.n1192 240.244
R5567 gnd.n1192 gnd.n1091 240.244
R5568 gnd.n1767 gnd.n1091 240.244
R5569 gnd.n1767 gnd.n1084 240.244
R5570 gnd.n1778 gnd.n1084 240.244
R5571 gnd.n1778 gnd.n1077 240.244
R5572 gnd.n1793 gnd.n1077 240.244
R5573 gnd.n1793 gnd.n1078 240.244
R5574 gnd.n1078 gnd.n1056 240.244
R5575 gnd.n1815 gnd.n1056 240.244
R5576 gnd.n1815 gnd.n1057 240.244
R5577 gnd.n1057 gnd.n1038 240.244
R5578 gnd.n1854 gnd.n1038 240.244
R5579 gnd.n1854 gnd.n1031 240.244
R5580 gnd.n1865 gnd.n1031 240.244
R5581 gnd.n1865 gnd.n1024 240.244
R5582 gnd.n1880 gnd.n1024 240.244
R5583 gnd.n1880 gnd.n1025 240.244
R5584 gnd.n1025 gnd.n1002 240.244
R5585 gnd.n1902 gnd.n1002 240.244
R5586 gnd.n1902 gnd.n1004 240.244
R5587 gnd.n1004 gnd.n984 240.244
R5588 gnd.n1943 gnd.n984 240.244
R5589 gnd.n1943 gnd.n977 240.244
R5590 gnd.n1954 gnd.n977 240.244
R5591 gnd.n1954 gnd.n970 240.244
R5592 gnd.n2223 gnd.n970 240.244
R5593 gnd.n2223 gnd.n971 240.244
R5594 gnd.n971 gnd.n952 240.244
R5595 gnd.n2246 gnd.n952 240.244
R5596 gnd.n2621 gnd.n2575 240.244
R5597 gnd.n2678 gnd.n2622 240.244
R5598 gnd.n2632 gnd.n2631 240.244
R5599 gnd.n2680 gnd.n2639 240.244
R5600 gnd.n2683 gnd.n2640 240.244
R5601 gnd.n2650 gnd.n2649 240.244
R5602 gnd.n2685 gnd.n2657 240.244
R5603 gnd.n2688 gnd.n2658 240.244
R5604 gnd.n2675 gnd.n2670 240.244
R5605 gnd.n4165 gnd.n2365 240.244
R5606 gnd.n4165 gnd.n2376 240.244
R5607 gnd.n4161 gnd.n2376 240.244
R5608 gnd.n4161 gnd.n2388 240.244
R5609 gnd.n4153 gnd.n2388 240.244
R5610 gnd.n4153 gnd.n2399 240.244
R5611 gnd.n4149 gnd.n2399 240.244
R5612 gnd.n4149 gnd.n2409 240.244
R5613 gnd.n4141 gnd.n2409 240.244
R5614 gnd.n4141 gnd.n2420 240.244
R5615 gnd.n4198 gnd.n2420 240.244
R5616 gnd.n4198 gnd.n2429 240.244
R5617 gnd.n4204 gnd.n2429 240.244
R5618 gnd.n4204 gnd.n2440 240.244
R5619 gnd.n4212 gnd.n2440 240.244
R5620 gnd.n4212 gnd.n2450 240.244
R5621 gnd.n4219 gnd.n2450 240.244
R5622 gnd.n4219 gnd.n2459 240.244
R5623 gnd.n4263 gnd.n2459 240.244
R5624 gnd.n4263 gnd.n2468 240.244
R5625 gnd.n3804 gnd.n2468 240.244
R5626 gnd.n3804 gnd.n2476 240.244
R5627 gnd.n3807 gnd.n2476 240.244
R5628 gnd.n3807 gnd.n2485 240.244
R5629 gnd.n4252 gnd.n2485 240.244
R5630 gnd.n4252 gnd.n2493 240.244
R5631 gnd.n4284 gnd.n2493 240.244
R5632 gnd.n4284 gnd.n2502 240.244
R5633 gnd.n4290 gnd.n2502 240.244
R5634 gnd.n4290 gnd.n2513 240.244
R5635 gnd.n4330 gnd.n2513 240.244
R5636 gnd.n4330 gnd.n2522 240.244
R5637 gnd.n3774 gnd.n2522 240.244
R5638 gnd.n3774 gnd.n2533 240.244
R5639 gnd.n3775 gnd.n2533 240.244
R5640 gnd.n3775 gnd.n2542 240.244
R5641 gnd.n3778 gnd.n2542 240.244
R5642 gnd.n3778 gnd.n2553 240.244
R5643 gnd.n4315 gnd.n2553 240.244
R5644 gnd.n4315 gnd.n2563 240.244
R5645 gnd.n6159 gnd.n2563 240.244
R5646 gnd.n6159 gnd.n2573 240.244
R5647 gnd.n3905 gnd.n3904 240.244
R5648 gnd.n3901 gnd.n3900 240.244
R5649 gnd.n3898 gnd.n3847 240.244
R5650 gnd.n3894 gnd.n3892 240.244
R5651 gnd.n3890 gnd.n3853 240.244
R5652 gnd.n3886 gnd.n3884 240.244
R5653 gnd.n3882 gnd.n3859 240.244
R5654 gnd.n3878 gnd.n3876 240.244
R5655 gnd.n3874 gnd.n3865 240.244
R5656 gnd.n2378 gnd.n2367 240.244
R5657 gnd.n6289 gnd.n2378 240.244
R5658 gnd.n6289 gnd.n2379 240.244
R5659 gnd.n6285 gnd.n2379 240.244
R5660 gnd.n6285 gnd.n2385 240.244
R5661 gnd.n6277 gnd.n2385 240.244
R5662 gnd.n6277 gnd.n2401 240.244
R5663 gnd.n6273 gnd.n2401 240.244
R5664 gnd.n6273 gnd.n2406 240.244
R5665 gnd.n6265 gnd.n2406 240.244
R5666 gnd.n6265 gnd.n2422 240.244
R5667 gnd.n6261 gnd.n2422 240.244
R5668 gnd.n6261 gnd.n2427 240.244
R5669 gnd.n6253 gnd.n2427 240.244
R5670 gnd.n6253 gnd.n2442 240.244
R5671 gnd.n6249 gnd.n2442 240.244
R5672 gnd.n6249 gnd.n2447 240.244
R5673 gnd.n6240 gnd.n2447 240.244
R5674 gnd.n6240 gnd.n2461 240.244
R5675 gnd.n6236 gnd.n2461 240.244
R5676 gnd.n6236 gnd.n2466 240.244
R5677 gnd.n6227 gnd.n2466 240.244
R5678 gnd.n6227 gnd.n2477 240.244
R5679 gnd.n6223 gnd.n2477 240.244
R5680 gnd.n6223 gnd.n2482 240.244
R5681 gnd.n6214 gnd.n2482 240.244
R5682 gnd.n6214 gnd.n2495 240.244
R5683 gnd.n6210 gnd.n2495 240.244
R5684 gnd.n6210 gnd.n2500 240.244
R5685 gnd.n6202 gnd.n2500 240.244
R5686 gnd.n6202 gnd.n2514 240.244
R5687 gnd.n6198 gnd.n2514 240.244
R5688 gnd.n6198 gnd.n2519 240.244
R5689 gnd.n6190 gnd.n2519 240.244
R5690 gnd.n6190 gnd.n2535 240.244
R5691 gnd.n6186 gnd.n2535 240.244
R5692 gnd.n6186 gnd.n2540 240.244
R5693 gnd.n6178 gnd.n2540 240.244
R5694 gnd.n6178 gnd.n2555 240.244
R5695 gnd.n6174 gnd.n2555 240.244
R5696 gnd.n6174 gnd.n2560 240.244
R5697 gnd.n6166 gnd.n2560 240.244
R5698 gnd.n6499 gnd.n704 240.244
R5699 gnd.n6503 gnd.n704 240.244
R5700 gnd.n6503 gnd.n700 240.244
R5701 gnd.n6509 gnd.n700 240.244
R5702 gnd.n6509 gnd.n698 240.244
R5703 gnd.n6513 gnd.n698 240.244
R5704 gnd.n6513 gnd.n694 240.244
R5705 gnd.n6519 gnd.n694 240.244
R5706 gnd.n6519 gnd.n692 240.244
R5707 gnd.n6523 gnd.n692 240.244
R5708 gnd.n6523 gnd.n688 240.244
R5709 gnd.n6529 gnd.n688 240.244
R5710 gnd.n6529 gnd.n686 240.244
R5711 gnd.n6533 gnd.n686 240.244
R5712 gnd.n6533 gnd.n682 240.244
R5713 gnd.n6539 gnd.n682 240.244
R5714 gnd.n6539 gnd.n680 240.244
R5715 gnd.n6543 gnd.n680 240.244
R5716 gnd.n6543 gnd.n676 240.244
R5717 gnd.n6549 gnd.n676 240.244
R5718 gnd.n6549 gnd.n674 240.244
R5719 gnd.n6553 gnd.n674 240.244
R5720 gnd.n6553 gnd.n670 240.244
R5721 gnd.n6559 gnd.n670 240.244
R5722 gnd.n6559 gnd.n668 240.244
R5723 gnd.n6563 gnd.n668 240.244
R5724 gnd.n6563 gnd.n664 240.244
R5725 gnd.n6569 gnd.n664 240.244
R5726 gnd.n6569 gnd.n662 240.244
R5727 gnd.n6573 gnd.n662 240.244
R5728 gnd.n6573 gnd.n658 240.244
R5729 gnd.n6579 gnd.n658 240.244
R5730 gnd.n6579 gnd.n656 240.244
R5731 gnd.n6583 gnd.n656 240.244
R5732 gnd.n6583 gnd.n652 240.244
R5733 gnd.n6589 gnd.n652 240.244
R5734 gnd.n6589 gnd.n650 240.244
R5735 gnd.n6593 gnd.n650 240.244
R5736 gnd.n6593 gnd.n646 240.244
R5737 gnd.n6599 gnd.n646 240.244
R5738 gnd.n6599 gnd.n644 240.244
R5739 gnd.n6603 gnd.n644 240.244
R5740 gnd.n6603 gnd.n640 240.244
R5741 gnd.n6609 gnd.n640 240.244
R5742 gnd.n6609 gnd.n638 240.244
R5743 gnd.n6613 gnd.n638 240.244
R5744 gnd.n6613 gnd.n634 240.244
R5745 gnd.n6619 gnd.n634 240.244
R5746 gnd.n6619 gnd.n632 240.244
R5747 gnd.n6623 gnd.n632 240.244
R5748 gnd.n6623 gnd.n628 240.244
R5749 gnd.n6629 gnd.n628 240.244
R5750 gnd.n6629 gnd.n626 240.244
R5751 gnd.n6633 gnd.n626 240.244
R5752 gnd.n6633 gnd.n622 240.244
R5753 gnd.n6639 gnd.n622 240.244
R5754 gnd.n6639 gnd.n620 240.244
R5755 gnd.n6643 gnd.n620 240.244
R5756 gnd.n6643 gnd.n616 240.244
R5757 gnd.n6649 gnd.n616 240.244
R5758 gnd.n6649 gnd.n614 240.244
R5759 gnd.n6653 gnd.n614 240.244
R5760 gnd.n6653 gnd.n610 240.244
R5761 gnd.n6659 gnd.n610 240.244
R5762 gnd.n6659 gnd.n608 240.244
R5763 gnd.n6663 gnd.n608 240.244
R5764 gnd.n6663 gnd.n604 240.244
R5765 gnd.n6669 gnd.n604 240.244
R5766 gnd.n6669 gnd.n602 240.244
R5767 gnd.n6673 gnd.n602 240.244
R5768 gnd.n6673 gnd.n598 240.244
R5769 gnd.n6679 gnd.n598 240.244
R5770 gnd.n6679 gnd.n596 240.244
R5771 gnd.n6683 gnd.n596 240.244
R5772 gnd.n6683 gnd.n592 240.244
R5773 gnd.n6689 gnd.n592 240.244
R5774 gnd.n6689 gnd.n590 240.244
R5775 gnd.n6693 gnd.n590 240.244
R5776 gnd.n6693 gnd.n586 240.244
R5777 gnd.n6699 gnd.n586 240.244
R5778 gnd.n6699 gnd.n584 240.244
R5779 gnd.n6703 gnd.n584 240.244
R5780 gnd.n6703 gnd.n580 240.244
R5781 gnd.n6709 gnd.n580 240.244
R5782 gnd.n6709 gnd.n578 240.244
R5783 gnd.n6713 gnd.n578 240.244
R5784 gnd.n6713 gnd.n574 240.244
R5785 gnd.n6719 gnd.n574 240.244
R5786 gnd.n6719 gnd.n572 240.244
R5787 gnd.n6723 gnd.n572 240.244
R5788 gnd.n6723 gnd.n568 240.244
R5789 gnd.n6729 gnd.n568 240.244
R5790 gnd.n6729 gnd.n566 240.244
R5791 gnd.n6733 gnd.n566 240.244
R5792 gnd.n6733 gnd.n562 240.244
R5793 gnd.n6739 gnd.n562 240.244
R5794 gnd.n6739 gnd.n560 240.244
R5795 gnd.n6743 gnd.n560 240.244
R5796 gnd.n6743 gnd.n556 240.244
R5797 gnd.n6749 gnd.n556 240.244
R5798 gnd.n6749 gnd.n554 240.244
R5799 gnd.n6753 gnd.n554 240.244
R5800 gnd.n6753 gnd.n550 240.244
R5801 gnd.n6759 gnd.n550 240.244
R5802 gnd.n6759 gnd.n548 240.244
R5803 gnd.n6763 gnd.n548 240.244
R5804 gnd.n6763 gnd.n544 240.244
R5805 gnd.n6769 gnd.n544 240.244
R5806 gnd.n6769 gnd.n542 240.244
R5807 gnd.n6773 gnd.n542 240.244
R5808 gnd.n6773 gnd.n538 240.244
R5809 gnd.n6779 gnd.n538 240.244
R5810 gnd.n6779 gnd.n536 240.244
R5811 gnd.n6783 gnd.n536 240.244
R5812 gnd.n6783 gnd.n532 240.244
R5813 gnd.n6789 gnd.n532 240.244
R5814 gnd.n6789 gnd.n530 240.244
R5815 gnd.n6793 gnd.n530 240.244
R5816 gnd.n6793 gnd.n526 240.244
R5817 gnd.n6799 gnd.n526 240.244
R5818 gnd.n6799 gnd.n524 240.244
R5819 gnd.n6803 gnd.n524 240.244
R5820 gnd.n6803 gnd.n520 240.244
R5821 gnd.n6809 gnd.n520 240.244
R5822 gnd.n6809 gnd.n518 240.244
R5823 gnd.n6813 gnd.n518 240.244
R5824 gnd.n6813 gnd.n514 240.244
R5825 gnd.n6819 gnd.n514 240.244
R5826 gnd.n6819 gnd.n512 240.244
R5827 gnd.n6823 gnd.n512 240.244
R5828 gnd.n6823 gnd.n508 240.244
R5829 gnd.n6829 gnd.n508 240.244
R5830 gnd.n6829 gnd.n506 240.244
R5831 gnd.n6833 gnd.n506 240.244
R5832 gnd.n6833 gnd.n502 240.244
R5833 gnd.n6839 gnd.n502 240.244
R5834 gnd.n6839 gnd.n500 240.244
R5835 gnd.n6843 gnd.n500 240.244
R5836 gnd.n6843 gnd.n496 240.244
R5837 gnd.n6849 gnd.n496 240.244
R5838 gnd.n6849 gnd.n494 240.244
R5839 gnd.n6853 gnd.n494 240.244
R5840 gnd.n6853 gnd.n490 240.244
R5841 gnd.n6859 gnd.n490 240.244
R5842 gnd.n6859 gnd.n488 240.244
R5843 gnd.n6863 gnd.n488 240.244
R5844 gnd.n6863 gnd.n484 240.244
R5845 gnd.n6869 gnd.n484 240.244
R5846 gnd.n6869 gnd.n482 240.244
R5847 gnd.n6873 gnd.n482 240.244
R5848 gnd.n6873 gnd.n478 240.244
R5849 gnd.n6879 gnd.n478 240.244
R5850 gnd.n6879 gnd.n476 240.244
R5851 gnd.n6883 gnd.n476 240.244
R5852 gnd.n6883 gnd.n472 240.244
R5853 gnd.n6889 gnd.n472 240.244
R5854 gnd.n6889 gnd.n470 240.244
R5855 gnd.n6893 gnd.n470 240.244
R5856 gnd.n6893 gnd.n466 240.244
R5857 gnd.n6899 gnd.n466 240.244
R5858 gnd.n6899 gnd.n464 240.244
R5859 gnd.n6903 gnd.n464 240.244
R5860 gnd.n6903 gnd.n460 240.244
R5861 gnd.n6909 gnd.n460 240.244
R5862 gnd.n6909 gnd.n458 240.244
R5863 gnd.n6913 gnd.n458 240.244
R5864 gnd.n6913 gnd.n454 240.244
R5865 gnd.n6919 gnd.n454 240.244
R5866 gnd.n6919 gnd.n452 240.244
R5867 gnd.n6923 gnd.n452 240.244
R5868 gnd.n6923 gnd.n448 240.244
R5869 gnd.n6929 gnd.n448 240.244
R5870 gnd.n6929 gnd.n446 240.244
R5871 gnd.n6933 gnd.n446 240.244
R5872 gnd.n6933 gnd.n442 240.244
R5873 gnd.n6939 gnd.n442 240.244
R5874 gnd.n6939 gnd.n440 240.244
R5875 gnd.n6943 gnd.n440 240.244
R5876 gnd.n6943 gnd.n436 240.244
R5877 gnd.n6949 gnd.n436 240.244
R5878 gnd.n6949 gnd.n434 240.244
R5879 gnd.n6953 gnd.n434 240.244
R5880 gnd.n6953 gnd.n430 240.244
R5881 gnd.n6959 gnd.n430 240.244
R5882 gnd.n6959 gnd.n428 240.244
R5883 gnd.n6963 gnd.n428 240.244
R5884 gnd.n6963 gnd.n424 240.244
R5885 gnd.n6969 gnd.n424 240.244
R5886 gnd.n6969 gnd.n422 240.244
R5887 gnd.n6973 gnd.n422 240.244
R5888 gnd.n6973 gnd.n418 240.244
R5889 gnd.n6979 gnd.n418 240.244
R5890 gnd.n6979 gnd.n416 240.244
R5891 gnd.n6983 gnd.n416 240.244
R5892 gnd.n6983 gnd.n412 240.244
R5893 gnd.n6989 gnd.n412 240.244
R5894 gnd.n6989 gnd.n410 240.244
R5895 gnd.n6993 gnd.n410 240.244
R5896 gnd.n6993 gnd.n406 240.244
R5897 gnd.n6999 gnd.n406 240.244
R5898 gnd.n6999 gnd.n404 240.244
R5899 gnd.n7003 gnd.n404 240.244
R5900 gnd.n7003 gnd.n400 240.244
R5901 gnd.n7010 gnd.n400 240.244
R5902 gnd.n7010 gnd.n398 240.244
R5903 gnd.n7014 gnd.n398 240.244
R5904 gnd.n7014 gnd.n395 240.244
R5905 gnd.n7020 gnd.n393 240.244
R5906 gnd.n7024 gnd.n393 240.244
R5907 gnd.n7024 gnd.n389 240.244
R5908 gnd.n7030 gnd.n389 240.244
R5909 gnd.n7030 gnd.n387 240.244
R5910 gnd.n7034 gnd.n387 240.244
R5911 gnd.n7034 gnd.n383 240.244
R5912 gnd.n7040 gnd.n383 240.244
R5913 gnd.n7040 gnd.n381 240.244
R5914 gnd.n7044 gnd.n381 240.244
R5915 gnd.n7044 gnd.n377 240.244
R5916 gnd.n7050 gnd.n377 240.244
R5917 gnd.n7050 gnd.n375 240.244
R5918 gnd.n7054 gnd.n375 240.244
R5919 gnd.n7054 gnd.n371 240.244
R5920 gnd.n7060 gnd.n371 240.244
R5921 gnd.n7060 gnd.n369 240.244
R5922 gnd.n7064 gnd.n369 240.244
R5923 gnd.n7064 gnd.n365 240.244
R5924 gnd.n7070 gnd.n365 240.244
R5925 gnd.n7070 gnd.n363 240.244
R5926 gnd.n7074 gnd.n363 240.244
R5927 gnd.n7074 gnd.n359 240.244
R5928 gnd.n7080 gnd.n359 240.244
R5929 gnd.n7080 gnd.n357 240.244
R5930 gnd.n7084 gnd.n357 240.244
R5931 gnd.n7084 gnd.n353 240.244
R5932 gnd.n7090 gnd.n353 240.244
R5933 gnd.n7090 gnd.n351 240.244
R5934 gnd.n7094 gnd.n351 240.244
R5935 gnd.n7094 gnd.n347 240.244
R5936 gnd.n7100 gnd.n347 240.244
R5937 gnd.n7100 gnd.n345 240.244
R5938 gnd.n7104 gnd.n345 240.244
R5939 gnd.n7104 gnd.n341 240.244
R5940 gnd.n7110 gnd.n341 240.244
R5941 gnd.n7110 gnd.n339 240.244
R5942 gnd.n7114 gnd.n339 240.244
R5943 gnd.n7114 gnd.n335 240.244
R5944 gnd.n7120 gnd.n335 240.244
R5945 gnd.n7120 gnd.n333 240.244
R5946 gnd.n7124 gnd.n333 240.244
R5947 gnd.n7124 gnd.n329 240.244
R5948 gnd.n7130 gnd.n329 240.244
R5949 gnd.n7130 gnd.n327 240.244
R5950 gnd.n7134 gnd.n327 240.244
R5951 gnd.n7134 gnd.n323 240.244
R5952 gnd.n7140 gnd.n323 240.244
R5953 gnd.n7140 gnd.n321 240.244
R5954 gnd.n7144 gnd.n321 240.244
R5955 gnd.n7144 gnd.n317 240.244
R5956 gnd.n7150 gnd.n317 240.244
R5957 gnd.n7150 gnd.n315 240.244
R5958 gnd.n7154 gnd.n315 240.244
R5959 gnd.n7154 gnd.n311 240.244
R5960 gnd.n7160 gnd.n311 240.244
R5961 gnd.n7160 gnd.n309 240.244
R5962 gnd.n7164 gnd.n309 240.244
R5963 gnd.n7164 gnd.n305 240.244
R5964 gnd.n7170 gnd.n305 240.244
R5965 gnd.n7170 gnd.n303 240.244
R5966 gnd.n7174 gnd.n303 240.244
R5967 gnd.n7174 gnd.n299 240.244
R5968 gnd.n7180 gnd.n299 240.244
R5969 gnd.n7180 gnd.n297 240.244
R5970 gnd.n7184 gnd.n297 240.244
R5971 gnd.n7184 gnd.n293 240.244
R5972 gnd.n7190 gnd.n293 240.244
R5973 gnd.n7190 gnd.n291 240.244
R5974 gnd.n7194 gnd.n291 240.244
R5975 gnd.n7194 gnd.n287 240.244
R5976 gnd.n7200 gnd.n287 240.244
R5977 gnd.n7200 gnd.n285 240.244
R5978 gnd.n7204 gnd.n285 240.244
R5979 gnd.n7204 gnd.n281 240.244
R5980 gnd.n7210 gnd.n281 240.244
R5981 gnd.n7210 gnd.n279 240.244
R5982 gnd.n7214 gnd.n279 240.244
R5983 gnd.n7214 gnd.n275 240.244
R5984 gnd.n7220 gnd.n275 240.244
R5985 gnd.n7220 gnd.n273 240.244
R5986 gnd.n7224 gnd.n273 240.244
R5987 gnd.n7224 gnd.n269 240.244
R5988 gnd.n7231 gnd.n269 240.244
R5989 gnd.n6323 gnd.n876 240.244
R5990 gnd.n6319 gnd.n876 240.244
R5991 gnd.n6319 gnd.n2341 240.244
R5992 gnd.n6315 gnd.n2341 240.244
R5993 gnd.n6315 gnd.n2346 240.244
R5994 gnd.n6311 gnd.n2346 240.244
R5995 gnd.n6311 gnd.n2348 240.244
R5996 gnd.n6307 gnd.n2348 240.244
R5997 gnd.n6307 gnd.n2354 240.244
R5998 gnd.n6303 gnd.n2354 240.244
R5999 gnd.n6303 gnd.n2356 240.244
R6000 gnd.n6299 gnd.n2356 240.244
R6001 gnd.n6299 gnd.n2362 240.244
R6002 gnd.n3833 gnd.n2362 240.244
R6003 gnd.n4168 gnd.n3833 240.244
R6004 gnd.n4168 gnd.n3828 240.244
R6005 gnd.n4174 gnd.n3828 240.244
R6006 gnd.n4175 gnd.n4174 240.244
R6007 gnd.n4176 gnd.n4175 240.244
R6008 gnd.n4176 gnd.n3824 240.244
R6009 gnd.n4182 gnd.n3824 240.244
R6010 gnd.n4183 gnd.n4182 240.244
R6011 gnd.n4184 gnd.n4183 240.244
R6012 gnd.n4184 gnd.n3819 240.244
R6013 gnd.n4195 gnd.n3819 240.244
R6014 gnd.n4195 gnd.n3820 240.244
R6015 gnd.n4191 gnd.n3820 240.244
R6016 gnd.n4191 gnd.n3796 240.244
R6017 gnd.n4272 gnd.n3796 240.244
R6018 gnd.n4272 gnd.n4271 240.244
R6019 gnd.n4271 gnd.n4270 240.244
R6020 gnd.n4270 gnd.n4267 240.244
R6021 gnd.n4267 gnd.n4266 240.244
R6022 gnd.n4266 gnd.n3797 240.244
R6023 gnd.n4231 gnd.n3797 240.244
R6024 gnd.n4240 gnd.n4231 240.244
R6025 gnd.n4240 gnd.n4237 240.244
R6026 gnd.n4237 gnd.n4234 240.244
R6027 gnd.n4234 gnd.n4233 240.244
R6028 gnd.n4233 gnd.n3785 240.244
R6029 gnd.n4281 gnd.n3785 240.244
R6030 gnd.n4281 gnd.n3786 240.244
R6031 gnd.n3786 gnd.n3768 240.244
R6032 gnd.n4333 gnd.n3768 240.244
R6033 gnd.n4333 gnd.n3764 240.244
R6034 gnd.n4339 gnd.n3764 240.244
R6035 gnd.n4340 gnd.n4339 240.244
R6036 gnd.n4341 gnd.n4340 240.244
R6037 gnd.n4341 gnd.n3760 240.244
R6038 gnd.n4347 gnd.n3760 240.244
R6039 gnd.n4348 gnd.n4347 240.244
R6040 gnd.n4349 gnd.n4348 240.244
R6041 gnd.n4349 gnd.n3756 240.244
R6042 gnd.n4355 gnd.n3756 240.244
R6043 gnd.n4356 gnd.n4355 240.244
R6044 gnd.n4357 gnd.n4356 240.244
R6045 gnd.n4357 gnd.n3752 240.244
R6046 gnd.n4363 gnd.n3752 240.244
R6047 gnd.n4365 gnd.n4363 240.244
R6048 gnd.n4366 gnd.n4365 240.244
R6049 gnd.n4366 gnd.n3748 240.244
R6050 gnd.n4372 gnd.n3748 240.244
R6051 gnd.n4372 gnd.n3747 240.244
R6052 gnd.n4394 gnd.n3747 240.244
R6053 gnd.n4394 gnd.n3742 240.244
R6054 gnd.n4402 gnd.n3742 240.244
R6055 gnd.n4402 gnd.n3743 240.244
R6056 gnd.n3743 gnd.n3722 240.244
R6057 gnd.n4424 gnd.n3722 240.244
R6058 gnd.n4424 gnd.n3717 240.244
R6059 gnd.n4432 gnd.n3717 240.244
R6060 gnd.n4432 gnd.n3718 240.244
R6061 gnd.n3718 gnd.n3697 240.244
R6062 gnd.n4454 gnd.n3697 240.244
R6063 gnd.n4454 gnd.n3692 240.244
R6064 gnd.n4472 gnd.n3692 240.244
R6065 gnd.n4472 gnd.n3693 240.244
R6066 gnd.n4468 gnd.n3693 240.244
R6067 gnd.n4468 gnd.n4467 240.244
R6068 gnd.n4467 gnd.n4465 240.244
R6069 gnd.n4465 gnd.n3603 240.244
R6070 gnd.n4529 gnd.n3603 240.244
R6071 gnd.n4529 gnd.n3598 240.244
R6072 gnd.n4537 gnd.n3598 240.244
R6073 gnd.n4537 gnd.n3599 240.244
R6074 gnd.n3599 gnd.n3577 240.244
R6075 gnd.n4591 gnd.n3577 240.244
R6076 gnd.n4591 gnd.n3573 240.244
R6077 gnd.n4597 gnd.n3573 240.244
R6078 gnd.n4597 gnd.n3559 240.244
R6079 gnd.n4618 gnd.n3559 240.244
R6080 gnd.n4618 gnd.n3554 240.244
R6081 gnd.n4626 gnd.n3554 240.244
R6082 gnd.n4626 gnd.n3555 240.244
R6083 gnd.n3555 gnd.n3526 240.244
R6084 gnd.n4669 gnd.n3526 240.244
R6085 gnd.n4669 gnd.n3522 240.244
R6086 gnd.n4675 gnd.n3522 240.244
R6087 gnd.n4675 gnd.n3503 240.244
R6088 gnd.n4709 gnd.n3503 240.244
R6089 gnd.n4709 gnd.n3499 240.244
R6090 gnd.n4715 gnd.n3499 240.244
R6091 gnd.n4715 gnd.n3481 240.244
R6092 gnd.n4765 gnd.n3481 240.244
R6093 gnd.n4765 gnd.n3477 240.244
R6094 gnd.n4771 gnd.n3477 240.244
R6095 gnd.n4771 gnd.n3462 240.244
R6096 gnd.n4790 gnd.n3462 240.244
R6097 gnd.n4790 gnd.n3458 240.244
R6098 gnd.n4796 gnd.n3458 240.244
R6099 gnd.n4796 gnd.n3442 240.244
R6100 gnd.n4850 gnd.n3442 240.244
R6101 gnd.n4850 gnd.n3438 240.244
R6102 gnd.n4856 gnd.n3438 240.244
R6103 gnd.n4856 gnd.n3420 240.244
R6104 gnd.n4879 gnd.n3420 240.244
R6105 gnd.n4879 gnd.n3415 240.244
R6106 gnd.n4887 gnd.n3415 240.244
R6107 gnd.n4887 gnd.n3416 240.244
R6108 gnd.n3416 gnd.n3392 240.244
R6109 gnd.n4924 gnd.n3392 240.244
R6110 gnd.n4924 gnd.n3387 240.244
R6111 gnd.n4936 gnd.n3387 240.244
R6112 gnd.n4936 gnd.n3388 240.244
R6113 gnd.n4932 gnd.n3388 240.244
R6114 gnd.n4932 gnd.n3313 240.244
R6115 gnd.n5223 gnd.n3313 240.244
R6116 gnd.n5223 gnd.n3314 240.244
R6117 gnd.n5219 gnd.n3314 240.244
R6118 gnd.n5219 gnd.n3320 240.244
R6119 gnd.n5212 gnd.n3320 240.244
R6120 gnd.n5212 gnd.n3324 240.244
R6121 gnd.n5208 gnd.n3324 240.244
R6122 gnd.n5208 gnd.n3330 240.244
R6123 gnd.n5201 gnd.n3330 240.244
R6124 gnd.n5201 gnd.n3336 240.244
R6125 gnd.n5197 gnd.n3336 240.244
R6126 gnd.n5197 gnd.n3342 240.244
R6127 gnd.n5190 gnd.n3342 240.244
R6128 gnd.n5190 gnd.n3348 240.244
R6129 gnd.n5186 gnd.n3348 240.244
R6130 gnd.n5186 gnd.n3354 240.244
R6131 gnd.n5179 gnd.n3354 240.244
R6132 gnd.n5179 gnd.n3003 240.244
R6133 gnd.n5857 gnd.n3003 240.244
R6134 gnd.n5857 gnd.n3004 240.244
R6135 gnd.n5853 gnd.n3004 240.244
R6136 gnd.n5853 gnd.n3010 240.244
R6137 gnd.n5849 gnd.n3010 240.244
R6138 gnd.n5849 gnd.n3013 240.244
R6139 gnd.n5845 gnd.n3013 240.244
R6140 gnd.n5845 gnd.n3019 240.244
R6141 gnd.n5609 gnd.n3019 240.244
R6142 gnd.n5609 gnd.n5606 240.244
R6143 gnd.n5615 gnd.n5606 240.244
R6144 gnd.n5616 gnd.n5615 240.244
R6145 gnd.n5617 gnd.n5616 240.244
R6146 gnd.n5617 gnd.n5602 240.244
R6147 gnd.n5623 gnd.n5602 240.244
R6148 gnd.n5624 gnd.n5623 240.244
R6149 gnd.n5625 gnd.n5624 240.244
R6150 gnd.n5625 gnd.n3212 240.244
R6151 gnd.n5643 gnd.n3212 240.244
R6152 gnd.n5643 gnd.n3213 240.244
R6153 gnd.n5639 gnd.n3213 240.244
R6154 gnd.n5639 gnd.n5638 240.244
R6155 gnd.n5638 gnd.n5637 240.244
R6156 gnd.n5637 gnd.n3114 240.244
R6157 gnd.n5789 gnd.n3114 240.244
R6158 gnd.n5789 gnd.n3115 240.244
R6159 gnd.n5784 gnd.n3115 240.244
R6160 gnd.n5784 gnd.n3118 240.244
R6161 gnd.n3142 gnd.n3118 240.244
R6162 gnd.n3143 gnd.n3142 240.244
R6163 gnd.n3143 gnd.n3138 240.244
R6164 gnd.n5768 gnd.n3138 240.244
R6165 gnd.n5768 gnd.n3139 240.244
R6166 gnd.n5763 gnd.n3139 240.244
R6167 gnd.n5763 gnd.n5762 240.244
R6168 gnd.n5762 gnd.n5761 240.244
R6169 gnd.n5761 gnd.n3149 240.244
R6170 gnd.n5757 gnd.n3149 240.244
R6171 gnd.n5757 gnd.n3190 240.244
R6172 gnd.n3190 gnd.n3189 240.244
R6173 gnd.n3189 gnd.n3155 240.244
R6174 gnd.n3185 gnd.n3155 240.244
R6175 gnd.n3185 gnd.n3184 240.244
R6176 gnd.n3184 gnd.n3183 240.244
R6177 gnd.n3183 gnd.n3161 240.244
R6178 gnd.n3179 gnd.n3161 240.244
R6179 gnd.n3179 gnd.n3178 240.244
R6180 gnd.n3178 gnd.n3177 240.244
R6181 gnd.n3177 gnd.n3167 240.244
R6182 gnd.n3173 gnd.n3167 240.244
R6183 gnd.n3173 gnd.n244 240.244
R6184 gnd.n7255 gnd.n244 240.244
R6185 gnd.n7255 gnd.n245 240.244
R6186 gnd.n7251 gnd.n245 240.244
R6187 gnd.n7251 gnd.n251 240.244
R6188 gnd.n7247 gnd.n251 240.244
R6189 gnd.n7247 gnd.n253 240.244
R6190 gnd.n7243 gnd.n253 240.244
R6191 gnd.n7243 gnd.n259 240.244
R6192 gnd.n7239 gnd.n259 240.244
R6193 gnd.n7239 gnd.n261 240.244
R6194 gnd.n7235 gnd.n261 240.244
R6195 gnd.n7235 gnd.n267 240.244
R6196 gnd.n6493 gnd.n706 240.244
R6197 gnd.n6493 gnd.n709 240.244
R6198 gnd.n6489 gnd.n709 240.244
R6199 gnd.n6489 gnd.n711 240.244
R6200 gnd.n6485 gnd.n711 240.244
R6201 gnd.n6485 gnd.n717 240.244
R6202 gnd.n6481 gnd.n717 240.244
R6203 gnd.n6481 gnd.n719 240.244
R6204 gnd.n6477 gnd.n719 240.244
R6205 gnd.n6477 gnd.n725 240.244
R6206 gnd.n6473 gnd.n725 240.244
R6207 gnd.n6473 gnd.n727 240.244
R6208 gnd.n6469 gnd.n727 240.244
R6209 gnd.n6469 gnd.n733 240.244
R6210 gnd.n6465 gnd.n733 240.244
R6211 gnd.n6465 gnd.n735 240.244
R6212 gnd.n6461 gnd.n735 240.244
R6213 gnd.n6461 gnd.n741 240.244
R6214 gnd.n6457 gnd.n741 240.244
R6215 gnd.n6457 gnd.n743 240.244
R6216 gnd.n6453 gnd.n743 240.244
R6217 gnd.n6453 gnd.n749 240.244
R6218 gnd.n6449 gnd.n749 240.244
R6219 gnd.n6449 gnd.n751 240.244
R6220 gnd.n6445 gnd.n751 240.244
R6221 gnd.n6445 gnd.n757 240.244
R6222 gnd.n6441 gnd.n757 240.244
R6223 gnd.n6441 gnd.n759 240.244
R6224 gnd.n6437 gnd.n759 240.244
R6225 gnd.n6437 gnd.n765 240.244
R6226 gnd.n6433 gnd.n765 240.244
R6227 gnd.n6433 gnd.n767 240.244
R6228 gnd.n6429 gnd.n767 240.244
R6229 gnd.n6429 gnd.n773 240.244
R6230 gnd.n6425 gnd.n773 240.244
R6231 gnd.n6425 gnd.n775 240.244
R6232 gnd.n6421 gnd.n775 240.244
R6233 gnd.n6421 gnd.n781 240.244
R6234 gnd.n6417 gnd.n781 240.244
R6235 gnd.n6417 gnd.n783 240.244
R6236 gnd.n6413 gnd.n783 240.244
R6237 gnd.n6413 gnd.n789 240.244
R6238 gnd.n6409 gnd.n789 240.244
R6239 gnd.n6409 gnd.n791 240.244
R6240 gnd.n6405 gnd.n791 240.244
R6241 gnd.n6405 gnd.n797 240.244
R6242 gnd.n6401 gnd.n797 240.244
R6243 gnd.n6401 gnd.n799 240.244
R6244 gnd.n6397 gnd.n799 240.244
R6245 gnd.n6397 gnd.n805 240.244
R6246 gnd.n6393 gnd.n805 240.244
R6247 gnd.n6393 gnd.n807 240.244
R6248 gnd.n6389 gnd.n807 240.244
R6249 gnd.n6389 gnd.n813 240.244
R6250 gnd.n6385 gnd.n813 240.244
R6251 gnd.n6385 gnd.n815 240.244
R6252 gnd.n6381 gnd.n815 240.244
R6253 gnd.n6381 gnd.n821 240.244
R6254 gnd.n6377 gnd.n821 240.244
R6255 gnd.n6377 gnd.n823 240.244
R6256 gnd.n6373 gnd.n823 240.244
R6257 gnd.n6373 gnd.n829 240.244
R6258 gnd.n6369 gnd.n829 240.244
R6259 gnd.n6369 gnd.n831 240.244
R6260 gnd.n6365 gnd.n831 240.244
R6261 gnd.n6365 gnd.n837 240.244
R6262 gnd.n6361 gnd.n837 240.244
R6263 gnd.n6361 gnd.n839 240.244
R6264 gnd.n6357 gnd.n839 240.244
R6265 gnd.n6357 gnd.n845 240.244
R6266 gnd.n6353 gnd.n845 240.244
R6267 gnd.n6353 gnd.n847 240.244
R6268 gnd.n6349 gnd.n847 240.244
R6269 gnd.n6349 gnd.n853 240.244
R6270 gnd.n6345 gnd.n853 240.244
R6271 gnd.n6345 gnd.n855 240.244
R6272 gnd.n6341 gnd.n855 240.244
R6273 gnd.n6341 gnd.n861 240.244
R6274 gnd.n6337 gnd.n861 240.244
R6275 gnd.n6337 gnd.n863 240.244
R6276 gnd.n6333 gnd.n863 240.244
R6277 gnd.n6333 gnd.n869 240.244
R6278 gnd.n6329 gnd.n869 240.244
R6279 gnd.n6329 gnd.n871 240.244
R6280 gnd.n4380 gnd.n2604 240.244
R6281 gnd.n4380 gnd.n3738 240.244
R6282 gnd.n4405 gnd.n3738 240.244
R6283 gnd.n4405 gnd.n3731 240.244
R6284 gnd.n4412 gnd.n3731 240.244
R6285 gnd.n4412 gnd.n3733 240.244
R6286 gnd.n3733 gnd.n3713 240.244
R6287 gnd.n4435 gnd.n3713 240.244
R6288 gnd.n4435 gnd.n3707 240.244
R6289 gnd.n4442 gnd.n3707 240.244
R6290 gnd.n4442 gnd.n3708 240.244
R6291 gnd.n3708 gnd.n3688 240.244
R6292 gnd.n4475 gnd.n3688 240.244
R6293 gnd.n4475 gnd.n3682 240.244
R6294 gnd.n4482 gnd.n3682 240.244
R6295 gnd.n4482 gnd.n3683 240.244
R6296 gnd.n3683 gnd.n2915 240.244
R6297 gnd.n5958 gnd.n2915 240.244
R6298 gnd.n5958 gnd.n2916 240.244
R6299 gnd.n2921 gnd.n2916 240.244
R6300 gnd.n2922 gnd.n2921 240.244
R6301 gnd.n2923 gnd.n2922 240.244
R6302 gnd.n4567 gnd.n2923 240.244
R6303 gnd.n4567 gnd.n2926 240.244
R6304 gnd.n2927 gnd.n2926 240.244
R6305 gnd.n2928 gnd.n2927 240.244
R6306 gnd.n4547 gnd.n2928 240.244
R6307 gnd.n4547 gnd.n2931 240.244
R6308 gnd.n2932 gnd.n2931 240.244
R6309 gnd.n2933 gnd.n2932 240.244
R6310 gnd.n4637 gnd.n2933 240.244
R6311 gnd.n4637 gnd.n2936 240.244
R6312 gnd.n2937 gnd.n2936 240.244
R6313 gnd.n2938 gnd.n2937 240.244
R6314 gnd.n4649 gnd.n2938 240.244
R6315 gnd.n4649 gnd.n2941 240.244
R6316 gnd.n2942 gnd.n2941 240.244
R6317 gnd.n2943 gnd.n2942 240.244
R6318 gnd.n4688 gnd.n2943 240.244
R6319 gnd.n4688 gnd.n2946 240.244
R6320 gnd.n2947 gnd.n2946 240.244
R6321 gnd.n2948 gnd.n2947 240.244
R6322 gnd.n4729 gnd.n2948 240.244
R6323 gnd.n4729 gnd.n2951 240.244
R6324 gnd.n2952 gnd.n2951 240.244
R6325 gnd.n2953 gnd.n2952 240.244
R6326 gnd.n4799 gnd.n2953 240.244
R6327 gnd.n4799 gnd.n2956 240.244
R6328 gnd.n2957 gnd.n2956 240.244
R6329 gnd.n2958 gnd.n2957 240.244
R6330 gnd.n4858 gnd.n2958 240.244
R6331 gnd.n4858 gnd.n2961 240.244
R6332 gnd.n2962 gnd.n2961 240.244
R6333 gnd.n2963 gnd.n2962 240.244
R6334 gnd.n4889 gnd.n2963 240.244
R6335 gnd.n4889 gnd.n2966 240.244
R6336 gnd.n2967 gnd.n2966 240.244
R6337 gnd.n2968 gnd.n2967 240.244
R6338 gnd.n4921 gnd.n2968 240.244
R6339 gnd.n4921 gnd.n2971 240.244
R6340 gnd.n2972 gnd.n2971 240.244
R6341 gnd.n2973 gnd.n2972 240.244
R6342 gnd.n4954 gnd.n2973 240.244
R6343 gnd.n4954 gnd.n2976 240.244
R6344 gnd.n2977 gnd.n2976 240.244
R6345 gnd.n2978 gnd.n2977 240.244
R6346 gnd.n5216 gnd.n2978 240.244
R6347 gnd.n5216 gnd.n2981 240.244
R6348 gnd.n2982 gnd.n2981 240.244
R6349 gnd.n2983 gnd.n2982 240.244
R6350 gnd.n5205 gnd.n2983 240.244
R6351 gnd.n5205 gnd.n2986 240.244
R6352 gnd.n2987 gnd.n2986 240.244
R6353 gnd.n2988 gnd.n2987 240.244
R6354 gnd.n5194 gnd.n2988 240.244
R6355 gnd.n5194 gnd.n2991 240.244
R6356 gnd.n2992 gnd.n2991 240.244
R6357 gnd.n2993 gnd.n2992 240.244
R6358 gnd.n5183 gnd.n2993 240.244
R6359 gnd.n5183 gnd.n2996 240.244
R6360 gnd.n2997 gnd.n2996 240.244
R6361 gnd.n5860 gnd.n2997 240.244
R6362 gnd.n2603 gnd.n2602 240.244
R6363 gnd.n2608 gnd.n2602 240.244
R6364 gnd.n2610 gnd.n2609 240.244
R6365 gnd.n2614 gnd.n2613 240.244
R6366 gnd.n2616 gnd.n2615 240.244
R6367 gnd.n2626 gnd.n2625 240.244
R6368 gnd.n2628 gnd.n2627 240.244
R6369 gnd.n2636 gnd.n2635 240.244
R6370 gnd.n2644 gnd.n2643 240.244
R6371 gnd.n2646 gnd.n2645 240.244
R6372 gnd.n2654 gnd.n2653 240.244
R6373 gnd.n2662 gnd.n2661 240.244
R6374 gnd.n2667 gnd.n2663 240.244
R6375 gnd.n2599 gnd.n2585 240.244
R6376 gnd.n4382 gnd.n2586 240.244
R6377 gnd.n4391 gnd.n4382 240.244
R6378 gnd.n4391 gnd.n3740 240.244
R6379 gnd.n3740 gnd.n3728 240.244
R6380 gnd.n4414 gnd.n3728 240.244
R6381 gnd.n4414 gnd.n3723 240.244
R6382 gnd.n4421 gnd.n3723 240.244
R6383 gnd.n4421 gnd.n3715 240.244
R6384 gnd.n3715 gnd.n3704 240.244
R6385 gnd.n4444 gnd.n3704 240.244
R6386 gnd.n4444 gnd.n3699 240.244
R6387 gnd.n4451 gnd.n3699 240.244
R6388 gnd.n4451 gnd.n3690 240.244
R6389 gnd.n3690 gnd.n3679 240.244
R6390 gnd.n4484 gnd.n3679 240.244
R6391 gnd.n4484 gnd.n3674 240.244
R6392 gnd.n4494 gnd.n3674 240.244
R6393 gnd.n4494 gnd.n2913 240.244
R6394 gnd.n4488 gnd.n2913 240.244
R6395 gnd.n4488 gnd.n3595 240.244
R6396 gnd.n4540 gnd.n3595 240.244
R6397 gnd.n4540 gnd.n3590 240.244
R6398 gnd.n4566 gnd.n3590 240.244
R6399 gnd.n4566 gnd.n3586 240.244
R6400 gnd.n3586 gnd.n3578 240.244
R6401 gnd.n4545 gnd.n3578 240.244
R6402 gnd.n4549 gnd.n4545 240.244
R6403 gnd.n4550 gnd.n4549 240.244
R6404 gnd.n4550 gnd.n3561 240.244
R6405 gnd.n3561 gnd.n3543 240.244
R6406 gnd.n4639 gnd.n3543 240.244
R6407 gnd.n4640 gnd.n4639 240.244
R6408 gnd.n4642 gnd.n4640 240.244
R6409 gnd.n4642 gnd.n3539 240.244
R6410 gnd.n4648 gnd.n3539 240.244
R6411 gnd.n4648 gnd.n3513 240.244
R6412 gnd.n4696 gnd.n3513 240.244
R6413 gnd.n4696 gnd.n3514 240.244
R6414 gnd.n4690 gnd.n3514 240.244
R6415 gnd.n4690 gnd.n3491 240.244
R6416 gnd.n4754 gnd.n3491 240.244
R6417 gnd.n4754 gnd.n3483 240.244
R6418 gnd.n4731 gnd.n3483 240.244
R6419 gnd.n4732 gnd.n4731 240.244
R6420 gnd.n4733 gnd.n4732 240.244
R6421 gnd.n4733 gnd.n3464 240.244
R6422 gnd.n3464 gnd.n3457 240.244
R6423 gnd.n4736 gnd.n3457 240.244
R6424 gnd.n4739 gnd.n4736 240.244
R6425 gnd.n4739 gnd.n3435 240.244
R6426 gnd.n4860 gnd.n3435 240.244
R6427 gnd.n4860 gnd.n3429 240.244
R6428 gnd.n4867 gnd.n3429 240.244
R6429 gnd.n4867 gnd.n3430 240.244
R6430 gnd.n3430 gnd.n3406 240.244
R6431 gnd.n4899 gnd.n3406 240.244
R6432 gnd.n4899 gnd.n3401 240.244
R6433 gnd.n4912 gnd.n3401 240.244
R6434 gnd.n4912 gnd.n3394 240.244
R6435 gnd.n4904 gnd.n3394 240.244
R6436 gnd.n4905 gnd.n4904 240.244
R6437 gnd.n4905 gnd.n3371 240.244
R6438 gnd.n4956 gnd.n3371 240.244
R6439 gnd.n4956 gnd.n3312 240.244
R6440 gnd.n4962 gnd.n3312 240.244
R6441 gnd.n4963 gnd.n4962 240.244
R6442 gnd.n4963 gnd.n3321 240.244
R6443 gnd.n3322 gnd.n3321 240.244
R6444 gnd.n4970 gnd.n3322 240.244
R6445 gnd.n4971 gnd.n4970 240.244
R6446 gnd.n4971 gnd.n3333 240.244
R6447 gnd.n3334 gnd.n3333 240.244
R6448 gnd.n4978 gnd.n3334 240.244
R6449 gnd.n4979 gnd.n4978 240.244
R6450 gnd.n4979 gnd.n3345 240.244
R6451 gnd.n3346 gnd.n3345 240.244
R6452 gnd.n4986 gnd.n3346 240.244
R6453 gnd.n4987 gnd.n4986 240.244
R6454 gnd.n4987 gnd.n3357 240.244
R6455 gnd.n3358 gnd.n3357 240.244
R6456 gnd.n5173 gnd.n3358 240.244
R6457 gnd.n5173 gnd.n3001 240.244
R6458 gnd.n5060 gnd.n5059 240.244
R6459 gnd.n5063 gnd.n5062 240.244
R6460 gnd.n5071 gnd.n5070 240.244
R6461 gnd.n5074 gnd.n5073 240.244
R6462 gnd.n5086 gnd.n5085 240.244
R6463 gnd.n5089 gnd.n5088 240.244
R6464 gnd.n5105 gnd.n5104 240.244
R6465 gnd.n5108 gnd.n5107 240.244
R6466 gnd.n5124 gnd.n5123 240.244
R6467 gnd.n5127 gnd.n5126 240.244
R6468 gnd.n5143 gnd.n5142 240.244
R6469 gnd.n5145 gnd.n5001 240.244
R6470 gnd.n5162 gnd.n5001 240.244
R6471 gnd.n5165 gnd.n5164 240.244
R6472 gnd.n2895 gnd.n2894 240.132
R6473 gnd.n5242 gnd.n5241 240.132
R6474 gnd.n6501 gnd.n6500 225.874
R6475 gnd.n6502 gnd.n6501 225.874
R6476 gnd.n6502 gnd.n699 225.874
R6477 gnd.n6510 gnd.n699 225.874
R6478 gnd.n6511 gnd.n6510 225.874
R6479 gnd.n6512 gnd.n6511 225.874
R6480 gnd.n6512 gnd.n693 225.874
R6481 gnd.n6520 gnd.n693 225.874
R6482 gnd.n6521 gnd.n6520 225.874
R6483 gnd.n6522 gnd.n6521 225.874
R6484 gnd.n6522 gnd.n687 225.874
R6485 gnd.n6530 gnd.n687 225.874
R6486 gnd.n6531 gnd.n6530 225.874
R6487 gnd.n6532 gnd.n6531 225.874
R6488 gnd.n6532 gnd.n681 225.874
R6489 gnd.n6540 gnd.n681 225.874
R6490 gnd.n6541 gnd.n6540 225.874
R6491 gnd.n6542 gnd.n6541 225.874
R6492 gnd.n6542 gnd.n675 225.874
R6493 gnd.n6550 gnd.n675 225.874
R6494 gnd.n6551 gnd.n6550 225.874
R6495 gnd.n6552 gnd.n6551 225.874
R6496 gnd.n6552 gnd.n669 225.874
R6497 gnd.n6560 gnd.n669 225.874
R6498 gnd.n6561 gnd.n6560 225.874
R6499 gnd.n6562 gnd.n6561 225.874
R6500 gnd.n6562 gnd.n663 225.874
R6501 gnd.n6570 gnd.n663 225.874
R6502 gnd.n6571 gnd.n6570 225.874
R6503 gnd.n6572 gnd.n6571 225.874
R6504 gnd.n6572 gnd.n657 225.874
R6505 gnd.n6580 gnd.n657 225.874
R6506 gnd.n6581 gnd.n6580 225.874
R6507 gnd.n6582 gnd.n6581 225.874
R6508 gnd.n6582 gnd.n651 225.874
R6509 gnd.n6590 gnd.n651 225.874
R6510 gnd.n6591 gnd.n6590 225.874
R6511 gnd.n6592 gnd.n6591 225.874
R6512 gnd.n6592 gnd.n645 225.874
R6513 gnd.n6600 gnd.n645 225.874
R6514 gnd.n6601 gnd.n6600 225.874
R6515 gnd.n6602 gnd.n6601 225.874
R6516 gnd.n6602 gnd.n639 225.874
R6517 gnd.n6610 gnd.n639 225.874
R6518 gnd.n6611 gnd.n6610 225.874
R6519 gnd.n6612 gnd.n6611 225.874
R6520 gnd.n6612 gnd.n633 225.874
R6521 gnd.n6620 gnd.n633 225.874
R6522 gnd.n6621 gnd.n6620 225.874
R6523 gnd.n6622 gnd.n6621 225.874
R6524 gnd.n6622 gnd.n627 225.874
R6525 gnd.n6630 gnd.n627 225.874
R6526 gnd.n6631 gnd.n6630 225.874
R6527 gnd.n6632 gnd.n6631 225.874
R6528 gnd.n6632 gnd.n621 225.874
R6529 gnd.n6640 gnd.n621 225.874
R6530 gnd.n6641 gnd.n6640 225.874
R6531 gnd.n6642 gnd.n6641 225.874
R6532 gnd.n6642 gnd.n615 225.874
R6533 gnd.n6650 gnd.n615 225.874
R6534 gnd.n6651 gnd.n6650 225.874
R6535 gnd.n6652 gnd.n6651 225.874
R6536 gnd.n6652 gnd.n609 225.874
R6537 gnd.n6660 gnd.n609 225.874
R6538 gnd.n6661 gnd.n6660 225.874
R6539 gnd.n6662 gnd.n6661 225.874
R6540 gnd.n6662 gnd.n603 225.874
R6541 gnd.n6670 gnd.n603 225.874
R6542 gnd.n6671 gnd.n6670 225.874
R6543 gnd.n6672 gnd.n6671 225.874
R6544 gnd.n6672 gnd.n597 225.874
R6545 gnd.n6680 gnd.n597 225.874
R6546 gnd.n6681 gnd.n6680 225.874
R6547 gnd.n6682 gnd.n6681 225.874
R6548 gnd.n6682 gnd.n591 225.874
R6549 gnd.n6690 gnd.n591 225.874
R6550 gnd.n6691 gnd.n6690 225.874
R6551 gnd.n6692 gnd.n6691 225.874
R6552 gnd.n6692 gnd.n585 225.874
R6553 gnd.n6700 gnd.n585 225.874
R6554 gnd.n6701 gnd.n6700 225.874
R6555 gnd.n6702 gnd.n6701 225.874
R6556 gnd.n6702 gnd.n579 225.874
R6557 gnd.n6710 gnd.n579 225.874
R6558 gnd.n6711 gnd.n6710 225.874
R6559 gnd.n6712 gnd.n6711 225.874
R6560 gnd.n6712 gnd.n573 225.874
R6561 gnd.n6720 gnd.n573 225.874
R6562 gnd.n6721 gnd.n6720 225.874
R6563 gnd.n6722 gnd.n6721 225.874
R6564 gnd.n6722 gnd.n567 225.874
R6565 gnd.n6730 gnd.n567 225.874
R6566 gnd.n6731 gnd.n6730 225.874
R6567 gnd.n6732 gnd.n6731 225.874
R6568 gnd.n6732 gnd.n561 225.874
R6569 gnd.n6740 gnd.n561 225.874
R6570 gnd.n6741 gnd.n6740 225.874
R6571 gnd.n6742 gnd.n6741 225.874
R6572 gnd.n6742 gnd.n555 225.874
R6573 gnd.n6750 gnd.n555 225.874
R6574 gnd.n6751 gnd.n6750 225.874
R6575 gnd.n6752 gnd.n6751 225.874
R6576 gnd.n6752 gnd.n549 225.874
R6577 gnd.n6760 gnd.n549 225.874
R6578 gnd.n6761 gnd.n6760 225.874
R6579 gnd.n6762 gnd.n6761 225.874
R6580 gnd.n6762 gnd.n543 225.874
R6581 gnd.n6770 gnd.n543 225.874
R6582 gnd.n6771 gnd.n6770 225.874
R6583 gnd.n6772 gnd.n6771 225.874
R6584 gnd.n6772 gnd.n537 225.874
R6585 gnd.n6780 gnd.n537 225.874
R6586 gnd.n6781 gnd.n6780 225.874
R6587 gnd.n6782 gnd.n6781 225.874
R6588 gnd.n6782 gnd.n531 225.874
R6589 gnd.n6790 gnd.n531 225.874
R6590 gnd.n6791 gnd.n6790 225.874
R6591 gnd.n6792 gnd.n6791 225.874
R6592 gnd.n6792 gnd.n525 225.874
R6593 gnd.n6800 gnd.n525 225.874
R6594 gnd.n6801 gnd.n6800 225.874
R6595 gnd.n6802 gnd.n6801 225.874
R6596 gnd.n6802 gnd.n519 225.874
R6597 gnd.n6810 gnd.n519 225.874
R6598 gnd.n6811 gnd.n6810 225.874
R6599 gnd.n6812 gnd.n6811 225.874
R6600 gnd.n6812 gnd.n513 225.874
R6601 gnd.n6820 gnd.n513 225.874
R6602 gnd.n6821 gnd.n6820 225.874
R6603 gnd.n6822 gnd.n6821 225.874
R6604 gnd.n6822 gnd.n507 225.874
R6605 gnd.n6830 gnd.n507 225.874
R6606 gnd.n6831 gnd.n6830 225.874
R6607 gnd.n6832 gnd.n6831 225.874
R6608 gnd.n6832 gnd.n501 225.874
R6609 gnd.n6840 gnd.n501 225.874
R6610 gnd.n6841 gnd.n6840 225.874
R6611 gnd.n6842 gnd.n6841 225.874
R6612 gnd.n6842 gnd.n495 225.874
R6613 gnd.n6850 gnd.n495 225.874
R6614 gnd.n6851 gnd.n6850 225.874
R6615 gnd.n6852 gnd.n6851 225.874
R6616 gnd.n6852 gnd.n489 225.874
R6617 gnd.n6860 gnd.n489 225.874
R6618 gnd.n6861 gnd.n6860 225.874
R6619 gnd.n6862 gnd.n6861 225.874
R6620 gnd.n6862 gnd.n483 225.874
R6621 gnd.n6870 gnd.n483 225.874
R6622 gnd.n6871 gnd.n6870 225.874
R6623 gnd.n6872 gnd.n6871 225.874
R6624 gnd.n6872 gnd.n477 225.874
R6625 gnd.n6880 gnd.n477 225.874
R6626 gnd.n6881 gnd.n6880 225.874
R6627 gnd.n6882 gnd.n6881 225.874
R6628 gnd.n6882 gnd.n471 225.874
R6629 gnd.n6890 gnd.n471 225.874
R6630 gnd.n6891 gnd.n6890 225.874
R6631 gnd.n6892 gnd.n6891 225.874
R6632 gnd.n6892 gnd.n465 225.874
R6633 gnd.n6900 gnd.n465 225.874
R6634 gnd.n6901 gnd.n6900 225.874
R6635 gnd.n6902 gnd.n6901 225.874
R6636 gnd.n6902 gnd.n459 225.874
R6637 gnd.n6910 gnd.n459 225.874
R6638 gnd.n6911 gnd.n6910 225.874
R6639 gnd.n6912 gnd.n6911 225.874
R6640 gnd.n6912 gnd.n453 225.874
R6641 gnd.n6920 gnd.n453 225.874
R6642 gnd.n6921 gnd.n6920 225.874
R6643 gnd.n6922 gnd.n6921 225.874
R6644 gnd.n6922 gnd.n447 225.874
R6645 gnd.n6930 gnd.n447 225.874
R6646 gnd.n6931 gnd.n6930 225.874
R6647 gnd.n6932 gnd.n6931 225.874
R6648 gnd.n6932 gnd.n441 225.874
R6649 gnd.n6940 gnd.n441 225.874
R6650 gnd.n6941 gnd.n6940 225.874
R6651 gnd.n6942 gnd.n6941 225.874
R6652 gnd.n6942 gnd.n435 225.874
R6653 gnd.n6950 gnd.n435 225.874
R6654 gnd.n6951 gnd.n6950 225.874
R6655 gnd.n6952 gnd.n6951 225.874
R6656 gnd.n6952 gnd.n429 225.874
R6657 gnd.n6960 gnd.n429 225.874
R6658 gnd.n6961 gnd.n6960 225.874
R6659 gnd.n6962 gnd.n6961 225.874
R6660 gnd.n6962 gnd.n423 225.874
R6661 gnd.n6970 gnd.n423 225.874
R6662 gnd.n6971 gnd.n6970 225.874
R6663 gnd.n6972 gnd.n6971 225.874
R6664 gnd.n6972 gnd.n417 225.874
R6665 gnd.n6980 gnd.n417 225.874
R6666 gnd.n6981 gnd.n6980 225.874
R6667 gnd.n6982 gnd.n6981 225.874
R6668 gnd.n6982 gnd.n411 225.874
R6669 gnd.n6990 gnd.n411 225.874
R6670 gnd.n6991 gnd.n6990 225.874
R6671 gnd.n6992 gnd.n6991 225.874
R6672 gnd.n6992 gnd.n405 225.874
R6673 gnd.n7000 gnd.n405 225.874
R6674 gnd.n7001 gnd.n7000 225.874
R6675 gnd.n7002 gnd.n7001 225.874
R6676 gnd.n7002 gnd.n399 225.874
R6677 gnd.n7011 gnd.n399 225.874
R6678 gnd.n7012 gnd.n7011 225.874
R6679 gnd.n7013 gnd.n7012 225.874
R6680 gnd.n7013 gnd.n394 225.874
R6681 gnd.n1430 gnd.t185 224.174
R6682 gnd.n942 gnd.t180 224.174
R6683 gnd.n5483 gnd.n5482 199.319
R6684 gnd.n5484 gnd.n5483 199.319
R6685 gnd.n2752 gnd.n2707 199.319
R6686 gnd.n2752 gnd.n2706 199.319
R6687 gnd.n2896 gnd.n2893 186.49
R6688 gnd.n5243 gnd.n5240 186.49
R6689 gnd.n2207 gnd.n2206 185
R6690 gnd.n2205 gnd.n2204 185
R6691 gnd.n2184 gnd.n2183 185
R6692 gnd.n2199 gnd.n2198 185
R6693 gnd.n2197 gnd.n2196 185
R6694 gnd.n2188 gnd.n2187 185
R6695 gnd.n2191 gnd.n2190 185
R6696 gnd.n2175 gnd.n2174 185
R6697 gnd.n2173 gnd.n2172 185
R6698 gnd.n2152 gnd.n2151 185
R6699 gnd.n2167 gnd.n2166 185
R6700 gnd.n2165 gnd.n2164 185
R6701 gnd.n2156 gnd.n2155 185
R6702 gnd.n2159 gnd.n2158 185
R6703 gnd.n2143 gnd.n2142 185
R6704 gnd.n2141 gnd.n2140 185
R6705 gnd.n2120 gnd.n2119 185
R6706 gnd.n2135 gnd.n2134 185
R6707 gnd.n2133 gnd.n2132 185
R6708 gnd.n2124 gnd.n2123 185
R6709 gnd.n2127 gnd.n2126 185
R6710 gnd.n2112 gnd.n2111 185
R6711 gnd.n2110 gnd.n2109 185
R6712 gnd.n2089 gnd.n2088 185
R6713 gnd.n2104 gnd.n2103 185
R6714 gnd.n2102 gnd.n2101 185
R6715 gnd.n2093 gnd.n2092 185
R6716 gnd.n2096 gnd.n2095 185
R6717 gnd.n2080 gnd.n2079 185
R6718 gnd.n2078 gnd.n2077 185
R6719 gnd.n2057 gnd.n2056 185
R6720 gnd.n2072 gnd.n2071 185
R6721 gnd.n2070 gnd.n2069 185
R6722 gnd.n2061 gnd.n2060 185
R6723 gnd.n2064 gnd.n2063 185
R6724 gnd.n2048 gnd.n2047 185
R6725 gnd.n2046 gnd.n2045 185
R6726 gnd.n2025 gnd.n2024 185
R6727 gnd.n2040 gnd.n2039 185
R6728 gnd.n2038 gnd.n2037 185
R6729 gnd.n2029 gnd.n2028 185
R6730 gnd.n2032 gnd.n2031 185
R6731 gnd.n2016 gnd.n2015 185
R6732 gnd.n2014 gnd.n2013 185
R6733 gnd.n1993 gnd.n1992 185
R6734 gnd.n2008 gnd.n2007 185
R6735 gnd.n2006 gnd.n2005 185
R6736 gnd.n1997 gnd.n1996 185
R6737 gnd.n2000 gnd.n1999 185
R6738 gnd.n1985 gnd.n1984 185
R6739 gnd.n1983 gnd.n1982 185
R6740 gnd.n1962 gnd.n1961 185
R6741 gnd.n1977 gnd.n1976 185
R6742 gnd.n1975 gnd.n1974 185
R6743 gnd.n1966 gnd.n1965 185
R6744 gnd.n1969 gnd.n1968 185
R6745 gnd.n1431 gnd.t184 178.987
R6746 gnd.n943 gnd.t181 178.987
R6747 gnd.n1 gnd.t305 170.774
R6748 gnd.n7 gnd.t317 170.103
R6749 gnd.n6 gnd.t309 170.103
R6750 gnd.n5 gnd.t103 170.103
R6751 gnd.n4 gnd.t315 170.103
R6752 gnd.n3 gnd.t106 170.103
R6753 gnd.n2 gnd.t88 170.103
R6754 gnd.n1 gnd.t76 170.103
R6755 gnd.n5311 gnd.n5310 163.367
R6756 gnd.n5307 gnd.n5306 163.367
R6757 gnd.n5303 gnd.n5302 163.367
R6758 gnd.n5299 gnd.n5298 163.367
R6759 gnd.n5295 gnd.n5294 163.367
R6760 gnd.n5291 gnd.n5290 163.367
R6761 gnd.n5287 gnd.n5286 163.367
R6762 gnd.n5283 gnd.n5282 163.367
R6763 gnd.n5279 gnd.n5278 163.367
R6764 gnd.n5275 gnd.n5274 163.367
R6765 gnd.n5271 gnd.n5270 163.367
R6766 gnd.n5267 gnd.n5266 163.367
R6767 gnd.n5263 gnd.n5262 163.367
R6768 gnd.n5259 gnd.n5258 163.367
R6769 gnd.n5254 gnd.n5253 163.367
R6770 gnd.n5386 gnd.n3266 163.367
R6771 gnd.n5383 gnd.n5382 163.367
R6772 gnd.n5380 gnd.n3299 163.367
R6773 gnd.n5375 gnd.n5374 163.367
R6774 gnd.n5371 gnd.n5370 163.367
R6775 gnd.n5367 gnd.n5366 163.367
R6776 gnd.n5363 gnd.n5362 163.367
R6777 gnd.n5359 gnd.n5358 163.367
R6778 gnd.n5355 gnd.n5354 163.367
R6779 gnd.n5351 gnd.n5350 163.367
R6780 gnd.n5347 gnd.n5346 163.367
R6781 gnd.n5343 gnd.n5342 163.367
R6782 gnd.n5339 gnd.n5338 163.367
R6783 gnd.n5335 gnd.n5334 163.367
R6784 gnd.n5331 gnd.n5330 163.367
R6785 gnd.n5327 gnd.n5326 163.367
R6786 gnd.n5323 gnd.n5322 163.367
R6787 gnd.n4497 gnd.n2912 163.367
R6788 gnd.n4501 gnd.n2912 163.367
R6789 gnd.n4504 gnd.n4501 163.367
R6790 gnd.n4504 gnd.n3605 163.367
R6791 gnd.n4511 gnd.n3605 163.367
R6792 gnd.n4511 gnd.n3608 163.367
R6793 gnd.n4507 gnd.n3608 163.367
R6794 gnd.n4507 gnd.n3588 163.367
R6795 gnd.n4570 gnd.n3588 163.367
R6796 gnd.n4570 gnd.n3585 163.367
R6797 gnd.n4579 gnd.n3585 163.367
R6798 gnd.n4579 gnd.n3579 163.367
R6799 gnd.n4575 gnd.n3579 163.367
R6800 gnd.n4575 gnd.n3572 163.367
R6801 gnd.n3572 gnd.n3564 163.367
R6802 gnd.n4607 gnd.n3564 163.367
R6803 gnd.n4607 gnd.n3562 163.367
R6804 gnd.n4614 gnd.n3562 163.367
R6805 gnd.n4614 gnd.n3552 163.367
R6806 gnd.n3553 gnd.n3552 163.367
R6807 gnd.n3553 gnd.n3545 163.367
R6808 gnd.n3545 gnd.n3535 163.367
R6809 gnd.n4657 gnd.n3535 163.367
R6810 gnd.n4657 gnd.n3536 163.367
R6811 gnd.n3536 gnd.n3528 163.367
R6812 gnd.n4652 gnd.n3528 163.367
R6813 gnd.n4652 gnd.n3520 163.367
R6814 gnd.n4679 gnd.n3520 163.367
R6815 gnd.n4679 gnd.n3512 163.367
R6816 gnd.n4682 gnd.n3512 163.367
R6817 gnd.n4682 gnd.n3505 163.367
R6818 gnd.n4686 gnd.n3505 163.367
R6819 gnd.n4686 gnd.n3497 163.367
R6820 gnd.n4719 gnd.n3497 163.367
R6821 gnd.n4719 gnd.n3490 163.367
R6822 gnd.n4722 gnd.n3490 163.367
R6823 gnd.n4722 gnd.n3484 163.367
R6824 gnd.n4727 gnd.n3484 163.367
R6825 gnd.n4727 gnd.n3474 163.367
R6826 gnd.n3474 gnd.n3467 163.367
R6827 gnd.n4781 gnd.n3467 163.367
R6828 gnd.n4781 gnd.n3465 163.367
R6829 gnd.n4786 gnd.n3465 163.367
R6830 gnd.n4786 gnd.n3456 163.367
R6831 gnd.n3456 gnd.n3448 163.367
R6832 gnd.n4816 gnd.n3448 163.367
R6833 gnd.n4816 gnd.n3445 163.367
R6834 gnd.n4848 gnd.n3445 163.367
R6835 gnd.n4848 gnd.n3446 163.367
R6836 gnd.n4844 gnd.n3446 163.367
R6837 gnd.n4844 gnd.n4843 163.367
R6838 gnd.n4843 gnd.n3427 163.367
R6839 gnd.n3428 gnd.n3427 163.367
R6840 gnd.n3428 gnd.n3421 163.367
R6841 gnd.n4837 gnd.n3421 163.367
R6842 gnd.n4837 gnd.n3414 163.367
R6843 gnd.n4833 gnd.n3414 163.367
R6844 gnd.n4833 gnd.n3408 163.367
R6845 gnd.n4830 gnd.n3408 163.367
R6846 gnd.n4830 gnd.n3400 163.367
R6847 gnd.n4824 gnd.n3400 163.367
R6848 gnd.n4824 gnd.n3395 163.367
R6849 gnd.n4821 gnd.n3395 163.367
R6850 gnd.n4821 gnd.n3384 163.367
R6851 gnd.n3384 gnd.n3375 163.367
R6852 gnd.n4946 gnd.n3375 163.367
R6853 gnd.n4946 gnd.n3373 163.367
R6854 gnd.n4952 gnd.n3373 163.367
R6855 gnd.n4952 gnd.n3311 163.367
R6856 gnd.n3311 gnd.n3303 163.367
R6857 gnd.n5318 gnd.n3303 163.367
R6858 gnd.n2887 gnd.n2886 163.367
R6859 gnd.n6023 gnd.n2886 163.367
R6860 gnd.n6021 gnd.n6020 163.367
R6861 gnd.n6017 gnd.n6016 163.367
R6862 gnd.n6013 gnd.n6012 163.367
R6863 gnd.n6009 gnd.n6008 163.367
R6864 gnd.n6005 gnd.n6004 163.367
R6865 gnd.n6001 gnd.n6000 163.367
R6866 gnd.n5997 gnd.n5996 163.367
R6867 gnd.n5993 gnd.n5992 163.367
R6868 gnd.n5989 gnd.n5988 163.367
R6869 gnd.n5985 gnd.n5984 163.367
R6870 gnd.n5981 gnd.n5980 163.367
R6871 gnd.n5977 gnd.n5976 163.367
R6872 gnd.n5973 gnd.n5972 163.367
R6873 gnd.n5969 gnd.n5968 163.367
R6874 gnd.n6032 gnd.n2853 163.367
R6875 gnd.n3613 gnd.n3612 163.367
R6876 gnd.n3618 gnd.n3617 163.367
R6877 gnd.n3622 gnd.n3621 163.367
R6878 gnd.n3626 gnd.n3625 163.367
R6879 gnd.n3630 gnd.n3629 163.367
R6880 gnd.n3634 gnd.n3633 163.367
R6881 gnd.n3638 gnd.n3637 163.367
R6882 gnd.n3642 gnd.n3641 163.367
R6883 gnd.n3646 gnd.n3645 163.367
R6884 gnd.n3650 gnd.n3649 163.367
R6885 gnd.n3654 gnd.n3653 163.367
R6886 gnd.n3658 gnd.n3657 163.367
R6887 gnd.n3662 gnd.n3661 163.367
R6888 gnd.n3666 gnd.n3665 163.367
R6889 gnd.n3670 gnd.n3669 163.367
R6890 gnd.n5961 gnd.n2888 163.367
R6891 gnd.n5961 gnd.n2910 163.367
R6892 gnd.n3607 gnd.n2910 163.367
R6893 gnd.n4526 gnd.n3607 163.367
R6894 gnd.n4526 gnd.n4514 163.367
R6895 gnd.n4522 gnd.n4514 163.367
R6896 gnd.n4522 gnd.n4521 163.367
R6897 gnd.n4521 gnd.n4520 163.367
R6898 gnd.n4520 gnd.n3583 163.367
R6899 gnd.n4583 gnd.n3583 163.367
R6900 gnd.n4583 gnd.n3581 163.367
R6901 gnd.n4587 gnd.n3581 163.367
R6902 gnd.n4587 gnd.n3570 163.367
R6903 gnd.n4600 gnd.n3570 163.367
R6904 gnd.n4600 gnd.n3567 163.367
R6905 gnd.n4605 gnd.n3567 163.367
R6906 gnd.n4605 gnd.n3568 163.367
R6907 gnd.n3568 gnd.n3550 163.367
R6908 gnd.n4631 gnd.n3550 163.367
R6909 gnd.n4631 gnd.n3548 163.367
R6910 gnd.n4635 gnd.n3548 163.367
R6911 gnd.n4635 gnd.n3533 163.367
R6912 gnd.n4659 gnd.n3533 163.367
R6913 gnd.n4659 gnd.n3530 163.367
R6914 gnd.n4666 gnd.n3530 163.367
R6915 gnd.n4666 gnd.n3531 163.367
R6916 gnd.n4662 gnd.n3531 163.367
R6917 gnd.n4662 gnd.n3510 163.367
R6918 gnd.n4699 gnd.n3510 163.367
R6919 gnd.n4699 gnd.n3507 163.367
R6920 gnd.n4706 gnd.n3507 163.367
R6921 gnd.n4706 gnd.n3508 163.367
R6922 gnd.n4702 gnd.n3508 163.367
R6923 gnd.n4702 gnd.n3488 163.367
R6924 gnd.n4757 gnd.n3488 163.367
R6925 gnd.n4757 gnd.n3486 163.367
R6926 gnd.n4761 gnd.n3486 163.367
R6927 gnd.n4761 gnd.n3473 163.367
R6928 gnd.n4774 gnd.n3473 163.367
R6929 gnd.n4774 gnd.n3470 163.367
R6930 gnd.n4779 gnd.n3470 163.367
R6931 gnd.n4779 gnd.n3471 163.367
R6932 gnd.n3471 gnd.n3454 163.367
R6933 gnd.n4802 gnd.n3454 163.367
R6934 gnd.n4802 gnd.n3451 163.367
R6935 gnd.n4814 gnd.n3451 163.367
R6936 gnd.n4814 gnd.n3452 163.367
R6937 gnd.n3452 gnd.n3443 163.367
R6938 gnd.n4809 gnd.n3443 163.367
R6939 gnd.n4809 gnd.n4806 163.367
R6940 gnd.n4806 gnd.n3425 163.367
R6941 gnd.n4872 gnd.n3425 163.367
R6942 gnd.n4872 gnd.n3423 163.367
R6943 gnd.n4876 gnd.n3423 163.367
R6944 gnd.n4876 gnd.n3412 163.367
R6945 gnd.n4892 gnd.n3412 163.367
R6946 gnd.n4892 gnd.n3410 163.367
R6947 gnd.n4896 gnd.n3410 163.367
R6948 gnd.n4896 gnd.n3399 163.367
R6949 gnd.n4915 gnd.n3399 163.367
R6950 gnd.n4915 gnd.n3397 163.367
R6951 gnd.n4919 gnd.n3397 163.367
R6952 gnd.n4919 gnd.n3382 163.367
R6953 gnd.n4939 gnd.n3382 163.367
R6954 gnd.n4939 gnd.n3377 163.367
R6955 gnd.n4944 gnd.n3377 163.367
R6956 gnd.n4944 gnd.n3380 163.367
R6957 gnd.n3380 gnd.n3309 163.367
R6958 gnd.n5228 gnd.n3309 163.367
R6959 gnd.n5228 gnd.n3306 163.367
R6960 gnd.n5316 gnd.n3306 163.367
R6961 gnd.n5249 gnd.n5248 156.462
R6962 gnd.n2147 gnd.n2115 153.042
R6963 gnd.n2211 gnd.n2210 152.079
R6964 gnd.n2179 gnd.n2178 152.079
R6965 gnd.n2147 gnd.n2146 152.079
R6966 gnd.n2901 gnd.n2900 152
R6967 gnd.n2902 gnd.n2891 152
R6968 gnd.n2904 gnd.n2903 152
R6969 gnd.n2906 gnd.n2889 152
R6970 gnd.n2908 gnd.n2907 152
R6971 gnd.n5247 gnd.n5231 152
R6972 gnd.n5239 gnd.n5232 152
R6973 gnd.n5238 gnd.n5237 152
R6974 gnd.n5236 gnd.n5233 152
R6975 gnd.n5234 gnd.t200 150.546
R6976 gnd.t38 gnd.n2189 147.661
R6977 gnd.t9 gnd.n2157 147.661
R6978 gnd.t40 gnd.n2125 147.661
R6979 gnd.t142 gnd.n2094 147.661
R6980 gnd.t138 gnd.n2062 147.661
R6981 gnd.t121 gnd.n2030 147.661
R6982 gnd.t112 gnd.n1998 147.661
R6983 gnd.t29 gnd.n1967 147.661
R6984 gnd.n5385 gnd.n3265 143.351
R6985 gnd.n2868 gnd.n2852 143.351
R6986 gnd.n6031 gnd.n2852 143.351
R6987 gnd.n5388 gnd.n5387 131.649
R6988 gnd.n6034 gnd.n6033 131.649
R6989 gnd.n2898 gnd.t251 130.484
R6990 gnd.n2907 gnd.t214 126.766
R6991 gnd.n2905 gnd.t171 126.766
R6992 gnd.n2891 gnd.t224 126.766
R6993 gnd.n2899 gnd.t288 126.766
R6994 gnd.n5235 gnd.t197 126.766
R6995 gnd.n5237 gnd.t266 126.766
R6996 gnd.n5246 gnd.t241 126.766
R6997 gnd.n5248 gnd.t282 126.766
R6998 gnd.n2206 gnd.n2205 104.615
R6999 gnd.n2205 gnd.n2183 104.615
R7000 gnd.n2198 gnd.n2183 104.615
R7001 gnd.n2198 gnd.n2197 104.615
R7002 gnd.n2197 gnd.n2187 104.615
R7003 gnd.n2190 gnd.n2187 104.615
R7004 gnd.n2174 gnd.n2173 104.615
R7005 gnd.n2173 gnd.n2151 104.615
R7006 gnd.n2166 gnd.n2151 104.615
R7007 gnd.n2166 gnd.n2165 104.615
R7008 gnd.n2165 gnd.n2155 104.615
R7009 gnd.n2158 gnd.n2155 104.615
R7010 gnd.n2142 gnd.n2141 104.615
R7011 gnd.n2141 gnd.n2119 104.615
R7012 gnd.n2134 gnd.n2119 104.615
R7013 gnd.n2134 gnd.n2133 104.615
R7014 gnd.n2133 gnd.n2123 104.615
R7015 gnd.n2126 gnd.n2123 104.615
R7016 gnd.n2111 gnd.n2110 104.615
R7017 gnd.n2110 gnd.n2088 104.615
R7018 gnd.n2103 gnd.n2088 104.615
R7019 gnd.n2103 gnd.n2102 104.615
R7020 gnd.n2102 gnd.n2092 104.615
R7021 gnd.n2095 gnd.n2092 104.615
R7022 gnd.n2079 gnd.n2078 104.615
R7023 gnd.n2078 gnd.n2056 104.615
R7024 gnd.n2071 gnd.n2056 104.615
R7025 gnd.n2071 gnd.n2070 104.615
R7026 gnd.n2070 gnd.n2060 104.615
R7027 gnd.n2063 gnd.n2060 104.615
R7028 gnd.n2047 gnd.n2046 104.615
R7029 gnd.n2046 gnd.n2024 104.615
R7030 gnd.n2039 gnd.n2024 104.615
R7031 gnd.n2039 gnd.n2038 104.615
R7032 gnd.n2038 gnd.n2028 104.615
R7033 gnd.n2031 gnd.n2028 104.615
R7034 gnd.n2015 gnd.n2014 104.615
R7035 gnd.n2014 gnd.n1992 104.615
R7036 gnd.n2007 gnd.n1992 104.615
R7037 gnd.n2007 gnd.n2006 104.615
R7038 gnd.n2006 gnd.n1996 104.615
R7039 gnd.n1999 gnd.n1996 104.615
R7040 gnd.n1984 gnd.n1983 104.615
R7041 gnd.n1983 gnd.n1961 104.615
R7042 gnd.n1976 gnd.n1961 104.615
R7043 gnd.n1976 gnd.n1975 104.615
R7044 gnd.n1975 gnd.n1965 104.615
R7045 gnd.n1968 gnd.n1965 104.615
R7046 gnd.n1356 gnd.t247 100.632
R7047 gnd.n916 gnd.t274 100.632
R7048 gnd.n7468 gnd.n7467 99.6594
R7049 gnd.n7463 gnd.n7284 99.6594
R7050 gnd.n7459 gnd.n7283 99.6594
R7051 gnd.n7455 gnd.n7282 99.6594
R7052 gnd.n7451 gnd.n7281 99.6594
R7053 gnd.n7447 gnd.n7280 99.6594
R7054 gnd.n7443 gnd.n7279 99.6594
R7055 gnd.n7439 gnd.n7278 99.6594
R7056 gnd.n7432 gnd.n7277 99.6594
R7057 gnd.n7428 gnd.n7276 99.6594
R7058 gnd.n7424 gnd.n7275 99.6594
R7059 gnd.n7420 gnd.n7274 99.6594
R7060 gnd.n7416 gnd.n7273 99.6594
R7061 gnd.n7412 gnd.n7272 99.6594
R7062 gnd.n7408 gnd.n7271 99.6594
R7063 gnd.n7404 gnd.n7270 99.6594
R7064 gnd.n7400 gnd.n7269 99.6594
R7065 gnd.n7396 gnd.n7268 99.6594
R7066 gnd.n7388 gnd.n7267 99.6594
R7067 gnd.n7386 gnd.n7266 99.6594
R7068 gnd.n7382 gnd.n7265 99.6594
R7069 gnd.n7378 gnd.n7264 99.6594
R7070 gnd.n7374 gnd.n7263 99.6594
R7071 gnd.n7370 gnd.n7262 99.6594
R7072 gnd.n7366 gnd.n7261 99.6594
R7073 gnd.n7362 gnd.n7260 99.6594
R7074 gnd.n7358 gnd.n7259 99.6594
R7075 gnd.n7354 gnd.n7258 99.6594
R7076 gnd.n7346 gnd.n7257 99.6594
R7077 gnd.n5417 gnd.n3025 99.6594
R7078 gnd.n5421 gnd.n5420 99.6594
R7079 gnd.n5428 gnd.n5427 99.6594
R7080 gnd.n5431 gnd.n5430 99.6594
R7081 gnd.n5438 gnd.n5437 99.6594
R7082 gnd.n5441 gnd.n5440 99.6594
R7083 gnd.n5448 gnd.n5447 99.6594
R7084 gnd.n5451 gnd.n5450 99.6594
R7085 gnd.n5461 gnd.n5460 99.6594
R7086 gnd.n5464 gnd.n5463 99.6594
R7087 gnd.n5471 gnd.n5470 99.6594
R7088 gnd.n5474 gnd.n5473 99.6594
R7089 gnd.n5482 gnd.n5481 99.6594
R7090 gnd.n5487 gnd.n5486 99.6594
R7091 gnd.n5494 gnd.n5493 99.6594
R7092 gnd.n5497 gnd.n5496 99.6594
R7093 gnd.n5504 gnd.n5503 99.6594
R7094 gnd.n5507 gnd.n5506 99.6594
R7095 gnd.n5516 gnd.n5515 99.6594
R7096 gnd.n5519 gnd.n5518 99.6594
R7097 gnd.n5526 gnd.n5525 99.6594
R7098 gnd.n5529 gnd.n5528 99.6594
R7099 gnd.n5536 gnd.n5535 99.6594
R7100 gnd.n5539 gnd.n5538 99.6594
R7101 gnd.n5546 gnd.n5545 99.6594
R7102 gnd.n5549 gnd.n5548 99.6594
R7103 gnd.n5557 gnd.n5556 99.6594
R7104 gnd.n5560 gnd.n5559 99.6594
R7105 gnd.n6083 gnd.n6082 99.6594
R7106 gnd.n6078 gnd.n2718 99.6594
R7107 gnd.n6074 gnd.n2717 99.6594
R7108 gnd.n6070 gnd.n2716 99.6594
R7109 gnd.n6066 gnd.n2715 99.6594
R7110 gnd.n6062 gnd.n2714 99.6594
R7111 gnd.n6058 gnd.n2713 99.6594
R7112 gnd.n6054 gnd.n2712 99.6594
R7113 gnd.n6049 gnd.n2711 99.6594
R7114 gnd.n6045 gnd.n2710 99.6594
R7115 gnd.n6041 gnd.n2709 99.6594
R7116 gnd.n6037 gnd.n2708 99.6594
R7117 gnd.n2844 gnd.n2706 99.6594
R7118 gnd.n2842 gnd.n2705 99.6594
R7119 gnd.n2838 gnd.n2704 99.6594
R7120 gnd.n2834 gnd.n2703 99.6594
R7121 gnd.n2830 gnd.n2702 99.6594
R7122 gnd.n2822 gnd.n2701 99.6594
R7123 gnd.n2820 gnd.n2700 99.6594
R7124 gnd.n2816 gnd.n2699 99.6594
R7125 gnd.n2812 gnd.n2698 99.6594
R7126 gnd.n2808 gnd.n2697 99.6594
R7127 gnd.n2804 gnd.n2696 99.6594
R7128 gnd.n2800 gnd.n2695 99.6594
R7129 gnd.n2796 gnd.n2694 99.6594
R7130 gnd.n2792 gnd.n2693 99.6594
R7131 gnd.n2788 gnd.n2692 99.6594
R7132 gnd.n2780 gnd.n2691 99.6594
R7133 gnd.n3974 gnd.n2368 99.6594
R7134 gnd.n3982 gnd.n3981 99.6594
R7135 gnd.n3985 gnd.n3984 99.6594
R7136 gnd.n3992 gnd.n3991 99.6594
R7137 gnd.n3995 gnd.n3994 99.6594
R7138 gnd.n4002 gnd.n4001 99.6594
R7139 gnd.n4005 gnd.n4004 99.6594
R7140 gnd.n4012 gnd.n4011 99.6594
R7141 gnd.n4015 gnd.n4014 99.6594
R7142 gnd.n4022 gnd.n4021 99.6594
R7143 gnd.n4025 gnd.n4024 99.6594
R7144 gnd.n4032 gnd.n4031 99.6594
R7145 gnd.n4035 gnd.n4034 99.6594
R7146 gnd.n4042 gnd.n4041 99.6594
R7147 gnd.n4045 gnd.n4044 99.6594
R7148 gnd.n4052 gnd.n4051 99.6594
R7149 gnd.n4055 gnd.n4054 99.6594
R7150 gnd.n4062 gnd.n4061 99.6594
R7151 gnd.n4065 gnd.n4064 99.6594
R7152 gnd.n4074 gnd.n4073 99.6594
R7153 gnd.n4077 gnd.n4076 99.6594
R7154 gnd.n4084 gnd.n4083 99.6594
R7155 gnd.n4087 gnd.n4086 99.6594
R7156 gnd.n4094 gnd.n4093 99.6594
R7157 gnd.n4097 gnd.n4096 99.6594
R7158 gnd.n4104 gnd.n4103 99.6594
R7159 gnd.n4107 gnd.n4106 99.6594
R7160 gnd.n4115 gnd.n4114 99.6594
R7161 gnd.n4118 gnd.n4117 99.6594
R7162 gnd.n2329 gnd.n899 99.6594
R7163 gnd.n2327 gnd.n898 99.6594
R7164 gnd.n2323 gnd.n897 99.6594
R7165 gnd.n2319 gnd.n896 99.6594
R7166 gnd.n2315 gnd.n895 99.6594
R7167 gnd.n2311 gnd.n894 99.6594
R7168 gnd.n2307 gnd.n893 99.6594
R7169 gnd.n2239 gnd.n892 99.6594
R7170 gnd.n1568 gnd.n1299 99.6594
R7171 gnd.n1325 gnd.n1306 99.6594
R7172 gnd.n1327 gnd.n1307 99.6594
R7173 gnd.n1335 gnd.n1308 99.6594
R7174 gnd.n1337 gnd.n1309 99.6594
R7175 gnd.n1345 gnd.n1310 99.6594
R7176 gnd.n1347 gnd.n1311 99.6594
R7177 gnd.n1355 gnd.n1312 99.6594
R7178 gnd.n206 gnd.n185 99.6594
R7179 gnd.n212 gnd.n186 99.6594
R7180 gnd.n216 gnd.n187 99.6594
R7181 gnd.n222 gnd.n188 99.6594
R7182 gnd.n226 gnd.n189 99.6594
R7183 gnd.n232 gnd.n190 99.6594
R7184 gnd.n235 gnd.n191 99.6594
R7185 gnd.n242 gnd.n241 99.6594
R7186 gnd.n7471 gnd.n7470 99.6594
R7187 gnd.n5079 gnd.n5078 99.6594
R7188 gnd.n5095 gnd.n5094 99.6594
R7189 gnd.n5098 gnd.n5097 99.6594
R7190 gnd.n5114 gnd.n5113 99.6594
R7191 gnd.n5117 gnd.n5116 99.6594
R7192 gnd.n5133 gnd.n5132 99.6594
R7193 gnd.n5136 gnd.n5135 99.6594
R7194 gnd.n5153 gnd.n5152 99.6594
R7195 gnd.n5156 gnd.n5155 99.6594
R7196 gnd.n2297 gnd.n879 99.6594
R7197 gnd.n2293 gnd.n880 99.6594
R7198 gnd.n2289 gnd.n881 99.6594
R7199 gnd.n2285 gnd.n882 99.6594
R7200 gnd.n2281 gnd.n883 99.6594
R7201 gnd.n2277 gnd.n884 99.6594
R7202 gnd.n2273 gnd.n885 99.6594
R7203 gnd.n2269 gnd.n886 99.6594
R7204 gnd.n2265 gnd.n887 99.6594
R7205 gnd.n2261 gnd.n888 99.6594
R7206 gnd.n2257 gnd.n889 99.6594
R7207 gnd.n2253 gnd.n890 99.6594
R7208 gnd.n2249 gnd.n891 99.6594
R7209 gnd.n1483 gnd.n1482 99.6594
R7210 gnd.n1477 gnd.n1394 99.6594
R7211 gnd.n1474 gnd.n1395 99.6594
R7212 gnd.n1470 gnd.n1396 99.6594
R7213 gnd.n1466 gnd.n1397 99.6594
R7214 gnd.n1462 gnd.n1398 99.6594
R7215 gnd.n1458 gnd.n1399 99.6594
R7216 gnd.n1454 gnd.n1400 99.6594
R7217 gnd.n1450 gnd.n1401 99.6594
R7218 gnd.n1446 gnd.n1402 99.6594
R7219 gnd.n1442 gnd.n1403 99.6594
R7220 gnd.n1438 gnd.n1404 99.6594
R7221 gnd.n1485 gnd.n1393 99.6594
R7222 gnd.n2677 gnd.n2622 99.6594
R7223 gnd.n2679 gnd.n2631 99.6594
R7224 gnd.n2681 gnd.n2680 99.6594
R7225 gnd.n2682 gnd.n2640 99.6594
R7226 gnd.n2684 gnd.n2649 99.6594
R7227 gnd.n2686 gnd.n2685 99.6594
R7228 gnd.n2687 gnd.n2658 99.6594
R7229 gnd.n2689 gnd.n2670 99.6594
R7230 gnd.n6086 gnd.n6085 99.6594
R7231 gnd.n3907 gnd.n3906 99.6594
R7232 gnd.n3904 gnd.n3843 99.6594
R7233 gnd.n3900 gnd.n3899 99.6594
R7234 gnd.n3893 gnd.n3847 99.6594
R7235 gnd.n3892 gnd.n3891 99.6594
R7236 gnd.n3885 gnd.n3853 99.6594
R7237 gnd.n3884 gnd.n3883 99.6594
R7238 gnd.n3877 gnd.n3859 99.6594
R7239 gnd.n3876 gnd.n3875 99.6594
R7240 gnd.n3906 gnd.n3905 99.6594
R7241 gnd.n3901 gnd.n3843 99.6594
R7242 gnd.n3899 gnd.n3898 99.6594
R7243 gnd.n3894 gnd.n3893 99.6594
R7244 gnd.n3891 gnd.n3890 99.6594
R7245 gnd.n3886 gnd.n3885 99.6594
R7246 gnd.n3883 gnd.n3882 99.6594
R7247 gnd.n3878 gnd.n3877 99.6594
R7248 gnd.n3875 gnd.n3874 99.6594
R7249 gnd.n6085 gnd.n2675 99.6594
R7250 gnd.n2689 gnd.n2688 99.6594
R7251 gnd.n2687 gnd.n2657 99.6594
R7252 gnd.n2686 gnd.n2650 99.6594
R7253 gnd.n2684 gnd.n2683 99.6594
R7254 gnd.n2682 gnd.n2639 99.6594
R7255 gnd.n2681 gnd.n2632 99.6594
R7256 gnd.n2679 gnd.n2678 99.6594
R7257 gnd.n2677 gnd.n2621 99.6594
R7258 gnd.n1483 gnd.n1406 99.6594
R7259 gnd.n1475 gnd.n1394 99.6594
R7260 gnd.n1471 gnd.n1395 99.6594
R7261 gnd.n1467 gnd.n1396 99.6594
R7262 gnd.n1463 gnd.n1397 99.6594
R7263 gnd.n1459 gnd.n1398 99.6594
R7264 gnd.n1455 gnd.n1399 99.6594
R7265 gnd.n1451 gnd.n1400 99.6594
R7266 gnd.n1447 gnd.n1401 99.6594
R7267 gnd.n1443 gnd.n1402 99.6594
R7268 gnd.n1439 gnd.n1403 99.6594
R7269 gnd.n1435 gnd.n1404 99.6594
R7270 gnd.n1486 gnd.n1485 99.6594
R7271 gnd.n2252 gnd.n891 99.6594
R7272 gnd.n2256 gnd.n890 99.6594
R7273 gnd.n2260 gnd.n889 99.6594
R7274 gnd.n2264 gnd.n888 99.6594
R7275 gnd.n2268 gnd.n887 99.6594
R7276 gnd.n2272 gnd.n886 99.6594
R7277 gnd.n2276 gnd.n885 99.6594
R7278 gnd.n2280 gnd.n884 99.6594
R7279 gnd.n2284 gnd.n883 99.6594
R7280 gnd.n2288 gnd.n882 99.6594
R7281 gnd.n2292 gnd.n881 99.6594
R7282 gnd.n2296 gnd.n880 99.6594
R7283 gnd.n920 gnd.n879 99.6594
R7284 gnd.n5078 gnd.n5042 99.6594
R7285 gnd.n5096 gnd.n5095 99.6594
R7286 gnd.n5097 gnd.n5033 99.6594
R7287 gnd.n5115 gnd.n5114 99.6594
R7288 gnd.n5116 gnd.n5024 99.6594
R7289 gnd.n5134 gnd.n5133 99.6594
R7290 gnd.n5135 gnd.n5015 99.6594
R7291 gnd.n5154 gnd.n5153 99.6594
R7292 gnd.n5155 gnd.n5011 99.6594
R7293 gnd.n7470 gnd.n183 99.6594
R7294 gnd.n242 gnd.n192 99.6594
R7295 gnd.n233 gnd.n191 99.6594
R7296 gnd.n225 gnd.n190 99.6594
R7297 gnd.n223 gnd.n189 99.6594
R7298 gnd.n215 gnd.n188 99.6594
R7299 gnd.n213 gnd.n187 99.6594
R7300 gnd.n205 gnd.n186 99.6594
R7301 gnd.n203 gnd.n185 99.6594
R7302 gnd.n1569 gnd.n1568 99.6594
R7303 gnd.n1328 gnd.n1306 99.6594
R7304 gnd.n1334 gnd.n1307 99.6594
R7305 gnd.n1338 gnd.n1308 99.6594
R7306 gnd.n1344 gnd.n1309 99.6594
R7307 gnd.n1348 gnd.n1310 99.6594
R7308 gnd.n1354 gnd.n1311 99.6594
R7309 gnd.n1312 gnd.n1296 99.6594
R7310 gnd.n2306 gnd.n892 99.6594
R7311 gnd.n2310 gnd.n893 99.6594
R7312 gnd.n2314 gnd.n894 99.6594
R7313 gnd.n2318 gnd.n895 99.6594
R7314 gnd.n2322 gnd.n896 99.6594
R7315 gnd.n2326 gnd.n897 99.6594
R7316 gnd.n2330 gnd.n898 99.6594
R7317 gnd.n901 gnd.n899 99.6594
R7318 gnd.n3975 gnd.n3974 99.6594
R7319 gnd.n3983 gnd.n3982 99.6594
R7320 gnd.n3984 gnd.n3966 99.6594
R7321 gnd.n3993 gnd.n3992 99.6594
R7322 gnd.n3994 gnd.n3962 99.6594
R7323 gnd.n4003 gnd.n4002 99.6594
R7324 gnd.n4004 gnd.n3958 99.6594
R7325 gnd.n4013 gnd.n4012 99.6594
R7326 gnd.n4014 gnd.n3951 99.6594
R7327 gnd.n4023 gnd.n4022 99.6594
R7328 gnd.n4024 gnd.n3947 99.6594
R7329 gnd.n4033 gnd.n4032 99.6594
R7330 gnd.n4034 gnd.n3943 99.6594
R7331 gnd.n4043 gnd.n4042 99.6594
R7332 gnd.n4044 gnd.n3939 99.6594
R7333 gnd.n4053 gnd.n4052 99.6594
R7334 gnd.n4054 gnd.n3935 99.6594
R7335 gnd.n4063 gnd.n4062 99.6594
R7336 gnd.n4064 gnd.n3931 99.6594
R7337 gnd.n4075 gnd.n4074 99.6594
R7338 gnd.n4076 gnd.n3927 99.6594
R7339 gnd.n4085 gnd.n4084 99.6594
R7340 gnd.n4086 gnd.n3923 99.6594
R7341 gnd.n4095 gnd.n4094 99.6594
R7342 gnd.n4096 gnd.n3919 99.6594
R7343 gnd.n4105 gnd.n4104 99.6594
R7344 gnd.n4106 gnd.n3915 99.6594
R7345 gnd.n4116 gnd.n4115 99.6594
R7346 gnd.n4119 gnd.n4118 99.6594
R7347 gnd.n2787 gnd.n2691 99.6594
R7348 gnd.n2791 gnd.n2692 99.6594
R7349 gnd.n2795 gnd.n2693 99.6594
R7350 gnd.n2799 gnd.n2694 99.6594
R7351 gnd.n2803 gnd.n2695 99.6594
R7352 gnd.n2807 gnd.n2696 99.6594
R7353 gnd.n2811 gnd.n2697 99.6594
R7354 gnd.n2815 gnd.n2698 99.6594
R7355 gnd.n2819 gnd.n2699 99.6594
R7356 gnd.n2823 gnd.n2700 99.6594
R7357 gnd.n2829 gnd.n2701 99.6594
R7358 gnd.n2833 gnd.n2702 99.6594
R7359 gnd.n2837 gnd.n2703 99.6594
R7360 gnd.n2841 gnd.n2704 99.6594
R7361 gnd.n2845 gnd.n2705 99.6594
R7362 gnd.n6036 gnd.n2707 99.6594
R7363 gnd.n6040 gnd.n2708 99.6594
R7364 gnd.n6044 gnd.n2709 99.6594
R7365 gnd.n6048 gnd.n2710 99.6594
R7366 gnd.n6053 gnd.n2711 99.6594
R7367 gnd.n6057 gnd.n2712 99.6594
R7368 gnd.n6061 gnd.n2713 99.6594
R7369 gnd.n6065 gnd.n2714 99.6594
R7370 gnd.n6069 gnd.n2715 99.6594
R7371 gnd.n6073 gnd.n2716 99.6594
R7372 gnd.n6077 gnd.n2717 99.6594
R7373 gnd.n2720 gnd.n2718 99.6594
R7374 gnd.n6083 gnd.n2719 99.6594
R7375 gnd.n5418 gnd.n5417 99.6594
R7376 gnd.n5420 gnd.n5409 99.6594
R7377 gnd.n5429 gnd.n5428 99.6594
R7378 gnd.n5430 gnd.n5405 99.6594
R7379 gnd.n5439 gnd.n5438 99.6594
R7380 gnd.n5440 gnd.n5401 99.6594
R7381 gnd.n5449 gnd.n5448 99.6594
R7382 gnd.n5450 gnd.n5397 99.6594
R7383 gnd.n5462 gnd.n5461 99.6594
R7384 gnd.n5463 gnd.n5393 99.6594
R7385 gnd.n5472 gnd.n5471 99.6594
R7386 gnd.n5473 gnd.n5389 99.6594
R7387 gnd.n5485 gnd.n5484 99.6594
R7388 gnd.n5486 gnd.n3259 99.6594
R7389 gnd.n5495 gnd.n5494 99.6594
R7390 gnd.n5496 gnd.n3255 99.6594
R7391 gnd.n5505 gnd.n5504 99.6594
R7392 gnd.n5506 gnd.n3251 99.6594
R7393 gnd.n5517 gnd.n5516 99.6594
R7394 gnd.n5518 gnd.n3247 99.6594
R7395 gnd.n5527 gnd.n5526 99.6594
R7396 gnd.n5528 gnd.n3243 99.6594
R7397 gnd.n5537 gnd.n5536 99.6594
R7398 gnd.n5538 gnd.n3239 99.6594
R7399 gnd.n5547 gnd.n5546 99.6594
R7400 gnd.n5548 gnd.n3235 99.6594
R7401 gnd.n5558 gnd.n5557 99.6594
R7402 gnd.n5561 gnd.n5560 99.6594
R7403 gnd.n7353 gnd.n7257 99.6594
R7404 gnd.n7357 gnd.n7258 99.6594
R7405 gnd.n7361 gnd.n7259 99.6594
R7406 gnd.n7365 gnd.n7260 99.6594
R7407 gnd.n7369 gnd.n7261 99.6594
R7408 gnd.n7373 gnd.n7262 99.6594
R7409 gnd.n7377 gnd.n7263 99.6594
R7410 gnd.n7381 gnd.n7264 99.6594
R7411 gnd.n7385 gnd.n7265 99.6594
R7412 gnd.n7389 gnd.n7266 99.6594
R7413 gnd.n7395 gnd.n7267 99.6594
R7414 gnd.n7399 gnd.n7268 99.6594
R7415 gnd.n7403 gnd.n7269 99.6594
R7416 gnd.n7407 gnd.n7270 99.6594
R7417 gnd.n7411 gnd.n7271 99.6594
R7418 gnd.n7415 gnd.n7272 99.6594
R7419 gnd.n7419 gnd.n7273 99.6594
R7420 gnd.n7423 gnd.n7274 99.6594
R7421 gnd.n7427 gnd.n7275 99.6594
R7422 gnd.n7431 gnd.n7276 99.6594
R7423 gnd.n7438 gnd.n7277 99.6594
R7424 gnd.n7442 gnd.n7278 99.6594
R7425 gnd.n7446 gnd.n7279 99.6594
R7426 gnd.n7450 gnd.n7280 99.6594
R7427 gnd.n7454 gnd.n7281 99.6594
R7428 gnd.n7458 gnd.n7282 99.6594
R7429 gnd.n7462 gnd.n7283 99.6594
R7430 gnd.n7286 gnd.n7284 99.6594
R7431 gnd.n7468 gnd.n7285 99.6594
R7432 gnd.n6148 gnd.n6147 99.6594
R7433 gnd.n2608 gnd.n2588 99.6594
R7434 gnd.n2610 gnd.n2589 99.6594
R7435 gnd.n2614 gnd.n2590 99.6594
R7436 gnd.n2616 gnd.n2591 99.6594
R7437 gnd.n2626 gnd.n2592 99.6594
R7438 gnd.n2628 gnd.n2593 99.6594
R7439 gnd.n2636 gnd.n2594 99.6594
R7440 gnd.n2644 gnd.n2595 99.6594
R7441 gnd.n2646 gnd.n2596 99.6594
R7442 gnd.n2654 gnd.n2597 99.6594
R7443 gnd.n2662 gnd.n2598 99.6594
R7444 gnd.n2667 gnd.n2600 99.6594
R7445 gnd.n6150 gnd.n2585 99.6594
R7446 gnd.n6148 gnd.n2603 99.6594
R7447 gnd.n2609 gnd.n2588 99.6594
R7448 gnd.n2613 gnd.n2589 99.6594
R7449 gnd.n2615 gnd.n2590 99.6594
R7450 gnd.n2625 gnd.n2591 99.6594
R7451 gnd.n2627 gnd.n2592 99.6594
R7452 gnd.n2635 gnd.n2593 99.6594
R7453 gnd.n2643 gnd.n2594 99.6594
R7454 gnd.n2645 gnd.n2595 99.6594
R7455 gnd.n2653 gnd.n2596 99.6594
R7456 gnd.n2661 gnd.n2597 99.6594
R7457 gnd.n2663 gnd.n2598 99.6594
R7458 gnd.n2600 gnd.n2599 99.6594
R7459 gnd.n6151 gnd.n6150 99.6594
R7460 gnd.n5059 gnd.n5054 99.6594
R7461 gnd.n5063 gnd.n5061 99.6594
R7462 gnd.n5070 gnd.n5050 99.6594
R7463 gnd.n5074 gnd.n5072 99.6594
R7464 gnd.n5085 gnd.n5047 99.6594
R7465 gnd.n5089 gnd.n5087 99.6594
R7466 gnd.n5104 gnd.n5038 99.6594
R7467 gnd.n5108 gnd.n5106 99.6594
R7468 gnd.n5123 gnd.n5029 99.6594
R7469 gnd.n5127 gnd.n5125 99.6594
R7470 gnd.n5142 gnd.n5020 99.6594
R7471 gnd.n5145 gnd.n5144 99.6594
R7472 gnd.n5163 gnd.n5162 99.6594
R7473 gnd.n5166 gnd.n5165 99.6594
R7474 gnd.n5144 gnd.n5143 99.6594
R7475 gnd.n5126 gnd.n5020 99.6594
R7476 gnd.n5125 gnd.n5124 99.6594
R7477 gnd.n5107 gnd.n5029 99.6594
R7478 gnd.n5106 gnd.n5105 99.6594
R7479 gnd.n5088 gnd.n5038 99.6594
R7480 gnd.n5087 gnd.n5086 99.6594
R7481 gnd.n5073 gnd.n5047 99.6594
R7482 gnd.n5072 gnd.n5071 99.6594
R7483 gnd.n5062 gnd.n5050 99.6594
R7484 gnd.n5061 gnd.n5060 99.6594
R7485 gnd.n5054 gnd.n2999 99.6594
R7486 gnd.n5167 gnd.n5166 99.6594
R7487 gnd.n5164 gnd.n5163 99.6594
R7488 gnd.n2664 gnd.t240 98.63
R7489 gnd.n5012 gnd.t265 98.63
R7490 gnd.n2671 gnd.t286 98.63
R7491 gnd.n5456 gnd.t262 98.63
R7492 gnd.n5508 gnd.t250 98.63
R7493 gnd.n3231 gnd.t196 98.63
R7494 gnd.n7348 gnd.t176 98.63
R7495 gnd.n7327 gnd.t191 98.63
R7496 gnd.n7434 gnd.t255 98.63
R7497 gnd.n180 gnd.t277 98.63
R7498 gnd.n3955 gnd.t223 98.63
R7499 gnd.n4066 gnd.t205 98.63
R7500 gnd.n3911 gnd.t233 98.63
R7501 gnd.n3871 gnd.t189 98.63
R7502 gnd.n2741 gnd.t270 98.63
R7503 gnd.n2782 gnd.t212 98.63
R7504 gnd.n2761 gnd.t235 98.63
R7505 gnd.n5002 gnd.t219 98.63
R7506 gnd.n3609 gnd.t209 92.8196
R7507 gnd.n3300 gnd.t229 92.8196
R7508 gnd.n5965 gnd.t259 92.8118
R7509 gnd.n5250 gnd.t280 92.8118
R7510 gnd.n2898 gnd.n2897 81.8399
R7511 gnd.n1357 gnd.t246 74.8376
R7512 gnd.n917 gnd.t275 74.8376
R7513 gnd.n3610 gnd.t208 72.8438
R7514 gnd.n3301 gnd.t230 72.8438
R7515 gnd.n2899 gnd.n2892 72.8411
R7516 gnd.n2905 gnd.n2890 72.8411
R7517 gnd.n5246 gnd.n5245 72.8411
R7518 gnd.n2665 gnd.t239 72.836
R7519 gnd.n5966 gnd.t258 72.836
R7520 gnd.n5251 gnd.t281 72.836
R7521 gnd.n5013 gnd.t264 72.836
R7522 gnd.n2672 gnd.t287 72.836
R7523 gnd.n5457 gnd.t261 72.836
R7524 gnd.n5509 gnd.t249 72.836
R7525 gnd.n3232 gnd.t195 72.836
R7526 gnd.n7349 gnd.t177 72.836
R7527 gnd.n7328 gnd.t192 72.836
R7528 gnd.n7435 gnd.t256 72.836
R7529 gnd.n181 gnd.t278 72.836
R7530 gnd.n3956 gnd.t222 72.836
R7531 gnd.n4067 gnd.t204 72.836
R7532 gnd.n3912 gnd.t232 72.836
R7533 gnd.n3872 gnd.t188 72.836
R7534 gnd.n2742 gnd.t271 72.836
R7535 gnd.n2783 gnd.t213 72.836
R7536 gnd.n2762 gnd.t236 72.836
R7537 gnd.n5003 gnd.t220 72.836
R7538 gnd.n5311 gnd.n3268 71.676
R7539 gnd.n5307 gnd.n3269 71.676
R7540 gnd.n5303 gnd.n3270 71.676
R7541 gnd.n5299 gnd.n3271 71.676
R7542 gnd.n5295 gnd.n3272 71.676
R7543 gnd.n5291 gnd.n3273 71.676
R7544 gnd.n5287 gnd.n3274 71.676
R7545 gnd.n5283 gnd.n3275 71.676
R7546 gnd.n5279 gnd.n3276 71.676
R7547 gnd.n5275 gnd.n3277 71.676
R7548 gnd.n5271 gnd.n3278 71.676
R7549 gnd.n5267 gnd.n3279 71.676
R7550 gnd.n5263 gnd.n3280 71.676
R7551 gnd.n5259 gnd.n3281 71.676
R7552 gnd.n5254 gnd.n3282 71.676
R7553 gnd.n3283 gnd.n3266 71.676
R7554 gnd.n5383 gnd.n3265 71.676
R7555 gnd.n5381 gnd.n5380 71.676
R7556 gnd.n5375 gnd.n3298 71.676
R7557 gnd.n5371 gnd.n3297 71.676
R7558 gnd.n5367 gnd.n3296 71.676
R7559 gnd.n5363 gnd.n3295 71.676
R7560 gnd.n5359 gnd.n3294 71.676
R7561 gnd.n5355 gnd.n3293 71.676
R7562 gnd.n5351 gnd.n3292 71.676
R7563 gnd.n5347 gnd.n3291 71.676
R7564 gnd.n5343 gnd.n3290 71.676
R7565 gnd.n5339 gnd.n3289 71.676
R7566 gnd.n5335 gnd.n3288 71.676
R7567 gnd.n5331 gnd.n3287 71.676
R7568 gnd.n5327 gnd.n3286 71.676
R7569 gnd.n5323 gnd.n3285 71.676
R7570 gnd.n5319 gnd.n3284 71.676
R7571 gnd.n6029 gnd.n6028 71.676
R7572 gnd.n6023 gnd.n2854 71.676
R7573 gnd.n6020 gnd.n2855 71.676
R7574 gnd.n6016 gnd.n2856 71.676
R7575 gnd.n6012 gnd.n2857 71.676
R7576 gnd.n6008 gnd.n2858 71.676
R7577 gnd.n6004 gnd.n2859 71.676
R7578 gnd.n6000 gnd.n2860 71.676
R7579 gnd.n5996 gnd.n2861 71.676
R7580 gnd.n5992 gnd.n2862 71.676
R7581 gnd.n5988 gnd.n2863 71.676
R7582 gnd.n5984 gnd.n2864 71.676
R7583 gnd.n5980 gnd.n2865 71.676
R7584 gnd.n5976 gnd.n2866 71.676
R7585 gnd.n5972 gnd.n2867 71.676
R7586 gnd.n5968 gnd.n2868 71.676
R7587 gnd.n2869 gnd.n2853 71.676
R7588 gnd.n3613 gnd.n2870 71.676
R7589 gnd.n3618 gnd.n2871 71.676
R7590 gnd.n3622 gnd.n2872 71.676
R7591 gnd.n3626 gnd.n2873 71.676
R7592 gnd.n3630 gnd.n2874 71.676
R7593 gnd.n3634 gnd.n2875 71.676
R7594 gnd.n3638 gnd.n2876 71.676
R7595 gnd.n3642 gnd.n2877 71.676
R7596 gnd.n3646 gnd.n2878 71.676
R7597 gnd.n3650 gnd.n2879 71.676
R7598 gnd.n3654 gnd.n2880 71.676
R7599 gnd.n3658 gnd.n2881 71.676
R7600 gnd.n3662 gnd.n2882 71.676
R7601 gnd.n3666 gnd.n2883 71.676
R7602 gnd.n3670 gnd.n2884 71.676
R7603 gnd.n6029 gnd.n2887 71.676
R7604 gnd.n6021 gnd.n2854 71.676
R7605 gnd.n6017 gnd.n2855 71.676
R7606 gnd.n6013 gnd.n2856 71.676
R7607 gnd.n6009 gnd.n2857 71.676
R7608 gnd.n6005 gnd.n2858 71.676
R7609 gnd.n6001 gnd.n2859 71.676
R7610 gnd.n5997 gnd.n2860 71.676
R7611 gnd.n5993 gnd.n2861 71.676
R7612 gnd.n5989 gnd.n2862 71.676
R7613 gnd.n5985 gnd.n2863 71.676
R7614 gnd.n5981 gnd.n2864 71.676
R7615 gnd.n5977 gnd.n2865 71.676
R7616 gnd.n5973 gnd.n2866 71.676
R7617 gnd.n5969 gnd.n2867 71.676
R7618 gnd.n6032 gnd.n6031 71.676
R7619 gnd.n3612 gnd.n2869 71.676
R7620 gnd.n3617 gnd.n2870 71.676
R7621 gnd.n3621 gnd.n2871 71.676
R7622 gnd.n3625 gnd.n2872 71.676
R7623 gnd.n3629 gnd.n2873 71.676
R7624 gnd.n3633 gnd.n2874 71.676
R7625 gnd.n3637 gnd.n2875 71.676
R7626 gnd.n3641 gnd.n2876 71.676
R7627 gnd.n3645 gnd.n2877 71.676
R7628 gnd.n3649 gnd.n2878 71.676
R7629 gnd.n3653 gnd.n2879 71.676
R7630 gnd.n3657 gnd.n2880 71.676
R7631 gnd.n3661 gnd.n2881 71.676
R7632 gnd.n3665 gnd.n2882 71.676
R7633 gnd.n3669 gnd.n2883 71.676
R7634 gnd.n3673 gnd.n2884 71.676
R7635 gnd.n5322 gnd.n3284 71.676
R7636 gnd.n5326 gnd.n3285 71.676
R7637 gnd.n5330 gnd.n3286 71.676
R7638 gnd.n5334 gnd.n3287 71.676
R7639 gnd.n5338 gnd.n3288 71.676
R7640 gnd.n5342 gnd.n3289 71.676
R7641 gnd.n5346 gnd.n3290 71.676
R7642 gnd.n5350 gnd.n3291 71.676
R7643 gnd.n5354 gnd.n3292 71.676
R7644 gnd.n5358 gnd.n3293 71.676
R7645 gnd.n5362 gnd.n3294 71.676
R7646 gnd.n5366 gnd.n3295 71.676
R7647 gnd.n5370 gnd.n3296 71.676
R7648 gnd.n5374 gnd.n3297 71.676
R7649 gnd.n3299 gnd.n3298 71.676
R7650 gnd.n5382 gnd.n5381 71.676
R7651 gnd.n5386 gnd.n5385 71.676
R7652 gnd.n5253 gnd.n3283 71.676
R7653 gnd.n5258 gnd.n3282 71.676
R7654 gnd.n5262 gnd.n3281 71.676
R7655 gnd.n5266 gnd.n3280 71.676
R7656 gnd.n5270 gnd.n3279 71.676
R7657 gnd.n5274 gnd.n3278 71.676
R7658 gnd.n5278 gnd.n3277 71.676
R7659 gnd.n5282 gnd.n3276 71.676
R7660 gnd.n5286 gnd.n3275 71.676
R7661 gnd.n5290 gnd.n3274 71.676
R7662 gnd.n5294 gnd.n3273 71.676
R7663 gnd.n5298 gnd.n3272 71.676
R7664 gnd.n5302 gnd.n3271 71.676
R7665 gnd.n5306 gnd.n3270 71.676
R7666 gnd.n5310 gnd.n3269 71.676
R7667 gnd.n3307 gnd.n3268 71.676
R7668 gnd.n8 gnd.t135 69.1507
R7669 gnd.n14 gnd.t313 68.4792
R7670 gnd.n13 gnd.t311 68.4792
R7671 gnd.n12 gnd.t116 68.4792
R7672 gnd.n11 gnd.t78 68.4792
R7673 gnd.n10 gnd.t118 68.4792
R7674 gnd.n9 gnd.t90 68.4792
R7675 gnd.n8 gnd.t64 68.4792
R7676 gnd.n1484 gnd.n1388 64.369
R7677 gnd.n6322 gnd.n2339 59.5891
R7678 gnd.n7233 gnd.n7232 59.5891
R7679 gnd.n3615 gnd.n3610 59.5399
R7680 gnd.n5377 gnd.n3301 59.5399
R7681 gnd.n5967 gnd.n5966 59.5399
R7682 gnd.n5256 gnd.n5251 59.5399
R7683 gnd.n5964 gnd.n2908 59.1804
R7684 gnd.n2338 gnd.n877 57.3586
R7685 gnd.n1143 gnd.t55 56.407
R7686 gnd.n1108 gnd.t129 56.407
R7687 gnd.n1119 gnd.t146 56.407
R7688 gnd.n1131 gnd.t307 56.407
R7689 gnd.n52 gnd.t157 56.407
R7690 gnd.n17 gnd.t124 56.407
R7691 gnd.n28 gnd.t82 56.407
R7692 gnd.n40 gnd.t122 56.407
R7693 gnd.n1152 gnd.t319 55.8337
R7694 gnd.n1117 gnd.t148 55.8337
R7695 gnd.n1128 gnd.t161 55.8337
R7696 gnd.n1140 gnd.t127 55.8337
R7697 gnd.n61 gnd.t1 55.8337
R7698 gnd.n26 gnd.t22 55.8337
R7699 gnd.n37 gnd.t133 55.8337
R7700 gnd.n49 gnd.t301 55.8337
R7701 gnd.n2896 gnd.n2895 54.358
R7702 gnd.n5243 gnd.n5242 54.358
R7703 gnd.n1143 gnd.n1142 53.0052
R7704 gnd.n1145 gnd.n1144 53.0052
R7705 gnd.n1147 gnd.n1146 53.0052
R7706 gnd.n1149 gnd.n1148 53.0052
R7707 gnd.n1151 gnd.n1150 53.0052
R7708 gnd.n1108 gnd.n1107 53.0052
R7709 gnd.n1110 gnd.n1109 53.0052
R7710 gnd.n1112 gnd.n1111 53.0052
R7711 gnd.n1114 gnd.n1113 53.0052
R7712 gnd.n1116 gnd.n1115 53.0052
R7713 gnd.n1119 gnd.n1118 53.0052
R7714 gnd.n1121 gnd.n1120 53.0052
R7715 gnd.n1123 gnd.n1122 53.0052
R7716 gnd.n1125 gnd.n1124 53.0052
R7717 gnd.n1127 gnd.n1126 53.0052
R7718 gnd.n1131 gnd.n1130 53.0052
R7719 gnd.n1133 gnd.n1132 53.0052
R7720 gnd.n1135 gnd.n1134 53.0052
R7721 gnd.n1137 gnd.n1136 53.0052
R7722 gnd.n1139 gnd.n1138 53.0052
R7723 gnd.n60 gnd.n59 53.0052
R7724 gnd.n58 gnd.n57 53.0052
R7725 gnd.n56 gnd.n55 53.0052
R7726 gnd.n54 gnd.n53 53.0052
R7727 gnd.n52 gnd.n51 53.0052
R7728 gnd.n25 gnd.n24 53.0052
R7729 gnd.n23 gnd.n22 53.0052
R7730 gnd.n21 gnd.n20 53.0052
R7731 gnd.n19 gnd.n18 53.0052
R7732 gnd.n17 gnd.n16 53.0052
R7733 gnd.n36 gnd.n35 53.0052
R7734 gnd.n34 gnd.n33 53.0052
R7735 gnd.n32 gnd.n31 53.0052
R7736 gnd.n30 gnd.n29 53.0052
R7737 gnd.n28 gnd.n27 53.0052
R7738 gnd.n48 gnd.n47 53.0052
R7739 gnd.n46 gnd.n45 53.0052
R7740 gnd.n44 gnd.n43 53.0052
R7741 gnd.n42 gnd.n41 53.0052
R7742 gnd.n40 gnd.n39 53.0052
R7743 gnd.n5234 gnd.n5233 52.4801
R7744 gnd.n2190 gnd.t38 52.3082
R7745 gnd.n2158 gnd.t9 52.3082
R7746 gnd.n2126 gnd.t40 52.3082
R7747 gnd.n2095 gnd.t142 52.3082
R7748 gnd.n2063 gnd.t138 52.3082
R7749 gnd.n2031 gnd.t121 52.3082
R7750 gnd.n1999 gnd.t112 52.3082
R7751 gnd.n1968 gnd.t29 52.3082
R7752 gnd.n2020 gnd.n1988 51.4173
R7753 gnd.n2084 gnd.n2083 50.455
R7754 gnd.n2052 gnd.n2051 50.455
R7755 gnd.n2020 gnd.n2019 50.455
R7756 gnd.n1431 gnd.n1430 45.1884
R7757 gnd.n943 gnd.n942 45.1884
R7758 gnd.n5314 gnd.n5249 44.3322
R7759 gnd.n2899 gnd.n2898 44.3189
R7760 gnd.n6492 gnd.n705 43.8952
R7761 gnd.n6492 gnd.n6491 43.8952
R7762 gnd.n6491 gnd.n6490 43.8952
R7763 gnd.n6490 gnd.n710 43.8952
R7764 gnd.n6484 gnd.n710 43.8952
R7765 gnd.n6484 gnd.n6483 43.8952
R7766 gnd.n6483 gnd.n6482 43.8952
R7767 gnd.n6482 gnd.n718 43.8952
R7768 gnd.n6476 gnd.n718 43.8952
R7769 gnd.n6476 gnd.n6475 43.8952
R7770 gnd.n6475 gnd.n6474 43.8952
R7771 gnd.n6474 gnd.n726 43.8952
R7772 gnd.n6468 gnd.n726 43.8952
R7773 gnd.n6468 gnd.n6467 43.8952
R7774 gnd.n6467 gnd.n6466 43.8952
R7775 gnd.n6466 gnd.n734 43.8952
R7776 gnd.n6460 gnd.n734 43.8952
R7777 gnd.n6460 gnd.n6459 43.8952
R7778 gnd.n6459 gnd.n6458 43.8952
R7779 gnd.n6458 gnd.n742 43.8952
R7780 gnd.n6452 gnd.n742 43.8952
R7781 gnd.n6452 gnd.n6451 43.8952
R7782 gnd.n6451 gnd.n6450 43.8952
R7783 gnd.n6450 gnd.n750 43.8952
R7784 gnd.n6444 gnd.n750 43.8952
R7785 gnd.n6444 gnd.n6443 43.8952
R7786 gnd.n6443 gnd.n6442 43.8952
R7787 gnd.n6442 gnd.n758 43.8952
R7788 gnd.n6436 gnd.n758 43.8952
R7789 gnd.n6436 gnd.n6435 43.8952
R7790 gnd.n6435 gnd.n6434 43.8952
R7791 gnd.n6434 gnd.n766 43.8952
R7792 gnd.n6428 gnd.n766 43.8952
R7793 gnd.n6428 gnd.n6427 43.8952
R7794 gnd.n6427 gnd.n6426 43.8952
R7795 gnd.n6426 gnd.n774 43.8952
R7796 gnd.n6420 gnd.n774 43.8952
R7797 gnd.n6420 gnd.n6419 43.8952
R7798 gnd.n6419 gnd.n6418 43.8952
R7799 gnd.n6418 gnd.n782 43.8952
R7800 gnd.n6412 gnd.n782 43.8952
R7801 gnd.n6412 gnd.n6411 43.8952
R7802 gnd.n6411 gnd.n6410 43.8952
R7803 gnd.n6410 gnd.n790 43.8952
R7804 gnd.n6404 gnd.n790 43.8952
R7805 gnd.n6404 gnd.n6403 43.8952
R7806 gnd.n6403 gnd.n6402 43.8952
R7807 gnd.n6402 gnd.n798 43.8952
R7808 gnd.n6396 gnd.n798 43.8952
R7809 gnd.n6396 gnd.n6395 43.8952
R7810 gnd.n6395 gnd.n6394 43.8952
R7811 gnd.n6394 gnd.n806 43.8952
R7812 gnd.n6388 gnd.n806 43.8952
R7813 gnd.n6388 gnd.n6387 43.8952
R7814 gnd.n6387 gnd.n6386 43.8952
R7815 gnd.n6386 gnd.n814 43.8952
R7816 gnd.n6380 gnd.n814 43.8952
R7817 gnd.n6380 gnd.n6379 43.8952
R7818 gnd.n6379 gnd.n6378 43.8952
R7819 gnd.n6378 gnd.n822 43.8952
R7820 gnd.n6372 gnd.n822 43.8952
R7821 gnd.n6372 gnd.n6371 43.8952
R7822 gnd.n6371 gnd.n6370 43.8952
R7823 gnd.n6370 gnd.n830 43.8952
R7824 gnd.n6364 gnd.n830 43.8952
R7825 gnd.n6364 gnd.n6363 43.8952
R7826 gnd.n6363 gnd.n6362 43.8952
R7827 gnd.n6362 gnd.n838 43.8952
R7828 gnd.n6356 gnd.n838 43.8952
R7829 gnd.n6356 gnd.n6355 43.8952
R7830 gnd.n6355 gnd.n6354 43.8952
R7831 gnd.n6354 gnd.n846 43.8952
R7832 gnd.n6348 gnd.n846 43.8952
R7833 gnd.n6348 gnd.n6347 43.8952
R7834 gnd.n6347 gnd.n6346 43.8952
R7835 gnd.n6346 gnd.n854 43.8952
R7836 gnd.n6340 gnd.n854 43.8952
R7837 gnd.n6340 gnd.n6339 43.8952
R7838 gnd.n6339 gnd.n6338 43.8952
R7839 gnd.n6338 gnd.n862 43.8952
R7840 gnd.n6332 gnd.n862 43.8952
R7841 gnd.n6332 gnd.n6331 43.8952
R7842 gnd.n6331 gnd.n6330 43.8952
R7843 gnd.n2666 gnd.n2665 42.2793
R7844 gnd.n5158 gnd.n5013 42.2793
R7845 gnd.n1432 gnd.n1431 42.2793
R7846 gnd.n944 gnd.n943 42.2793
R7847 gnd.n1358 gnd.n1357 42.2793
R7848 gnd.n2305 gnd.n917 42.2793
R7849 gnd.n6088 gnd.n2672 42.2793
R7850 gnd.n5458 gnd.n5457 42.2793
R7851 gnd.n5510 gnd.n5509 42.2793
R7852 gnd.n3233 gnd.n3232 42.2793
R7853 gnd.n7352 gnd.n7349 42.2793
R7854 gnd.n7394 gnd.n7328 42.2793
R7855 gnd.n7436 gnd.n7435 42.2793
R7856 gnd.n182 gnd.n181 42.2793
R7857 gnd.n3957 gnd.n3956 42.2793
R7858 gnd.n4068 gnd.n4067 42.2793
R7859 gnd.n3913 gnd.n3912 42.2793
R7860 gnd.n3873 gnd.n3872 42.2793
R7861 gnd.n6051 gnd.n2742 42.2793
R7862 gnd.n2786 gnd.n2783 42.2793
R7863 gnd.n2828 gnd.n2762 42.2793
R7864 gnd.n5004 gnd.n5003 42.2793
R7865 gnd.n2897 gnd.n2896 41.6274
R7866 gnd.n5244 gnd.n5243 41.6274
R7867 gnd.n2906 gnd.n2905 40.8975
R7868 gnd.n5247 gnd.n5246 40.8975
R7869 gnd.n2905 gnd.n2904 35.055
R7870 gnd.n2900 gnd.n2899 35.055
R7871 gnd.n5236 gnd.n5235 35.055
R7872 gnd.n5246 gnd.n5232 35.055
R7873 gnd.n1494 gnd.n1388 31.8661
R7874 gnd.n1494 gnd.n1493 31.8661
R7875 gnd.n1502 gnd.n1377 31.8661
R7876 gnd.n1510 gnd.n1377 31.8661
R7877 gnd.n1510 gnd.n1371 31.8661
R7878 gnd.n1518 gnd.n1371 31.8661
R7879 gnd.n1518 gnd.n1364 31.8661
R7880 gnd.n1556 gnd.n1364 31.8661
R7881 gnd.n1566 gnd.n1297 31.8661
R7882 gnd.n6322 gnd.n6321 31.8661
R7883 gnd.n6321 gnd.n6320 31.8661
R7884 gnd.n6320 gnd.n2340 31.8661
R7885 gnd.n6314 gnd.n2340 31.8661
R7886 gnd.n6314 gnd.n6313 31.8661
R7887 gnd.n6313 gnd.n6312 31.8661
R7888 gnd.n6312 gnd.n2347 31.8661
R7889 gnd.n6306 gnd.n2347 31.8661
R7890 gnd.n6306 gnd.n6305 31.8661
R7891 gnd.n6305 gnd.n6304 31.8661
R7892 gnd.n6304 gnd.n2355 31.8661
R7893 gnd.n6298 gnd.n6297 31.8661
R7894 gnd.n2676 gnd.n2574 31.8661
R7895 gnd.n4364 gnd.n2690 31.8661
R7896 gnd.n4364 gnd.n2587 31.8661
R7897 gnd.n4373 gnd.n2601 31.8661
R7898 gnd.n5858 gnd.n3002 31.8661
R7899 gnd.n5852 gnd.n5851 31.8661
R7900 gnd.n5851 gnd.n5850 31.8661
R7901 gnd.n5844 gnd.n3020 31.8661
R7902 gnd.n184 gnd.n171 31.8661
R7903 gnd.n7256 gnd.n243 31.8661
R7904 gnd.n7250 gnd.n243 31.8661
R7905 gnd.n7250 gnd.n7249 31.8661
R7906 gnd.n7249 gnd.n7248 31.8661
R7907 gnd.n7248 gnd.n252 31.8661
R7908 gnd.n7242 gnd.n252 31.8661
R7909 gnd.n7242 gnd.n7241 31.8661
R7910 gnd.n7241 gnd.n7240 31.8661
R7911 gnd.n7240 gnd.n260 31.8661
R7912 gnd.n7234 gnd.n260 31.8661
R7913 gnd.n7234 gnd.n7233 31.8661
R7914 gnd.n5320 gnd.n3302 30.1273
R7915 gnd.n4498 gnd.n3672 30.1273
R7916 gnd.n6330 gnd.n870 26.3373
R7917 gnd.n2665 gnd.n2664 25.7944
R7918 gnd.n5013 gnd.n5012 25.7944
R7919 gnd.n1357 gnd.n1356 25.7944
R7920 gnd.n917 gnd.n916 25.7944
R7921 gnd.n2672 gnd.n2671 25.7944
R7922 gnd.n5457 gnd.n5456 25.7944
R7923 gnd.n5509 gnd.n5508 25.7944
R7924 gnd.n3232 gnd.n3231 25.7944
R7925 gnd.n7349 gnd.n7348 25.7944
R7926 gnd.n7328 gnd.n7327 25.7944
R7927 gnd.n7435 gnd.n7434 25.7944
R7928 gnd.n181 gnd.n180 25.7944
R7929 gnd.n3956 gnd.n3955 25.7944
R7930 gnd.n4067 gnd.n4066 25.7944
R7931 gnd.n3912 gnd.n3911 25.7944
R7932 gnd.n3872 gnd.n3871 25.7944
R7933 gnd.n2742 gnd.n2741 25.7944
R7934 gnd.n2783 gnd.n2782 25.7944
R7935 gnd.n2762 gnd.n2761 25.7944
R7936 gnd.n5003 gnd.n5002 25.7944
R7937 gnd.n1578 gnd.n1298 24.8557
R7938 gnd.n1588 gnd.n1281 24.8557
R7939 gnd.n1284 gnd.n1272 24.8557
R7940 gnd.n1609 gnd.n1273 24.8557
R7941 gnd.n1619 gnd.n1253 24.8557
R7942 gnd.n1629 gnd.n1628 24.8557
R7943 gnd.n1239 gnd.n1237 24.8557
R7944 gnd.n1660 gnd.n1659 24.8557
R7945 gnd.n1675 gnd.n1222 24.8557
R7946 gnd.n1729 gnd.n1161 24.8557
R7947 gnd.n1685 gnd.n1162 24.8557
R7948 gnd.n1722 gnd.n1173 24.8557
R7949 gnd.n1211 gnd.n1210 24.8557
R7950 gnd.n1716 gnd.n1715 24.8557
R7951 gnd.n1197 gnd.n1184 24.8557
R7952 gnd.n1755 gnd.n1754 24.8557
R7953 gnd.n1765 gnd.n1093 24.8557
R7954 gnd.n1777 gnd.n1085 24.8557
R7955 gnd.n1776 gnd.n1073 24.8557
R7956 gnd.n1795 gnd.n1794 24.8557
R7957 gnd.n1805 gnd.n1066 24.8557
R7958 gnd.n1816 gnd.n1054 24.8557
R7959 gnd.n1842 gnd.n1841 24.8557
R7960 gnd.n1852 gnd.n1040 24.8557
R7961 gnd.n1864 gnd.n1032 24.8557
R7962 gnd.n1882 gnd.n1881 24.8557
R7963 gnd.n1023 gnd.n1012 24.8557
R7964 gnd.n1903 gnd.n1000 24.8557
R7965 gnd.n1931 gnd.n1930 24.8557
R7966 gnd.n1942 gnd.n985 24.8557
R7967 gnd.n1953 gnd.n978 24.8557
R7968 gnd.n1952 gnd.n966 24.8557
R7969 gnd.n2225 gnd.n2224 24.8557
R7970 gnd.n2247 gnd.n951 24.8557
R7971 gnd.n1599 gnd.t28 23.2624
R7972 gnd.n1300 gnd.t245 22.6251
R7973 gnd.n2363 gnd.n2355 21.6691
R7974 gnd.n7469 gnd.n7256 21.6691
R7975 gnd.t141 gnd.n1305 21.3504
R7976 gnd.n6297 gnd.n6296 21.0318
R7977 gnd.n4166 gnd.n2366 21.0318
R7978 gnd.n4160 gnd.n2377 21.0318
R7979 gnd.n6284 gnd.n2386 21.0318
R7980 gnd.n4154 gnd.n2389 21.0318
R7981 gnd.n6278 gnd.n2397 21.0318
R7982 gnd.n6272 gnd.n2407 21.0318
R7983 gnd.n4142 gnd.n2410 21.0318
R7984 gnd.n6266 gnd.n2418 21.0318
R7985 gnd.n4197 gnd.n2421 21.0318
R7986 gnd.n4205 gnd.n2430 21.0318
R7987 gnd.n6254 gnd.n2438 21.0318
R7988 gnd.n6248 gnd.n2448 21.0318
R7989 gnd.n4220 gnd.n2451 21.0318
R7990 gnd.n6241 gnd.n2457 21.0318
R7991 gnd.n4264 gnd.n2460 21.0318
R7992 gnd.n4227 gnd.n2469 21.0318
R7993 gnd.n6228 gnd.n2474 21.0318
R7994 gnd.n4242 gnd.n4241 21.0318
R7995 gnd.n6222 gnd.n2483 21.0318
R7996 gnd.n6215 gnd.n2491 21.0318
R7997 gnd.n4283 gnd.n2494 21.0318
R7998 gnd.n4291 gnd.n2503 21.0318
R7999 gnd.n6203 gnd.n2511 21.0318
R8000 gnd.n4332 gnd.n4331 21.0318
R8001 gnd.n6197 gnd.n2520 21.0318
R8002 gnd.n6191 gnd.n2531 21.0318
R8003 gnd.n4303 gnd.n2534 21.0318
R8004 gnd.n4308 gnd.n2543 21.0318
R8005 gnd.n6179 gnd.n2551 21.0318
R8006 gnd.n4314 gnd.n2554 21.0318
R8007 gnd.n6173 gnd.n2561 21.0318
R8008 gnd.n6167 gnd.n2571 21.0318
R8009 gnd.n5843 gnd.n3023 21.0318
R8010 gnd.n5837 gnd.n3035 21.0318
R8011 gnd.n5572 gnd.n3044 21.0318
R8012 gnd.n5831 gnd.n3047 21.0318
R8013 gnd.n5580 gnd.n3055 21.0318
R8014 gnd.n5600 gnd.n3064 21.0318
R8015 gnd.n5819 gnd.n3067 21.0318
R8016 gnd.n5813 gnd.n3078 21.0318
R8017 gnd.n5645 gnd.n5644 21.0318
R8018 gnd.n5807 gnd.n3087 21.0318
R8019 gnd.n5652 gnd.n3095 21.0318
R8020 gnd.n5670 gnd.n3104 21.0318
R8021 gnd.n5795 gnd.n3107 21.0318
R8022 gnd.n3119 gnd.n3113 21.0318
R8023 gnd.n5783 gnd.n3120 21.0318
R8024 gnd.n5782 gnd.n3123 21.0318
R8025 gnd.n5777 gnd.n3130 21.0318
R8026 gnd.n7541 gnd.n71 21.0318
R8027 gnd.n5770 gnd.n5769 21.0318
R8028 gnd.n5697 gnd.n86 21.0318
R8029 gnd.n7533 gnd.n89 21.0318
R8030 gnd.n7527 gnd.n101 21.0318
R8031 gnd.n5712 gnd.n108 21.0318
R8032 gnd.n5755 gnd.n117 21.0318
R8033 gnd.n7515 gnd.n120 21.0318
R8034 gnd.n5749 gnd.n128 21.0318
R8035 gnd.n7509 gnd.n131 21.0318
R8036 gnd.n7503 gnd.n141 21.0318
R8037 gnd.n5737 gnd.n149 21.0318
R8038 gnd.n7497 gnd.n152 21.0318
R8039 gnd.n5731 gnd.n159 21.0318
R8040 gnd.n7478 gnd.n168 21.0318
R8041 gnd.n7485 gnd.n171 21.0318
R8042 gnd.t48 gnd.n1013 20.7131
R8043 gnd.n4211 gnd.t15 20.7131
R8044 gnd.t4 gnd.n2486 20.7131
R8045 gnd.t51 gnd.n5790 20.7131
R8046 gnd.n5703 gnd.t2 20.7131
R8047 gnd.n6084 gnd.n2676 20.3945
R8048 gnd.n3020 gnd.n3012 20.3945
R8049 gnd.t21 gnd.n1047 20.0758
R8050 gnd.n4148 gnd.t126 20.0758
R8051 gnd.t23 gnd.n2523 20.0758
R8052 gnd.t45 gnd.n3075 20.0758
R8053 gnd.n5743 gnd.t0 20.0758
R8054 gnd.n3610 gnd.n3609 19.9763
R8055 gnd.n3301 gnd.n3300 19.9763
R8056 gnd.n5966 gnd.n5965 19.9763
R8057 gnd.n5251 gnd.n5250 19.9763
R8058 gnd.n2894 gnd.t173 19.8005
R8059 gnd.n2894 gnd.t226 19.8005
R8060 gnd.n2893 gnd.t290 19.8005
R8061 gnd.n2893 gnd.t253 19.8005
R8062 gnd.n5241 gnd.t199 19.8005
R8063 gnd.n5241 gnd.t268 19.8005
R8064 gnd.n5240 gnd.t243 19.8005
R8065 gnd.n5240 gnd.t284 19.8005
R8066 gnd.n2890 gnd.n2889 19.5087
R8067 gnd.n2903 gnd.n2890 19.5087
R8068 gnd.n2901 gnd.n2892 19.5087
R8069 gnd.n5245 gnd.n5239 19.5087
R8070 gnd.n1766 gnd.t67 19.4385
R8071 gnd.n4385 gnd.n4383 19.3944
R8072 gnd.n4390 gnd.n4383 19.3944
R8073 gnd.n4390 gnd.n4384 19.3944
R8074 gnd.n4384 gnd.n3727 19.3944
R8075 gnd.n4415 gnd.n3727 19.3944
R8076 gnd.n4415 gnd.n3724 19.3944
R8077 gnd.n4420 gnd.n3724 19.3944
R8078 gnd.n4420 gnd.n3725 19.3944
R8079 gnd.n3725 gnd.n3703 19.3944
R8080 gnd.n4445 gnd.n3703 19.3944
R8081 gnd.n4445 gnd.n3700 19.3944
R8082 gnd.n4450 gnd.n3700 19.3944
R8083 gnd.n4450 gnd.n3701 19.3944
R8084 gnd.n3701 gnd.n3678 19.3944
R8085 gnd.n4485 gnd.n3678 19.3944
R8086 gnd.n4485 gnd.n3675 19.3944
R8087 gnd.n4493 gnd.n3675 19.3944
R8088 gnd.n4493 gnd.n3676 19.3944
R8089 gnd.n4489 gnd.n3676 19.3944
R8090 gnd.n4489 gnd.n3594 19.3944
R8091 gnd.n4541 gnd.n3594 19.3944
R8092 gnd.n4541 gnd.n3591 19.3944
R8093 gnd.n4565 gnd.n3591 19.3944
R8094 gnd.n4565 gnd.n3592 19.3944
R8095 gnd.n4561 gnd.n3592 19.3944
R8096 gnd.n4561 gnd.n4560 19.3944
R8097 gnd.n4560 gnd.n4559 19.3944
R8098 gnd.n4559 gnd.n4551 19.3944
R8099 gnd.n4555 gnd.n4551 19.3944
R8100 gnd.n4555 gnd.n4554 19.3944
R8101 gnd.n4554 gnd.n3544 19.3944
R8102 gnd.n3544 gnd.n3542 19.3944
R8103 gnd.n4643 gnd.n3542 19.3944
R8104 gnd.n4643 gnd.n3540 19.3944
R8105 gnd.n4647 gnd.n3540 19.3944
R8106 gnd.n4647 gnd.n3515 19.3944
R8107 gnd.n4695 gnd.n3515 19.3944
R8108 gnd.n4695 gnd.n3516 19.3944
R8109 gnd.n4691 gnd.n3516 19.3944
R8110 gnd.n4691 gnd.n3492 19.3944
R8111 gnd.n4753 gnd.n3492 19.3944
R8112 gnd.n4753 gnd.n3493 19.3944
R8113 gnd.n4749 gnd.n3493 19.3944
R8114 gnd.n4749 gnd.n4748 19.3944
R8115 gnd.n4748 gnd.n4747 19.3944
R8116 gnd.n4747 gnd.n4734 19.3944
R8117 gnd.n4743 gnd.n4734 19.3944
R8118 gnd.n4743 gnd.n4742 19.3944
R8119 gnd.n4742 gnd.n4741 19.3944
R8120 gnd.n4741 gnd.n3434 19.3944
R8121 gnd.n4861 gnd.n3434 19.3944
R8122 gnd.n4861 gnd.n3431 19.3944
R8123 gnd.n4866 gnd.n3431 19.3944
R8124 gnd.n4866 gnd.n3432 19.3944
R8125 gnd.n3432 gnd.n3405 19.3944
R8126 gnd.n4900 gnd.n3405 19.3944
R8127 gnd.n4900 gnd.n3402 19.3944
R8128 gnd.n4911 gnd.n3402 19.3944
R8129 gnd.n4911 gnd.n3403 19.3944
R8130 gnd.n4907 gnd.n3403 19.3944
R8131 gnd.n4907 gnd.n4906 19.3944
R8132 gnd.n4906 gnd.n3370 19.3944
R8133 gnd.n4957 gnd.n3370 19.3944
R8134 gnd.n4957 gnd.n3368 19.3944
R8135 gnd.n4961 gnd.n3368 19.3944
R8136 gnd.n4964 gnd.n4961 19.3944
R8137 gnd.n4965 gnd.n4964 19.3944
R8138 gnd.n4965 gnd.n3366 19.3944
R8139 gnd.n4969 gnd.n3366 19.3944
R8140 gnd.n4972 gnd.n4969 19.3944
R8141 gnd.n4973 gnd.n4972 19.3944
R8142 gnd.n4973 gnd.n3364 19.3944
R8143 gnd.n4977 gnd.n3364 19.3944
R8144 gnd.n4980 gnd.n4977 19.3944
R8145 gnd.n4981 gnd.n4980 19.3944
R8146 gnd.n4981 gnd.n3362 19.3944
R8147 gnd.n4985 gnd.n3362 19.3944
R8148 gnd.n4988 gnd.n4985 19.3944
R8149 gnd.n4989 gnd.n4988 19.3944
R8150 gnd.n4989 gnd.n3359 19.3944
R8151 gnd.n5172 gnd.n3359 19.3944
R8152 gnd.n5172 gnd.n3360 19.3944
R8153 gnd.n2668 gnd.n2584 19.3944
R8154 gnd.n6153 gnd.n2584 19.3944
R8155 gnd.n6153 gnd.n6152 19.3944
R8156 gnd.n6146 gnd.n6145 19.3944
R8157 gnd.n6145 gnd.n2606 19.3944
R8158 gnd.n6141 gnd.n2606 19.3944
R8159 gnd.n6141 gnd.n6140 19.3944
R8160 gnd.n6140 gnd.n6139 19.3944
R8161 gnd.n6139 gnd.n2611 19.3944
R8162 gnd.n6134 gnd.n2611 19.3944
R8163 gnd.n6134 gnd.n6133 19.3944
R8164 gnd.n6133 gnd.n6132 19.3944
R8165 gnd.n6132 gnd.n2617 19.3944
R8166 gnd.n6125 gnd.n2617 19.3944
R8167 gnd.n6125 gnd.n6124 19.3944
R8168 gnd.n6124 gnd.n2629 19.3944
R8169 gnd.n6117 gnd.n2629 19.3944
R8170 gnd.n6117 gnd.n6116 19.3944
R8171 gnd.n6116 gnd.n2637 19.3944
R8172 gnd.n6109 gnd.n2637 19.3944
R8173 gnd.n6109 gnd.n6108 19.3944
R8174 gnd.n6108 gnd.n2647 19.3944
R8175 gnd.n6101 gnd.n2647 19.3944
R8176 gnd.n6101 gnd.n6100 19.3944
R8177 gnd.n6100 gnd.n2655 19.3944
R8178 gnd.n6093 gnd.n2655 19.3944
R8179 gnd.n6093 gnd.n6092 19.3944
R8180 gnd.n5080 gnd.n5043 19.3944
R8181 gnd.n5093 gnd.n5043 19.3944
R8182 gnd.n5093 gnd.n5041 19.3944
R8183 gnd.n5099 gnd.n5041 19.3944
R8184 gnd.n5099 gnd.n5034 19.3944
R8185 gnd.n5112 gnd.n5034 19.3944
R8186 gnd.n5112 gnd.n5032 19.3944
R8187 gnd.n5118 gnd.n5032 19.3944
R8188 gnd.n5118 gnd.n5025 19.3944
R8189 gnd.n5131 gnd.n5025 19.3944
R8190 gnd.n5131 gnd.n5023 19.3944
R8191 gnd.n5137 gnd.n5023 19.3944
R8192 gnd.n5137 gnd.n5016 19.3944
R8193 gnd.n5151 gnd.n5016 19.3944
R8194 gnd.n5151 gnd.n5014 19.3944
R8195 gnd.n5157 gnd.n5014 19.3944
R8196 gnd.n1481 gnd.n1480 19.3944
R8197 gnd.n1480 gnd.n1479 19.3944
R8198 gnd.n1479 gnd.n1478 19.3944
R8199 gnd.n1478 gnd.n1476 19.3944
R8200 gnd.n1476 gnd.n1473 19.3944
R8201 gnd.n1473 gnd.n1472 19.3944
R8202 gnd.n1472 gnd.n1469 19.3944
R8203 gnd.n1469 gnd.n1468 19.3944
R8204 gnd.n1468 gnd.n1465 19.3944
R8205 gnd.n1465 gnd.n1464 19.3944
R8206 gnd.n1464 gnd.n1461 19.3944
R8207 gnd.n1461 gnd.n1460 19.3944
R8208 gnd.n1460 gnd.n1457 19.3944
R8209 gnd.n1457 gnd.n1456 19.3944
R8210 gnd.n1456 gnd.n1453 19.3944
R8211 gnd.n1453 gnd.n1452 19.3944
R8212 gnd.n1452 gnd.n1449 19.3944
R8213 gnd.n1449 gnd.n1448 19.3944
R8214 gnd.n1448 gnd.n1445 19.3944
R8215 gnd.n1445 gnd.n1444 19.3944
R8216 gnd.n1444 gnd.n1441 19.3944
R8217 gnd.n1441 gnd.n1440 19.3944
R8218 gnd.n1437 gnd.n1436 19.3944
R8219 gnd.n1436 gnd.n1392 19.3944
R8220 gnd.n1487 gnd.n1392 19.3944
R8221 gnd.n2255 gnd.n2254 19.3944
R8222 gnd.n2254 gnd.n2251 19.3944
R8223 gnd.n2251 gnd.n2250 19.3944
R8224 gnd.n2300 gnd.n2299 19.3944
R8225 gnd.n2299 gnd.n2298 19.3944
R8226 gnd.n2298 gnd.n2295 19.3944
R8227 gnd.n2295 gnd.n2294 19.3944
R8228 gnd.n2294 gnd.n2291 19.3944
R8229 gnd.n2291 gnd.n2290 19.3944
R8230 gnd.n2290 gnd.n2287 19.3944
R8231 gnd.n2287 gnd.n2286 19.3944
R8232 gnd.n2286 gnd.n2283 19.3944
R8233 gnd.n2283 gnd.n2282 19.3944
R8234 gnd.n2282 gnd.n2279 19.3944
R8235 gnd.n2279 gnd.n2278 19.3944
R8236 gnd.n2278 gnd.n2275 19.3944
R8237 gnd.n2275 gnd.n2274 19.3944
R8238 gnd.n2274 gnd.n2271 19.3944
R8239 gnd.n2271 gnd.n2270 19.3944
R8240 gnd.n2270 gnd.n2267 19.3944
R8241 gnd.n2267 gnd.n2266 19.3944
R8242 gnd.n2266 gnd.n2263 19.3944
R8243 gnd.n2263 gnd.n2262 19.3944
R8244 gnd.n2262 gnd.n2259 19.3944
R8245 gnd.n2259 gnd.n2258 19.3944
R8246 gnd.n1580 gnd.n1289 19.3944
R8247 gnd.n1590 gnd.n1289 19.3944
R8248 gnd.n1591 gnd.n1590 19.3944
R8249 gnd.n1591 gnd.n1270 19.3944
R8250 gnd.n1611 gnd.n1270 19.3944
R8251 gnd.n1611 gnd.n1262 19.3944
R8252 gnd.n1621 gnd.n1262 19.3944
R8253 gnd.n1622 gnd.n1621 19.3944
R8254 gnd.n1623 gnd.n1622 19.3944
R8255 gnd.n1623 gnd.n1245 19.3944
R8256 gnd.n1640 gnd.n1245 19.3944
R8257 gnd.n1643 gnd.n1640 19.3944
R8258 gnd.n1643 gnd.n1642 19.3944
R8259 gnd.n1642 gnd.n1218 19.3944
R8260 gnd.n1682 gnd.n1218 19.3944
R8261 gnd.n1682 gnd.n1215 19.3944
R8262 gnd.n1688 gnd.n1215 19.3944
R8263 gnd.n1689 gnd.n1688 19.3944
R8264 gnd.n1689 gnd.n1213 19.3944
R8265 gnd.n1695 gnd.n1213 19.3944
R8266 gnd.n1698 gnd.n1695 19.3944
R8267 gnd.n1700 gnd.n1698 19.3944
R8268 gnd.n1706 gnd.n1700 19.3944
R8269 gnd.n1706 gnd.n1705 19.3944
R8270 gnd.n1705 gnd.n1088 19.3944
R8271 gnd.n1772 gnd.n1088 19.3944
R8272 gnd.n1773 gnd.n1772 19.3944
R8273 gnd.n1773 gnd.n1081 19.3944
R8274 gnd.n1784 gnd.n1081 19.3944
R8275 gnd.n1785 gnd.n1784 19.3944
R8276 gnd.n1785 gnd.n1064 19.3944
R8277 gnd.n1064 gnd.n1062 19.3944
R8278 gnd.n1809 gnd.n1062 19.3944
R8279 gnd.n1810 gnd.n1809 19.3944
R8280 gnd.n1810 gnd.n1035 19.3944
R8281 gnd.n1859 gnd.n1035 19.3944
R8282 gnd.n1860 gnd.n1859 19.3944
R8283 gnd.n1860 gnd.n1028 19.3944
R8284 gnd.n1871 gnd.n1028 19.3944
R8285 gnd.n1872 gnd.n1871 19.3944
R8286 gnd.n1872 gnd.n1011 19.3944
R8287 gnd.n1011 gnd.n1009 19.3944
R8288 gnd.n1896 gnd.n1009 19.3944
R8289 gnd.n1897 gnd.n1896 19.3944
R8290 gnd.n1897 gnd.n981 19.3944
R8291 gnd.n1948 gnd.n981 19.3944
R8292 gnd.n1949 gnd.n1948 19.3944
R8293 gnd.n1949 gnd.n974 19.3944
R8294 gnd.n2216 gnd.n974 19.3944
R8295 gnd.n2217 gnd.n2216 19.3944
R8296 gnd.n2217 gnd.n955 19.3944
R8297 gnd.n2242 gnd.n955 19.3944
R8298 gnd.n2242 gnd.n956 19.3944
R8299 gnd.n1571 gnd.n1570 19.3944
R8300 gnd.n1570 gnd.n1303 19.3944
R8301 gnd.n1326 gnd.n1303 19.3944
R8302 gnd.n1329 gnd.n1326 19.3944
R8303 gnd.n1329 gnd.n1322 19.3944
R8304 gnd.n1333 gnd.n1322 19.3944
R8305 gnd.n1336 gnd.n1333 19.3944
R8306 gnd.n1339 gnd.n1336 19.3944
R8307 gnd.n1339 gnd.n1320 19.3944
R8308 gnd.n1343 gnd.n1320 19.3944
R8309 gnd.n1346 gnd.n1343 19.3944
R8310 gnd.n1349 gnd.n1346 19.3944
R8311 gnd.n1349 gnd.n1318 19.3944
R8312 gnd.n1353 gnd.n1318 19.3944
R8313 gnd.n1576 gnd.n1575 19.3944
R8314 gnd.n1575 gnd.n1279 19.3944
R8315 gnd.n1601 gnd.n1279 19.3944
R8316 gnd.n1601 gnd.n1277 19.3944
R8317 gnd.n1607 gnd.n1277 19.3944
R8318 gnd.n1607 gnd.n1606 19.3944
R8319 gnd.n1606 gnd.n1251 19.3944
R8320 gnd.n1631 gnd.n1251 19.3944
R8321 gnd.n1631 gnd.n1249 19.3944
R8322 gnd.n1635 gnd.n1249 19.3944
R8323 gnd.n1635 gnd.n1229 19.3944
R8324 gnd.n1662 gnd.n1229 19.3944
R8325 gnd.n1662 gnd.n1227 19.3944
R8326 gnd.n1672 gnd.n1227 19.3944
R8327 gnd.n1672 gnd.n1671 19.3944
R8328 gnd.n1671 gnd.n1670 19.3944
R8329 gnd.n1670 gnd.n1176 19.3944
R8330 gnd.n1720 gnd.n1176 19.3944
R8331 gnd.n1720 gnd.n1719 19.3944
R8332 gnd.n1719 gnd.n1718 19.3944
R8333 gnd.n1718 gnd.n1180 19.3944
R8334 gnd.n1200 gnd.n1180 19.3944
R8335 gnd.n1200 gnd.n1098 19.3944
R8336 gnd.n1757 gnd.n1098 19.3944
R8337 gnd.n1757 gnd.n1096 19.3944
R8338 gnd.n1763 gnd.n1096 19.3944
R8339 gnd.n1763 gnd.n1762 19.3944
R8340 gnd.n1762 gnd.n1071 19.3944
R8341 gnd.n1797 gnd.n1071 19.3944
R8342 gnd.n1797 gnd.n1069 19.3944
R8343 gnd.n1803 gnd.n1069 19.3944
R8344 gnd.n1803 gnd.n1802 19.3944
R8345 gnd.n1802 gnd.n1045 19.3944
R8346 gnd.n1844 gnd.n1045 19.3944
R8347 gnd.n1844 gnd.n1043 19.3944
R8348 gnd.n1850 gnd.n1043 19.3944
R8349 gnd.n1850 gnd.n1849 19.3944
R8350 gnd.n1849 gnd.n1018 19.3944
R8351 gnd.n1884 gnd.n1018 19.3944
R8352 gnd.n1884 gnd.n1016 19.3944
R8353 gnd.n1890 gnd.n1016 19.3944
R8354 gnd.n1890 gnd.n1889 19.3944
R8355 gnd.n1889 gnd.n991 19.3944
R8356 gnd.n1933 gnd.n991 19.3944
R8357 gnd.n1933 gnd.n989 19.3944
R8358 gnd.n1939 gnd.n989 19.3944
R8359 gnd.n1939 gnd.n1938 19.3944
R8360 gnd.n1938 gnd.n964 19.3944
R8361 gnd.n2227 gnd.n964 19.3944
R8362 gnd.n2227 gnd.n962 19.3944
R8363 gnd.n2235 gnd.n962 19.3944
R8364 gnd.n2235 gnd.n2234 19.3944
R8365 gnd.n2234 gnd.n2233 19.3944
R8366 gnd.n2336 gnd.n2335 19.3944
R8367 gnd.n2335 gnd.n903 19.3944
R8368 gnd.n2331 gnd.n903 19.3944
R8369 gnd.n2331 gnd.n2328 19.3944
R8370 gnd.n2328 gnd.n2325 19.3944
R8371 gnd.n2325 gnd.n2324 19.3944
R8372 gnd.n2324 gnd.n2321 19.3944
R8373 gnd.n2321 gnd.n2320 19.3944
R8374 gnd.n2320 gnd.n2317 19.3944
R8375 gnd.n2317 gnd.n2316 19.3944
R8376 gnd.n2316 gnd.n2313 19.3944
R8377 gnd.n2313 gnd.n2312 19.3944
R8378 gnd.n2312 gnd.n2309 19.3944
R8379 gnd.n2309 gnd.n2308 19.3944
R8380 gnd.n1491 gnd.n1390 19.3944
R8381 gnd.n1491 gnd.n1381 19.3944
R8382 gnd.n1504 gnd.n1381 19.3944
R8383 gnd.n1504 gnd.n1379 19.3944
R8384 gnd.n1508 gnd.n1379 19.3944
R8385 gnd.n1508 gnd.n1369 19.3944
R8386 gnd.n1520 gnd.n1369 19.3944
R8387 gnd.n1520 gnd.n1367 19.3944
R8388 gnd.n1554 gnd.n1367 19.3944
R8389 gnd.n1554 gnd.n1553 19.3944
R8390 gnd.n1553 gnd.n1552 19.3944
R8391 gnd.n1552 gnd.n1551 19.3944
R8392 gnd.n1551 gnd.n1548 19.3944
R8393 gnd.n1548 gnd.n1547 19.3944
R8394 gnd.n1547 gnd.n1546 19.3944
R8395 gnd.n1546 gnd.n1544 19.3944
R8396 gnd.n1544 gnd.n1543 19.3944
R8397 gnd.n1543 gnd.n1540 19.3944
R8398 gnd.n1540 gnd.n1539 19.3944
R8399 gnd.n1539 gnd.n1538 19.3944
R8400 gnd.n1538 gnd.n1536 19.3944
R8401 gnd.n1536 gnd.n1235 19.3944
R8402 gnd.n1651 gnd.n1235 19.3944
R8403 gnd.n1651 gnd.n1233 19.3944
R8404 gnd.n1657 gnd.n1233 19.3944
R8405 gnd.n1657 gnd.n1656 19.3944
R8406 gnd.n1656 gnd.n1157 19.3944
R8407 gnd.n1731 gnd.n1157 19.3944
R8408 gnd.n1731 gnd.n1158 19.3944
R8409 gnd.n1205 gnd.n1204 19.3944
R8410 gnd.n1208 gnd.n1207 19.3944
R8411 gnd.n1195 gnd.n1194 19.3944
R8412 gnd.n1750 gnd.n1103 19.3944
R8413 gnd.n1750 gnd.n1749 19.3944
R8414 gnd.n1749 gnd.n1748 19.3944
R8415 gnd.n1748 gnd.n1746 19.3944
R8416 gnd.n1746 gnd.n1745 19.3944
R8417 gnd.n1745 gnd.n1743 19.3944
R8418 gnd.n1743 gnd.n1742 19.3944
R8419 gnd.n1742 gnd.n1052 19.3944
R8420 gnd.n1818 gnd.n1052 19.3944
R8421 gnd.n1818 gnd.n1050 19.3944
R8422 gnd.n1837 gnd.n1050 19.3944
R8423 gnd.n1837 gnd.n1836 19.3944
R8424 gnd.n1836 gnd.n1835 19.3944
R8425 gnd.n1835 gnd.n1833 19.3944
R8426 gnd.n1833 gnd.n1832 19.3944
R8427 gnd.n1832 gnd.n1830 19.3944
R8428 gnd.n1830 gnd.n1829 19.3944
R8429 gnd.n1829 gnd.n998 19.3944
R8430 gnd.n1905 gnd.n998 19.3944
R8431 gnd.n1905 gnd.n996 19.3944
R8432 gnd.n1928 gnd.n996 19.3944
R8433 gnd.n1928 gnd.n1927 19.3944
R8434 gnd.n1927 gnd.n1926 19.3944
R8435 gnd.n1926 gnd.n1923 19.3944
R8436 gnd.n1923 gnd.n1922 19.3944
R8437 gnd.n1922 gnd.n1920 19.3944
R8438 gnd.n1920 gnd.n1919 19.3944
R8439 gnd.n1919 gnd.n1917 19.3944
R8440 gnd.n1917 gnd.n950 19.3944
R8441 gnd.n1496 gnd.n1386 19.3944
R8442 gnd.n1496 gnd.n1384 19.3944
R8443 gnd.n1500 gnd.n1384 19.3944
R8444 gnd.n1500 gnd.n1375 19.3944
R8445 gnd.n1512 gnd.n1375 19.3944
R8446 gnd.n1512 gnd.n1373 19.3944
R8447 gnd.n1516 gnd.n1373 19.3944
R8448 gnd.n1516 gnd.n1362 19.3944
R8449 gnd.n1558 gnd.n1362 19.3944
R8450 gnd.n1558 gnd.n1316 19.3944
R8451 gnd.n1564 gnd.n1316 19.3944
R8452 gnd.n1564 gnd.n1563 19.3944
R8453 gnd.n1563 gnd.n1294 19.3944
R8454 gnd.n1585 gnd.n1294 19.3944
R8455 gnd.n1585 gnd.n1287 19.3944
R8456 gnd.n1596 gnd.n1287 19.3944
R8457 gnd.n1596 gnd.n1595 19.3944
R8458 gnd.n1595 gnd.n1268 19.3944
R8459 gnd.n1616 gnd.n1268 19.3944
R8460 gnd.n1616 gnd.n1258 19.3944
R8461 gnd.n1626 gnd.n1258 19.3944
R8462 gnd.n1626 gnd.n1241 19.3944
R8463 gnd.n1647 gnd.n1241 19.3944
R8464 gnd.n1647 gnd.n1646 19.3944
R8465 gnd.n1646 gnd.n1220 19.3944
R8466 gnd.n1677 gnd.n1220 19.3944
R8467 gnd.n1677 gnd.n1165 19.3944
R8468 gnd.n1727 gnd.n1165 19.3944
R8469 gnd.n1727 gnd.n1726 19.3944
R8470 gnd.n1726 gnd.n1725 19.3944
R8471 gnd.n1725 gnd.n1169 19.3944
R8472 gnd.n1187 gnd.n1169 19.3944
R8473 gnd.n1713 gnd.n1187 19.3944
R8474 gnd.n1713 gnd.n1712 19.3944
R8475 gnd.n1712 gnd.n1711 19.3944
R8476 gnd.n1711 gnd.n1191 19.3944
R8477 gnd.n1191 gnd.n1090 19.3944
R8478 gnd.n1768 gnd.n1090 19.3944
R8479 gnd.n1768 gnd.n1083 19.3944
R8480 gnd.n1779 gnd.n1083 19.3944
R8481 gnd.n1779 gnd.n1079 19.3944
R8482 gnd.n1792 gnd.n1079 19.3944
R8483 gnd.n1792 gnd.n1791 19.3944
R8484 gnd.n1791 gnd.n1058 19.3944
R8485 gnd.n1814 gnd.n1058 19.3944
R8486 gnd.n1814 gnd.n1813 19.3944
R8487 gnd.n1813 gnd.n1037 19.3944
R8488 gnd.n1855 gnd.n1037 19.3944
R8489 gnd.n1855 gnd.n1030 19.3944
R8490 gnd.n1866 gnd.n1030 19.3944
R8491 gnd.n1866 gnd.n1026 19.3944
R8492 gnd.n1879 gnd.n1026 19.3944
R8493 gnd.n1879 gnd.n1878 19.3944
R8494 gnd.n1878 gnd.n1005 19.3944
R8495 gnd.n1901 gnd.n1005 19.3944
R8496 gnd.n1901 gnd.n1900 19.3944
R8497 gnd.n1900 gnd.n983 19.3944
R8498 gnd.n1944 gnd.n983 19.3944
R8499 gnd.n1944 gnd.n976 19.3944
R8500 gnd.n1955 gnd.n976 19.3944
R8501 gnd.n1955 gnd.n972 19.3944
R8502 gnd.n2222 gnd.n972 19.3944
R8503 gnd.n2222 gnd.n2221 19.3944
R8504 gnd.n2221 gnd.n953 19.3944
R8505 gnd.n2245 gnd.n953 19.3944
R8506 gnd.n6129 gnd.n2620 19.3944
R8507 gnd.n6129 gnd.n6128 19.3944
R8508 gnd.n6128 gnd.n2623 19.3944
R8509 gnd.n6121 gnd.n2623 19.3944
R8510 gnd.n6121 gnd.n6120 19.3944
R8511 gnd.n6120 gnd.n2633 19.3944
R8512 gnd.n6113 gnd.n2633 19.3944
R8513 gnd.n6113 gnd.n6112 19.3944
R8514 gnd.n6112 gnd.n2641 19.3944
R8515 gnd.n6105 gnd.n2641 19.3944
R8516 gnd.n6105 gnd.n6104 19.3944
R8517 gnd.n6104 gnd.n2651 19.3944
R8518 gnd.n6097 gnd.n2651 19.3944
R8519 gnd.n6097 gnd.n6096 19.3944
R8520 gnd.n6096 gnd.n2659 19.3944
R8521 gnd.n6089 gnd.n2659 19.3944
R8522 gnd.n7019 gnd.n392 19.3944
R8523 gnd.n7025 gnd.n392 19.3944
R8524 gnd.n7025 gnd.n390 19.3944
R8525 gnd.n7029 gnd.n390 19.3944
R8526 gnd.n7029 gnd.n386 19.3944
R8527 gnd.n7035 gnd.n386 19.3944
R8528 gnd.n7035 gnd.n384 19.3944
R8529 gnd.n7039 gnd.n384 19.3944
R8530 gnd.n7039 gnd.n380 19.3944
R8531 gnd.n7045 gnd.n380 19.3944
R8532 gnd.n7045 gnd.n378 19.3944
R8533 gnd.n7049 gnd.n378 19.3944
R8534 gnd.n7049 gnd.n374 19.3944
R8535 gnd.n7055 gnd.n374 19.3944
R8536 gnd.n7055 gnd.n372 19.3944
R8537 gnd.n7059 gnd.n372 19.3944
R8538 gnd.n7059 gnd.n368 19.3944
R8539 gnd.n7065 gnd.n368 19.3944
R8540 gnd.n7065 gnd.n366 19.3944
R8541 gnd.n7069 gnd.n366 19.3944
R8542 gnd.n7069 gnd.n362 19.3944
R8543 gnd.n7075 gnd.n362 19.3944
R8544 gnd.n7075 gnd.n360 19.3944
R8545 gnd.n7079 gnd.n360 19.3944
R8546 gnd.n7079 gnd.n356 19.3944
R8547 gnd.n7085 gnd.n356 19.3944
R8548 gnd.n7085 gnd.n354 19.3944
R8549 gnd.n7089 gnd.n354 19.3944
R8550 gnd.n7089 gnd.n350 19.3944
R8551 gnd.n7095 gnd.n350 19.3944
R8552 gnd.n7095 gnd.n348 19.3944
R8553 gnd.n7099 gnd.n348 19.3944
R8554 gnd.n7099 gnd.n344 19.3944
R8555 gnd.n7105 gnd.n344 19.3944
R8556 gnd.n7105 gnd.n342 19.3944
R8557 gnd.n7109 gnd.n342 19.3944
R8558 gnd.n7109 gnd.n338 19.3944
R8559 gnd.n7115 gnd.n338 19.3944
R8560 gnd.n7115 gnd.n336 19.3944
R8561 gnd.n7119 gnd.n336 19.3944
R8562 gnd.n7119 gnd.n332 19.3944
R8563 gnd.n7125 gnd.n332 19.3944
R8564 gnd.n7125 gnd.n330 19.3944
R8565 gnd.n7129 gnd.n330 19.3944
R8566 gnd.n7129 gnd.n326 19.3944
R8567 gnd.n7135 gnd.n326 19.3944
R8568 gnd.n7135 gnd.n324 19.3944
R8569 gnd.n7139 gnd.n324 19.3944
R8570 gnd.n7139 gnd.n320 19.3944
R8571 gnd.n7145 gnd.n320 19.3944
R8572 gnd.n7145 gnd.n318 19.3944
R8573 gnd.n7149 gnd.n318 19.3944
R8574 gnd.n7149 gnd.n314 19.3944
R8575 gnd.n7155 gnd.n314 19.3944
R8576 gnd.n7155 gnd.n312 19.3944
R8577 gnd.n7159 gnd.n312 19.3944
R8578 gnd.n7159 gnd.n308 19.3944
R8579 gnd.n7165 gnd.n308 19.3944
R8580 gnd.n7165 gnd.n306 19.3944
R8581 gnd.n7169 gnd.n306 19.3944
R8582 gnd.n7169 gnd.n302 19.3944
R8583 gnd.n7175 gnd.n302 19.3944
R8584 gnd.n7175 gnd.n300 19.3944
R8585 gnd.n7179 gnd.n300 19.3944
R8586 gnd.n7179 gnd.n296 19.3944
R8587 gnd.n7185 gnd.n296 19.3944
R8588 gnd.n7185 gnd.n294 19.3944
R8589 gnd.n7189 gnd.n294 19.3944
R8590 gnd.n7189 gnd.n290 19.3944
R8591 gnd.n7195 gnd.n290 19.3944
R8592 gnd.n7195 gnd.n288 19.3944
R8593 gnd.n7199 gnd.n288 19.3944
R8594 gnd.n7199 gnd.n284 19.3944
R8595 gnd.n7205 gnd.n284 19.3944
R8596 gnd.n7205 gnd.n282 19.3944
R8597 gnd.n7209 gnd.n282 19.3944
R8598 gnd.n7209 gnd.n278 19.3944
R8599 gnd.n7215 gnd.n278 19.3944
R8600 gnd.n7215 gnd.n276 19.3944
R8601 gnd.n7219 gnd.n276 19.3944
R8602 gnd.n7219 gnd.n272 19.3944
R8603 gnd.n7225 gnd.n272 19.3944
R8604 gnd.n7225 gnd.n270 19.3944
R8605 gnd.n7230 gnd.n270 19.3944
R8606 gnd.n6498 gnd.n703 19.3944
R8607 gnd.n6504 gnd.n703 19.3944
R8608 gnd.n6504 gnd.n701 19.3944
R8609 gnd.n6508 gnd.n701 19.3944
R8610 gnd.n6508 gnd.n697 19.3944
R8611 gnd.n6514 gnd.n697 19.3944
R8612 gnd.n6514 gnd.n695 19.3944
R8613 gnd.n6518 gnd.n695 19.3944
R8614 gnd.n6518 gnd.n691 19.3944
R8615 gnd.n6524 gnd.n691 19.3944
R8616 gnd.n6524 gnd.n689 19.3944
R8617 gnd.n6528 gnd.n689 19.3944
R8618 gnd.n6528 gnd.n685 19.3944
R8619 gnd.n6534 gnd.n685 19.3944
R8620 gnd.n6534 gnd.n683 19.3944
R8621 gnd.n6538 gnd.n683 19.3944
R8622 gnd.n6538 gnd.n679 19.3944
R8623 gnd.n6544 gnd.n679 19.3944
R8624 gnd.n6544 gnd.n677 19.3944
R8625 gnd.n6548 gnd.n677 19.3944
R8626 gnd.n6548 gnd.n673 19.3944
R8627 gnd.n6554 gnd.n673 19.3944
R8628 gnd.n6554 gnd.n671 19.3944
R8629 gnd.n6558 gnd.n671 19.3944
R8630 gnd.n6558 gnd.n667 19.3944
R8631 gnd.n6564 gnd.n667 19.3944
R8632 gnd.n6564 gnd.n665 19.3944
R8633 gnd.n6568 gnd.n665 19.3944
R8634 gnd.n6568 gnd.n661 19.3944
R8635 gnd.n6574 gnd.n661 19.3944
R8636 gnd.n6574 gnd.n659 19.3944
R8637 gnd.n6578 gnd.n659 19.3944
R8638 gnd.n6578 gnd.n655 19.3944
R8639 gnd.n6584 gnd.n655 19.3944
R8640 gnd.n6584 gnd.n653 19.3944
R8641 gnd.n6588 gnd.n653 19.3944
R8642 gnd.n6588 gnd.n649 19.3944
R8643 gnd.n6594 gnd.n649 19.3944
R8644 gnd.n6594 gnd.n647 19.3944
R8645 gnd.n6598 gnd.n647 19.3944
R8646 gnd.n6598 gnd.n643 19.3944
R8647 gnd.n6604 gnd.n643 19.3944
R8648 gnd.n6604 gnd.n641 19.3944
R8649 gnd.n6608 gnd.n641 19.3944
R8650 gnd.n6608 gnd.n637 19.3944
R8651 gnd.n6614 gnd.n637 19.3944
R8652 gnd.n6614 gnd.n635 19.3944
R8653 gnd.n6618 gnd.n635 19.3944
R8654 gnd.n6618 gnd.n631 19.3944
R8655 gnd.n6624 gnd.n631 19.3944
R8656 gnd.n6624 gnd.n629 19.3944
R8657 gnd.n6628 gnd.n629 19.3944
R8658 gnd.n6628 gnd.n625 19.3944
R8659 gnd.n6634 gnd.n625 19.3944
R8660 gnd.n6634 gnd.n623 19.3944
R8661 gnd.n6638 gnd.n623 19.3944
R8662 gnd.n6638 gnd.n619 19.3944
R8663 gnd.n6644 gnd.n619 19.3944
R8664 gnd.n6644 gnd.n617 19.3944
R8665 gnd.n6648 gnd.n617 19.3944
R8666 gnd.n6648 gnd.n613 19.3944
R8667 gnd.n6654 gnd.n613 19.3944
R8668 gnd.n6654 gnd.n611 19.3944
R8669 gnd.n6658 gnd.n611 19.3944
R8670 gnd.n6658 gnd.n607 19.3944
R8671 gnd.n6664 gnd.n607 19.3944
R8672 gnd.n6664 gnd.n605 19.3944
R8673 gnd.n6668 gnd.n605 19.3944
R8674 gnd.n6668 gnd.n601 19.3944
R8675 gnd.n6674 gnd.n601 19.3944
R8676 gnd.n6674 gnd.n599 19.3944
R8677 gnd.n6678 gnd.n599 19.3944
R8678 gnd.n6678 gnd.n595 19.3944
R8679 gnd.n6684 gnd.n595 19.3944
R8680 gnd.n6684 gnd.n593 19.3944
R8681 gnd.n6688 gnd.n593 19.3944
R8682 gnd.n6688 gnd.n589 19.3944
R8683 gnd.n6694 gnd.n589 19.3944
R8684 gnd.n6694 gnd.n587 19.3944
R8685 gnd.n6698 gnd.n587 19.3944
R8686 gnd.n6698 gnd.n583 19.3944
R8687 gnd.n6704 gnd.n583 19.3944
R8688 gnd.n6704 gnd.n581 19.3944
R8689 gnd.n6708 gnd.n581 19.3944
R8690 gnd.n6708 gnd.n577 19.3944
R8691 gnd.n6714 gnd.n577 19.3944
R8692 gnd.n6714 gnd.n575 19.3944
R8693 gnd.n6718 gnd.n575 19.3944
R8694 gnd.n6718 gnd.n571 19.3944
R8695 gnd.n6724 gnd.n571 19.3944
R8696 gnd.n6724 gnd.n569 19.3944
R8697 gnd.n6728 gnd.n569 19.3944
R8698 gnd.n6728 gnd.n565 19.3944
R8699 gnd.n6734 gnd.n565 19.3944
R8700 gnd.n6734 gnd.n563 19.3944
R8701 gnd.n6738 gnd.n563 19.3944
R8702 gnd.n6738 gnd.n559 19.3944
R8703 gnd.n6744 gnd.n559 19.3944
R8704 gnd.n6744 gnd.n557 19.3944
R8705 gnd.n6748 gnd.n557 19.3944
R8706 gnd.n6748 gnd.n553 19.3944
R8707 gnd.n6754 gnd.n553 19.3944
R8708 gnd.n6754 gnd.n551 19.3944
R8709 gnd.n6758 gnd.n551 19.3944
R8710 gnd.n6758 gnd.n547 19.3944
R8711 gnd.n6764 gnd.n547 19.3944
R8712 gnd.n6764 gnd.n545 19.3944
R8713 gnd.n6768 gnd.n545 19.3944
R8714 gnd.n6768 gnd.n541 19.3944
R8715 gnd.n6774 gnd.n541 19.3944
R8716 gnd.n6774 gnd.n539 19.3944
R8717 gnd.n6778 gnd.n539 19.3944
R8718 gnd.n6778 gnd.n535 19.3944
R8719 gnd.n6784 gnd.n535 19.3944
R8720 gnd.n6784 gnd.n533 19.3944
R8721 gnd.n6788 gnd.n533 19.3944
R8722 gnd.n6788 gnd.n529 19.3944
R8723 gnd.n6794 gnd.n529 19.3944
R8724 gnd.n6794 gnd.n527 19.3944
R8725 gnd.n6798 gnd.n527 19.3944
R8726 gnd.n6798 gnd.n523 19.3944
R8727 gnd.n6804 gnd.n523 19.3944
R8728 gnd.n6804 gnd.n521 19.3944
R8729 gnd.n6808 gnd.n521 19.3944
R8730 gnd.n6808 gnd.n517 19.3944
R8731 gnd.n6814 gnd.n517 19.3944
R8732 gnd.n6814 gnd.n515 19.3944
R8733 gnd.n6818 gnd.n515 19.3944
R8734 gnd.n6818 gnd.n511 19.3944
R8735 gnd.n6824 gnd.n511 19.3944
R8736 gnd.n6824 gnd.n509 19.3944
R8737 gnd.n6828 gnd.n509 19.3944
R8738 gnd.n6828 gnd.n505 19.3944
R8739 gnd.n6834 gnd.n505 19.3944
R8740 gnd.n6834 gnd.n503 19.3944
R8741 gnd.n6838 gnd.n503 19.3944
R8742 gnd.n6838 gnd.n499 19.3944
R8743 gnd.n6844 gnd.n499 19.3944
R8744 gnd.n6844 gnd.n497 19.3944
R8745 gnd.n6848 gnd.n497 19.3944
R8746 gnd.n6848 gnd.n493 19.3944
R8747 gnd.n6854 gnd.n493 19.3944
R8748 gnd.n6854 gnd.n491 19.3944
R8749 gnd.n6858 gnd.n491 19.3944
R8750 gnd.n6858 gnd.n487 19.3944
R8751 gnd.n6864 gnd.n487 19.3944
R8752 gnd.n6864 gnd.n485 19.3944
R8753 gnd.n6868 gnd.n485 19.3944
R8754 gnd.n6868 gnd.n481 19.3944
R8755 gnd.n6874 gnd.n481 19.3944
R8756 gnd.n6874 gnd.n479 19.3944
R8757 gnd.n6878 gnd.n479 19.3944
R8758 gnd.n6878 gnd.n475 19.3944
R8759 gnd.n6884 gnd.n475 19.3944
R8760 gnd.n6884 gnd.n473 19.3944
R8761 gnd.n6888 gnd.n473 19.3944
R8762 gnd.n6888 gnd.n469 19.3944
R8763 gnd.n6894 gnd.n469 19.3944
R8764 gnd.n6894 gnd.n467 19.3944
R8765 gnd.n6898 gnd.n467 19.3944
R8766 gnd.n6898 gnd.n463 19.3944
R8767 gnd.n6904 gnd.n463 19.3944
R8768 gnd.n6904 gnd.n461 19.3944
R8769 gnd.n6908 gnd.n461 19.3944
R8770 gnd.n6908 gnd.n457 19.3944
R8771 gnd.n6914 gnd.n457 19.3944
R8772 gnd.n6914 gnd.n455 19.3944
R8773 gnd.n6918 gnd.n455 19.3944
R8774 gnd.n6918 gnd.n451 19.3944
R8775 gnd.n6924 gnd.n451 19.3944
R8776 gnd.n6924 gnd.n449 19.3944
R8777 gnd.n6928 gnd.n449 19.3944
R8778 gnd.n6928 gnd.n445 19.3944
R8779 gnd.n6934 gnd.n445 19.3944
R8780 gnd.n6934 gnd.n443 19.3944
R8781 gnd.n6938 gnd.n443 19.3944
R8782 gnd.n6938 gnd.n439 19.3944
R8783 gnd.n6944 gnd.n439 19.3944
R8784 gnd.n6944 gnd.n437 19.3944
R8785 gnd.n6948 gnd.n437 19.3944
R8786 gnd.n6948 gnd.n433 19.3944
R8787 gnd.n6954 gnd.n433 19.3944
R8788 gnd.n6954 gnd.n431 19.3944
R8789 gnd.n6958 gnd.n431 19.3944
R8790 gnd.n6958 gnd.n427 19.3944
R8791 gnd.n6964 gnd.n427 19.3944
R8792 gnd.n6964 gnd.n425 19.3944
R8793 gnd.n6968 gnd.n425 19.3944
R8794 gnd.n6968 gnd.n421 19.3944
R8795 gnd.n6974 gnd.n421 19.3944
R8796 gnd.n6974 gnd.n419 19.3944
R8797 gnd.n6978 gnd.n419 19.3944
R8798 gnd.n6978 gnd.n415 19.3944
R8799 gnd.n6984 gnd.n415 19.3944
R8800 gnd.n6984 gnd.n413 19.3944
R8801 gnd.n6988 gnd.n413 19.3944
R8802 gnd.n6988 gnd.n409 19.3944
R8803 gnd.n6994 gnd.n409 19.3944
R8804 gnd.n6994 gnd.n407 19.3944
R8805 gnd.n6998 gnd.n407 19.3944
R8806 gnd.n6998 gnd.n403 19.3944
R8807 gnd.n7004 gnd.n403 19.3944
R8808 gnd.n7004 gnd.n401 19.3944
R8809 gnd.n7009 gnd.n401 19.3944
R8810 gnd.n7009 gnd.n397 19.3944
R8811 gnd.n7015 gnd.n397 19.3944
R8812 gnd.n7016 gnd.n7015 19.3944
R8813 gnd.n5416 gnd.n5413 19.3944
R8814 gnd.n5416 gnd.n5412 19.3944
R8815 gnd.n5422 gnd.n5412 19.3944
R8816 gnd.n5422 gnd.n5410 19.3944
R8817 gnd.n5426 gnd.n5410 19.3944
R8818 gnd.n5426 gnd.n5408 19.3944
R8819 gnd.n5432 gnd.n5408 19.3944
R8820 gnd.n5432 gnd.n5406 19.3944
R8821 gnd.n5436 gnd.n5406 19.3944
R8822 gnd.n5436 gnd.n5404 19.3944
R8823 gnd.n5442 gnd.n5404 19.3944
R8824 gnd.n5442 gnd.n5402 19.3944
R8825 gnd.n5446 gnd.n5402 19.3944
R8826 gnd.n5446 gnd.n5400 19.3944
R8827 gnd.n5452 gnd.n5400 19.3944
R8828 gnd.n5452 gnd.n5398 19.3944
R8829 gnd.n5459 gnd.n5398 19.3944
R8830 gnd.n5465 gnd.n5396 19.3944
R8831 gnd.n5465 gnd.n5394 19.3944
R8832 gnd.n5469 gnd.n5394 19.3944
R8833 gnd.n5469 gnd.n5392 19.3944
R8834 gnd.n5475 gnd.n5392 19.3944
R8835 gnd.n5475 gnd.n5390 19.3944
R8836 gnd.n5480 gnd.n5390 19.3944
R8837 gnd.n5488 gnd.n3262 19.3944
R8838 gnd.n5488 gnd.n3260 19.3944
R8839 gnd.n5492 gnd.n3260 19.3944
R8840 gnd.n5492 gnd.n3258 19.3944
R8841 gnd.n5498 gnd.n3258 19.3944
R8842 gnd.n5498 gnd.n3256 19.3944
R8843 gnd.n5502 gnd.n3256 19.3944
R8844 gnd.n5502 gnd.n3254 19.3944
R8845 gnd.n5514 gnd.n3252 19.3944
R8846 gnd.n5514 gnd.n3250 19.3944
R8847 gnd.n5520 gnd.n3250 19.3944
R8848 gnd.n5520 gnd.n3248 19.3944
R8849 gnd.n5524 gnd.n3248 19.3944
R8850 gnd.n5524 gnd.n3246 19.3944
R8851 gnd.n5530 gnd.n3246 19.3944
R8852 gnd.n5530 gnd.n3244 19.3944
R8853 gnd.n5534 gnd.n3244 19.3944
R8854 gnd.n5534 gnd.n3242 19.3944
R8855 gnd.n5540 gnd.n3242 19.3944
R8856 gnd.n5540 gnd.n3240 19.3944
R8857 gnd.n5544 gnd.n3240 19.3944
R8858 gnd.n5544 gnd.n3238 19.3944
R8859 gnd.n5550 gnd.n3238 19.3944
R8860 gnd.n5550 gnd.n3236 19.3944
R8861 gnd.n5555 gnd.n3236 19.3944
R8862 gnd.n5555 gnd.n3234 19.3944
R8863 gnd.n5568 gnd.n3227 19.3944
R8864 gnd.n5569 gnd.n5568 19.3944
R8865 gnd.n5570 gnd.n5569 19.3944
R8866 gnd.n5570 gnd.n3222 19.3944
R8867 gnd.n5582 gnd.n3222 19.3944
R8868 gnd.n5583 gnd.n5582 19.3944
R8869 gnd.n5584 gnd.n5583 19.3944
R8870 gnd.n5585 gnd.n5584 19.3944
R8871 gnd.n5587 gnd.n5585 19.3944
R8872 gnd.n5587 gnd.n3210 19.3944
R8873 gnd.n5647 gnd.n3210 19.3944
R8874 gnd.n5648 gnd.n5647 19.3944
R8875 gnd.n5650 gnd.n5648 19.3944
R8876 gnd.n5650 gnd.n3204 19.3944
R8877 gnd.n5672 gnd.n3204 19.3944
R8878 gnd.n5673 gnd.n5672 19.3944
R8879 gnd.n5674 gnd.n5673 19.3944
R8880 gnd.n5677 gnd.n5674 19.3944
R8881 gnd.n5677 gnd.n3202 19.3944
R8882 gnd.n5685 gnd.n3202 19.3944
R8883 gnd.n5686 gnd.n5685 19.3944
R8884 gnd.n5689 gnd.n5686 19.3944
R8885 gnd.n5690 gnd.n5689 19.3944
R8886 gnd.n5691 gnd.n5690 19.3944
R8887 gnd.n5699 gnd.n5691 19.3944
R8888 gnd.n5700 gnd.n5699 19.3944
R8889 gnd.n5701 gnd.n5700 19.3944
R8890 gnd.n5701 gnd.n3197 19.3944
R8891 gnd.n5714 gnd.n3197 19.3944
R8892 gnd.n5715 gnd.n5714 19.3944
R8893 gnd.n5716 gnd.n5715 19.3944
R8894 gnd.n5717 gnd.n5716 19.3944
R8895 gnd.n5747 gnd.n5717 19.3944
R8896 gnd.n5747 gnd.n5746 19.3944
R8897 gnd.n5746 gnd.n5745 19.3944
R8898 gnd.n5745 gnd.n5719 19.3944
R8899 gnd.n5735 gnd.n5719 19.3944
R8900 gnd.n5735 gnd.n5734 19.3944
R8901 gnd.n5734 gnd.n5733 19.3944
R8902 gnd.n5733 gnd.n175 19.3944
R8903 gnd.n7480 gnd.n175 19.3944
R8904 gnd.n7481 gnd.n7480 19.3944
R8905 gnd.n5565 gnd.n3038 19.3944
R8906 gnd.n5835 gnd.n3038 19.3944
R8907 gnd.n5835 gnd.n5834 19.3944
R8908 gnd.n5834 gnd.n5833 19.3944
R8909 gnd.n5833 gnd.n3042 19.3944
R8910 gnd.n5823 gnd.n3042 19.3944
R8911 gnd.n5823 gnd.n5822 19.3944
R8912 gnd.n5822 gnd.n5821 19.3944
R8913 gnd.n5821 gnd.n3062 19.3944
R8914 gnd.n5811 gnd.n3062 19.3944
R8915 gnd.n5811 gnd.n5810 19.3944
R8916 gnd.n5810 gnd.n5809 19.3944
R8917 gnd.n5809 gnd.n3083 19.3944
R8918 gnd.n5799 gnd.n3083 19.3944
R8919 gnd.n5799 gnd.n5798 19.3944
R8920 gnd.n5798 gnd.n5797 19.3944
R8921 gnd.n5797 gnd.n3102 19.3944
R8922 gnd.n5679 gnd.n3102 19.3944
R8923 gnd.n5682 gnd.n5679 19.3944
R8924 gnd.n5682 gnd.n3132 19.3944
R8925 gnd.n5775 gnd.n3132 19.3944
R8926 gnd.n5775 gnd.n5774 19.3944
R8927 gnd.n5774 gnd.n5773 19.3944
R8928 gnd.n5773 gnd.n5772 19.3944
R8929 gnd.n5772 gnd.n92 19.3944
R8930 gnd.n7531 gnd.n92 19.3944
R8931 gnd.n7531 gnd.n7530 19.3944
R8932 gnd.n7530 gnd.n7529 19.3944
R8933 gnd.n7529 gnd.n96 19.3944
R8934 gnd.n7519 gnd.n96 19.3944
R8935 gnd.n7519 gnd.n7518 19.3944
R8936 gnd.n7518 gnd.n7517 19.3944
R8937 gnd.n7517 gnd.n115 19.3944
R8938 gnd.n7507 gnd.n115 19.3944
R8939 gnd.n7507 gnd.n7506 19.3944
R8940 gnd.n7506 gnd.n7505 19.3944
R8941 gnd.n7505 gnd.n136 19.3944
R8942 gnd.n7495 gnd.n136 19.3944
R8943 gnd.n7495 gnd.n7494 19.3944
R8944 gnd.n7494 gnd.n7493 19.3944
R8945 gnd.n7493 gnd.n157 19.3944
R8946 gnd.n7483 gnd.n157 19.3944
R8947 gnd.n7390 gnd.n7326 19.3944
R8948 gnd.n7390 gnd.n7387 19.3944
R8949 gnd.n7387 gnd.n7384 19.3944
R8950 gnd.n7384 gnd.n7383 19.3944
R8951 gnd.n7383 gnd.n7380 19.3944
R8952 gnd.n7380 gnd.n7379 19.3944
R8953 gnd.n7379 gnd.n7376 19.3944
R8954 gnd.n7376 gnd.n7375 19.3944
R8955 gnd.n7375 gnd.n7372 19.3944
R8956 gnd.n7372 gnd.n7371 19.3944
R8957 gnd.n7371 gnd.n7368 19.3944
R8958 gnd.n7368 gnd.n7367 19.3944
R8959 gnd.n7367 gnd.n7364 19.3944
R8960 gnd.n7364 gnd.n7363 19.3944
R8961 gnd.n7363 gnd.n7360 19.3944
R8962 gnd.n7360 gnd.n7359 19.3944
R8963 gnd.n7359 gnd.n7356 19.3944
R8964 gnd.n7356 gnd.n7355 19.3944
R8965 gnd.n7433 gnd.n7430 19.3944
R8966 gnd.n7430 gnd.n7429 19.3944
R8967 gnd.n7429 gnd.n7426 19.3944
R8968 gnd.n7426 gnd.n7425 19.3944
R8969 gnd.n7425 gnd.n7422 19.3944
R8970 gnd.n7422 gnd.n7421 19.3944
R8971 gnd.n7421 gnd.n7418 19.3944
R8972 gnd.n7418 gnd.n7417 19.3944
R8973 gnd.n7417 gnd.n7414 19.3944
R8974 gnd.n7414 gnd.n7413 19.3944
R8975 gnd.n7413 gnd.n7410 19.3944
R8976 gnd.n7410 gnd.n7409 19.3944
R8977 gnd.n7409 gnd.n7406 19.3944
R8978 gnd.n7406 gnd.n7405 19.3944
R8979 gnd.n7405 gnd.n7402 19.3944
R8980 gnd.n7402 gnd.n7401 19.3944
R8981 gnd.n7401 gnd.n7398 19.3944
R8982 gnd.n7398 gnd.n7397 19.3944
R8983 gnd.n7288 gnd.n7287 19.3944
R8984 gnd.n7466 gnd.n7287 19.3944
R8985 gnd.n7466 gnd.n7465 19.3944
R8986 gnd.n7465 gnd.n7464 19.3944
R8987 gnd.n7464 gnd.n7461 19.3944
R8988 gnd.n7461 gnd.n7460 19.3944
R8989 gnd.n7460 gnd.n7457 19.3944
R8990 gnd.n7457 gnd.n7456 19.3944
R8991 gnd.n7456 gnd.n7453 19.3944
R8992 gnd.n7453 gnd.n7452 19.3944
R8993 gnd.n7452 gnd.n7449 19.3944
R8994 gnd.n7449 gnd.n7448 19.3944
R8995 gnd.n7448 gnd.n7445 19.3944
R8996 gnd.n7445 gnd.n7444 19.3944
R8997 gnd.n7444 gnd.n7441 19.3944
R8998 gnd.n7441 gnd.n7440 19.3944
R8999 gnd.n7440 gnd.n7437 19.3944
R9000 gnd.n204 gnd.n202 19.3944
R9001 gnd.n207 gnd.n204 19.3944
R9002 gnd.n207 gnd.n199 19.3944
R9003 gnd.n211 gnd.n199 19.3944
R9004 gnd.n214 gnd.n211 19.3944
R9005 gnd.n217 gnd.n214 19.3944
R9006 gnd.n217 gnd.n197 19.3944
R9007 gnd.n221 gnd.n197 19.3944
R9008 gnd.n224 gnd.n221 19.3944
R9009 gnd.n227 gnd.n224 19.3944
R9010 gnd.n227 gnd.n195 19.3944
R9011 gnd.n231 gnd.n195 19.3944
R9012 gnd.n234 gnd.n231 19.3944
R9013 gnd.n236 gnd.n234 19.3944
R9014 gnd.n236 gnd.n193 19.3944
R9015 gnd.n240 gnd.n193 19.3944
R9016 gnd.n4996 gnd.n4995 19.3944
R9017 gnd.n4995 gnd.n3226 19.3944
R9018 gnd.n5574 gnd.n3226 19.3944
R9019 gnd.n5574 gnd.n3224 19.3944
R9020 gnd.n5578 gnd.n3224 19.3944
R9021 gnd.n5578 gnd.n3218 19.3944
R9022 gnd.n5598 gnd.n3218 19.3944
R9023 gnd.n5598 gnd.n3219 19.3944
R9024 gnd.n5594 gnd.n3219 19.3944
R9025 gnd.n5594 gnd.n5593 19.3944
R9026 gnd.n5593 gnd.n5592 19.3944
R9027 gnd.n5592 gnd.n3209 19.3944
R9028 gnd.n5654 gnd.n3209 19.3944
R9029 gnd.n5654 gnd.n3206 19.3944
R9030 gnd.n5668 gnd.n3206 19.3944
R9031 gnd.n5668 gnd.n3207 19.3944
R9032 gnd.n5664 gnd.n3207 19.3944
R9033 gnd.n5664 gnd.n5663 19.3944
R9034 gnd.n5663 gnd.n5662 19.3944
R9035 gnd.n5662 gnd.n5660 19.3944
R9036 gnd.n5660 gnd.n64 19.3944
R9037 gnd.n7544 gnd.n64 19.3944
R9038 gnd.n7544 gnd.n7543 19.3944
R9039 gnd.n7543 gnd.n67 19.3944
R9040 gnd.n5695 gnd.n67 19.3944
R9041 gnd.n5695 gnd.n3201 19.3944
R9042 gnd.n5705 gnd.n3201 19.3944
R9043 gnd.n5705 gnd.n3199 19.3944
R9044 gnd.n5710 gnd.n3199 19.3944
R9045 gnd.n5710 gnd.n3192 19.3944
R9046 gnd.n5753 gnd.n3192 19.3944
R9047 gnd.n5753 gnd.n5752 19.3944
R9048 gnd.n5752 gnd.n5751 19.3944
R9049 gnd.n5751 gnd.n3196 19.3944
R9050 gnd.n5741 gnd.n3196 19.3944
R9051 gnd.n5741 gnd.n5740 19.3944
R9052 gnd.n5740 gnd.n5739 19.3944
R9053 gnd.n5739 gnd.n5724 19.3944
R9054 gnd.n5729 gnd.n5724 19.3944
R9055 gnd.n5729 gnd.n177 19.3944
R9056 gnd.n7476 gnd.n177 19.3944
R9057 gnd.n7476 gnd.n7475 19.3944
R9058 gnd.n5841 gnd.n5840 19.3944
R9059 gnd.n5840 gnd.n5839 19.3944
R9060 gnd.n5839 gnd.n3030 19.3944
R9061 gnd.n5829 gnd.n3030 19.3944
R9062 gnd.n5829 gnd.n5828 19.3944
R9063 gnd.n5828 gnd.n5827 19.3944
R9064 gnd.n5827 gnd.n3053 19.3944
R9065 gnd.n5817 gnd.n3053 19.3944
R9066 gnd.n5817 gnd.n5816 19.3944
R9067 gnd.n5816 gnd.n5815 19.3944
R9068 gnd.n5815 gnd.n3073 19.3944
R9069 gnd.n5805 gnd.n3073 19.3944
R9070 gnd.n5805 gnd.n5804 19.3944
R9071 gnd.n5804 gnd.n5803 19.3944
R9072 gnd.n5803 gnd.n3093 19.3944
R9073 gnd.n5793 gnd.n3093 19.3944
R9074 gnd.n3110 gnd.n3109 19.3944
R9075 gnd.n5780 gnd.n5779 19.3944
R9076 gnd.n3127 gnd.n3126 19.3944
R9077 gnd.n7539 gnd.n7538 19.3944
R9078 gnd.n7535 gnd.n76 19.3944
R9079 gnd.n7535 gnd.n83 19.3944
R9080 gnd.n7525 gnd.n83 19.3944
R9081 gnd.n7525 gnd.n7524 19.3944
R9082 gnd.n7524 gnd.n7523 19.3944
R9083 gnd.n7523 gnd.n106 19.3944
R9084 gnd.n7513 gnd.n106 19.3944
R9085 gnd.n7513 gnd.n7512 19.3944
R9086 gnd.n7512 gnd.n7511 19.3944
R9087 gnd.n7511 gnd.n126 19.3944
R9088 gnd.n7501 gnd.n126 19.3944
R9089 gnd.n7501 gnd.n7500 19.3944
R9090 gnd.n7500 gnd.n7499 19.3944
R9091 gnd.n7499 gnd.n147 19.3944
R9092 gnd.n7489 gnd.n147 19.3944
R9093 gnd.n7489 gnd.n7488 19.3944
R9094 gnd.n7488 gnd.n7487 19.3944
R9095 gnd.n6324 gnd.n875 19.3944
R9096 gnd.n6318 gnd.n875 19.3944
R9097 gnd.n6318 gnd.n6317 19.3944
R9098 gnd.n6317 gnd.n6316 19.3944
R9099 gnd.n6316 gnd.n2345 19.3944
R9100 gnd.n6310 gnd.n2345 19.3944
R9101 gnd.n6310 gnd.n6309 19.3944
R9102 gnd.n6309 gnd.n6308 19.3944
R9103 gnd.n6308 gnd.n2353 19.3944
R9104 gnd.n6302 gnd.n2353 19.3944
R9105 gnd.n6302 gnd.n6301 19.3944
R9106 gnd.n6301 gnd.n6300 19.3944
R9107 gnd.n6300 gnd.n2361 19.3944
R9108 gnd.n3832 gnd.n2361 19.3944
R9109 gnd.n4169 gnd.n3832 19.3944
R9110 gnd.n4169 gnd.n3829 19.3944
R9111 gnd.n4173 gnd.n3829 19.3944
R9112 gnd.n4173 gnd.n3827 19.3944
R9113 gnd.n4177 gnd.n3827 19.3944
R9114 gnd.n4177 gnd.n3825 19.3944
R9115 gnd.n4181 gnd.n3825 19.3944
R9116 gnd.n4181 gnd.n3823 19.3944
R9117 gnd.n4185 gnd.n3823 19.3944
R9118 gnd.n4185 gnd.n3821 19.3944
R9119 gnd.n4194 gnd.n3821 19.3944
R9120 gnd.n4194 gnd.n4193 19.3944
R9121 gnd.n4193 gnd.n4192 19.3944
R9122 gnd.n4192 gnd.n3794 19.3944
R9123 gnd.n4273 gnd.n3794 19.3944
R9124 gnd.n4273 gnd.n3795 19.3944
R9125 gnd.n4269 gnd.n4268 19.3944
R9126 gnd.n3799 gnd.n3798 19.3944
R9127 gnd.n4239 gnd.n4238 19.3944
R9128 gnd.n4236 gnd.n4235 19.3944
R9129 gnd.n4232 gnd.n3787 19.3944
R9130 gnd.n4280 gnd.n3787 19.3944
R9131 gnd.n4280 gnd.n4279 19.3944
R9132 gnd.n4279 gnd.n3767 19.3944
R9133 gnd.n4334 gnd.n3767 19.3944
R9134 gnd.n4334 gnd.n3765 19.3944
R9135 gnd.n4338 gnd.n3765 19.3944
R9136 gnd.n4338 gnd.n3763 19.3944
R9137 gnd.n4342 gnd.n3763 19.3944
R9138 gnd.n4342 gnd.n3761 19.3944
R9139 gnd.n4346 gnd.n3761 19.3944
R9140 gnd.n4346 gnd.n3759 19.3944
R9141 gnd.n4350 gnd.n3759 19.3944
R9142 gnd.n4350 gnd.n3757 19.3944
R9143 gnd.n4354 gnd.n3757 19.3944
R9144 gnd.n4354 gnd.n3755 19.3944
R9145 gnd.n4358 gnd.n3755 19.3944
R9146 gnd.n4358 gnd.n3753 19.3944
R9147 gnd.n4362 gnd.n3753 19.3944
R9148 gnd.n4362 gnd.n3751 19.3944
R9149 gnd.n4367 gnd.n3751 19.3944
R9150 gnd.n4367 gnd.n3749 19.3944
R9151 gnd.n4371 gnd.n3749 19.3944
R9152 gnd.n4371 gnd.n3746 19.3944
R9153 gnd.n4395 gnd.n3746 19.3944
R9154 gnd.n4395 gnd.n3744 19.3944
R9155 gnd.n4401 gnd.n3744 19.3944
R9156 gnd.n4401 gnd.n4400 19.3944
R9157 gnd.n4400 gnd.n3721 19.3944
R9158 gnd.n4425 gnd.n3721 19.3944
R9159 gnd.n4425 gnd.n3719 19.3944
R9160 gnd.n4431 gnd.n3719 19.3944
R9161 gnd.n4431 gnd.n4430 19.3944
R9162 gnd.n4430 gnd.n3696 19.3944
R9163 gnd.n4455 gnd.n3696 19.3944
R9164 gnd.n4455 gnd.n3694 19.3944
R9165 gnd.n4471 gnd.n3694 19.3944
R9166 gnd.n4471 gnd.n4470 19.3944
R9167 gnd.n4470 gnd.n4469 19.3944
R9168 gnd.n4469 gnd.n4461 19.3944
R9169 gnd.n4464 gnd.n4461 19.3944
R9170 gnd.n4464 gnd.n3602 19.3944
R9171 gnd.n4530 gnd.n3602 19.3944
R9172 gnd.n4530 gnd.n3600 19.3944
R9173 gnd.n4536 gnd.n3600 19.3944
R9174 gnd.n4536 gnd.n4535 19.3944
R9175 gnd.n4535 gnd.n3576 19.3944
R9176 gnd.n4592 gnd.n3576 19.3944
R9177 gnd.n4592 gnd.n3574 19.3944
R9178 gnd.n4596 gnd.n3574 19.3944
R9179 gnd.n4596 gnd.n3558 19.3944
R9180 gnd.n4619 gnd.n3558 19.3944
R9181 gnd.n4619 gnd.n3556 19.3944
R9182 gnd.n4625 gnd.n3556 19.3944
R9183 gnd.n4625 gnd.n4624 19.3944
R9184 gnd.n4624 gnd.n3525 19.3944
R9185 gnd.n4670 gnd.n3525 19.3944
R9186 gnd.n4670 gnd.n3523 19.3944
R9187 gnd.n4674 gnd.n3523 19.3944
R9188 gnd.n4674 gnd.n3502 19.3944
R9189 gnd.n4710 gnd.n3502 19.3944
R9190 gnd.n4710 gnd.n3500 19.3944
R9191 gnd.n4714 gnd.n3500 19.3944
R9192 gnd.n4714 gnd.n3480 19.3944
R9193 gnd.n4766 gnd.n3480 19.3944
R9194 gnd.n4766 gnd.n3478 19.3944
R9195 gnd.n4770 gnd.n3478 19.3944
R9196 gnd.n4770 gnd.n3461 19.3944
R9197 gnd.n4791 gnd.n3461 19.3944
R9198 gnd.n4791 gnd.n3459 19.3944
R9199 gnd.n4795 gnd.n3459 19.3944
R9200 gnd.n4795 gnd.n3441 19.3944
R9201 gnd.n4851 gnd.n3441 19.3944
R9202 gnd.n4851 gnd.n3439 19.3944
R9203 gnd.n4855 gnd.n3439 19.3944
R9204 gnd.n4855 gnd.n3419 19.3944
R9205 gnd.n4880 gnd.n3419 19.3944
R9206 gnd.n4880 gnd.n3417 19.3944
R9207 gnd.n4886 gnd.n3417 19.3944
R9208 gnd.n4886 gnd.n4885 19.3944
R9209 gnd.n4885 gnd.n3391 19.3944
R9210 gnd.n4925 gnd.n3391 19.3944
R9211 gnd.n4925 gnd.n3389 19.3944
R9212 gnd.n4935 gnd.n3389 19.3944
R9213 gnd.n4935 gnd.n4934 19.3944
R9214 gnd.n4934 gnd.n4933 19.3944
R9215 gnd.n4933 gnd.n3315 19.3944
R9216 gnd.n5222 gnd.n3315 19.3944
R9217 gnd.n5222 gnd.n5221 19.3944
R9218 gnd.n5221 gnd.n5220 19.3944
R9219 gnd.n5220 gnd.n3319 19.3944
R9220 gnd.n5211 gnd.n3319 19.3944
R9221 gnd.n5211 gnd.n5210 19.3944
R9222 gnd.n5210 gnd.n5209 19.3944
R9223 gnd.n5209 gnd.n3329 19.3944
R9224 gnd.n5200 gnd.n3329 19.3944
R9225 gnd.n5200 gnd.n5199 19.3944
R9226 gnd.n5199 gnd.n5198 19.3944
R9227 gnd.n5198 gnd.n3341 19.3944
R9228 gnd.n5189 gnd.n3341 19.3944
R9229 gnd.n5189 gnd.n5188 19.3944
R9230 gnd.n5188 gnd.n5187 19.3944
R9231 gnd.n5187 gnd.n3353 19.3944
R9232 gnd.n5178 gnd.n3353 19.3944
R9233 gnd.n5178 gnd.n3005 19.3944
R9234 gnd.n5856 gnd.n3005 19.3944
R9235 gnd.n5856 gnd.n5855 19.3944
R9236 gnd.n5855 gnd.n5854 19.3944
R9237 gnd.n5854 gnd.n3009 19.3944
R9238 gnd.n5848 gnd.n3009 19.3944
R9239 gnd.n5848 gnd.n5847 19.3944
R9240 gnd.n5847 gnd.n5846 19.3944
R9241 gnd.n5846 gnd.n3018 19.3944
R9242 gnd.n5610 gnd.n3018 19.3944
R9243 gnd.n5610 gnd.n5607 19.3944
R9244 gnd.n5614 gnd.n5607 19.3944
R9245 gnd.n5614 gnd.n5605 19.3944
R9246 gnd.n5618 gnd.n5605 19.3944
R9247 gnd.n5618 gnd.n5603 19.3944
R9248 gnd.n5622 gnd.n5603 19.3944
R9249 gnd.n5622 gnd.n3216 19.3944
R9250 gnd.n5626 gnd.n3216 19.3944
R9251 gnd.n5626 gnd.n3214 19.3944
R9252 gnd.n5642 gnd.n3214 19.3944
R9253 gnd.n5642 gnd.n5641 19.3944
R9254 gnd.n5641 gnd.n5640 19.3944
R9255 gnd.n5640 gnd.n5632 19.3944
R9256 gnd.n5636 gnd.n5632 19.3944
R9257 gnd.n5636 gnd.n5635 19.3944
R9258 gnd.n5788 gnd.n5787 19.3944
R9259 gnd.n5785 gnd.n3117 19.3944
R9260 gnd.n3144 gnd.n3141 19.3944
R9261 gnd.n5767 gnd.n3146 19.3944
R9262 gnd.n5765 gnd.n5764 19.3944
R9263 gnd.n5764 gnd.n3148 19.3944
R9264 gnd.n5760 gnd.n3148 19.3944
R9265 gnd.n5760 gnd.n5759 19.3944
R9266 gnd.n5759 gnd.n5758 19.3944
R9267 gnd.n5758 gnd.n3154 19.3944
R9268 gnd.n3188 gnd.n3154 19.3944
R9269 gnd.n3188 gnd.n3187 19.3944
R9270 gnd.n3187 gnd.n3186 19.3944
R9271 gnd.n3186 gnd.n3160 19.3944
R9272 gnd.n3182 gnd.n3160 19.3944
R9273 gnd.n3182 gnd.n3181 19.3944
R9274 gnd.n3181 gnd.n3180 19.3944
R9275 gnd.n3180 gnd.n3166 19.3944
R9276 gnd.n3176 gnd.n3166 19.3944
R9277 gnd.n3176 gnd.n3175 19.3944
R9278 gnd.n3175 gnd.n3174 19.3944
R9279 gnd.n3174 gnd.n246 19.3944
R9280 gnd.n7254 gnd.n246 19.3944
R9281 gnd.n7254 gnd.n7253 19.3944
R9282 gnd.n7253 gnd.n7252 19.3944
R9283 gnd.n7252 gnd.n250 19.3944
R9284 gnd.n7246 gnd.n250 19.3944
R9285 gnd.n7246 gnd.n7245 19.3944
R9286 gnd.n7245 gnd.n7244 19.3944
R9287 gnd.n7244 gnd.n258 19.3944
R9288 gnd.n7238 gnd.n258 19.3944
R9289 gnd.n7238 gnd.n7237 19.3944
R9290 gnd.n7237 gnd.n7236 19.3944
R9291 gnd.n7236 gnd.n266 19.3944
R9292 gnd.n3976 gnd.n3973 19.3944
R9293 gnd.n3976 gnd.n3971 19.3944
R9294 gnd.n3980 gnd.n3971 19.3944
R9295 gnd.n3980 gnd.n3969 19.3944
R9296 gnd.n3986 gnd.n3969 19.3944
R9297 gnd.n3986 gnd.n3967 19.3944
R9298 gnd.n3990 gnd.n3967 19.3944
R9299 gnd.n3990 gnd.n3965 19.3944
R9300 gnd.n3996 gnd.n3965 19.3944
R9301 gnd.n3996 gnd.n3963 19.3944
R9302 gnd.n4000 gnd.n3963 19.3944
R9303 gnd.n4000 gnd.n3961 19.3944
R9304 gnd.n4006 gnd.n3961 19.3944
R9305 gnd.n4006 gnd.n3959 19.3944
R9306 gnd.n4010 gnd.n3959 19.3944
R9307 gnd.n4010 gnd.n3954 19.3944
R9308 gnd.n4016 gnd.n3954 19.3944
R9309 gnd.n4020 gnd.n3952 19.3944
R9310 gnd.n4020 gnd.n3950 19.3944
R9311 gnd.n4026 gnd.n3950 19.3944
R9312 gnd.n4026 gnd.n3948 19.3944
R9313 gnd.n4030 gnd.n3948 19.3944
R9314 gnd.n4030 gnd.n3946 19.3944
R9315 gnd.n4036 gnd.n3946 19.3944
R9316 gnd.n4036 gnd.n3944 19.3944
R9317 gnd.n4040 gnd.n3944 19.3944
R9318 gnd.n4040 gnd.n3942 19.3944
R9319 gnd.n4046 gnd.n3942 19.3944
R9320 gnd.n4046 gnd.n3940 19.3944
R9321 gnd.n4050 gnd.n3940 19.3944
R9322 gnd.n4050 gnd.n3938 19.3944
R9323 gnd.n4056 gnd.n3938 19.3944
R9324 gnd.n4056 gnd.n3936 19.3944
R9325 gnd.n4060 gnd.n3936 19.3944
R9326 gnd.n4060 gnd.n3934 19.3944
R9327 gnd.n4072 gnd.n3932 19.3944
R9328 gnd.n4072 gnd.n3930 19.3944
R9329 gnd.n4078 gnd.n3930 19.3944
R9330 gnd.n4078 gnd.n3928 19.3944
R9331 gnd.n4082 gnd.n3928 19.3944
R9332 gnd.n4082 gnd.n3926 19.3944
R9333 gnd.n4088 gnd.n3926 19.3944
R9334 gnd.n4088 gnd.n3924 19.3944
R9335 gnd.n4092 gnd.n3924 19.3944
R9336 gnd.n4092 gnd.n3922 19.3944
R9337 gnd.n4098 gnd.n3922 19.3944
R9338 gnd.n4098 gnd.n3920 19.3944
R9339 gnd.n4102 gnd.n3920 19.3944
R9340 gnd.n4102 gnd.n3918 19.3944
R9341 gnd.n4108 gnd.n3918 19.3944
R9342 gnd.n4108 gnd.n3916 19.3944
R9343 gnd.n4113 gnd.n3916 19.3944
R9344 gnd.n4113 gnd.n3914 19.3944
R9345 gnd.n3908 gnd.n3842 19.3944
R9346 gnd.n3903 gnd.n3842 19.3944
R9347 gnd.n3903 gnd.n3902 19.3944
R9348 gnd.n3902 gnd.n3846 19.3944
R9349 gnd.n3897 gnd.n3846 19.3944
R9350 gnd.n3897 gnd.n3896 19.3944
R9351 gnd.n3896 gnd.n3895 19.3944
R9352 gnd.n3895 gnd.n3852 19.3944
R9353 gnd.n3889 gnd.n3852 19.3944
R9354 gnd.n3889 gnd.n3888 19.3944
R9355 gnd.n3888 gnd.n3887 19.3944
R9356 gnd.n3887 gnd.n3858 19.3944
R9357 gnd.n3881 gnd.n3858 19.3944
R9358 gnd.n3881 gnd.n3880 19.3944
R9359 gnd.n3880 gnd.n3879 19.3944
R9360 gnd.n3879 gnd.n3864 19.3944
R9361 gnd.n4164 gnd.n3835 19.3944
R9362 gnd.n4164 gnd.n4163 19.3944
R9363 gnd.n4163 gnd.n4162 19.3944
R9364 gnd.n4162 gnd.n3839 19.3944
R9365 gnd.n4152 gnd.n3839 19.3944
R9366 gnd.n4152 gnd.n4151 19.3944
R9367 gnd.n4151 gnd.n4150 19.3944
R9368 gnd.n4150 gnd.n4134 19.3944
R9369 gnd.n4140 gnd.n4134 19.3944
R9370 gnd.n4140 gnd.n3817 19.3944
R9371 gnd.n4199 gnd.n3817 19.3944
R9372 gnd.n4199 gnd.n3815 19.3944
R9373 gnd.n4203 gnd.n3815 19.3944
R9374 gnd.n4203 gnd.n3812 19.3944
R9375 gnd.n4213 gnd.n3812 19.3944
R9376 gnd.n4213 gnd.n3810 19.3944
R9377 gnd.n4218 gnd.n3810 19.3944
R9378 gnd.n4218 gnd.n3801 19.3944
R9379 gnd.n4262 gnd.n3801 19.3944
R9380 gnd.n4262 gnd.n4261 19.3944
R9381 gnd.n4261 gnd.n4260 19.3944
R9382 gnd.n4260 gnd.n3805 19.3944
R9383 gnd.n4256 gnd.n3805 19.3944
R9384 gnd.n4256 gnd.n4255 19.3944
R9385 gnd.n4255 gnd.n4254 19.3944
R9386 gnd.n4254 gnd.n3783 19.3944
R9387 gnd.n4285 gnd.n3783 19.3944
R9388 gnd.n4285 gnd.n3781 19.3944
R9389 gnd.n4289 gnd.n3781 19.3944
R9390 gnd.n4289 gnd.n3770 19.3944
R9391 gnd.n4329 gnd.n3770 19.3944
R9392 gnd.n4329 gnd.n3771 19.3944
R9393 gnd.n4325 gnd.n3771 19.3944
R9394 gnd.n4325 gnd.n4324 19.3944
R9395 gnd.n4324 gnd.n4323 19.3944
R9396 gnd.n4323 gnd.n3776 19.3944
R9397 gnd.n4319 gnd.n3776 19.3944
R9398 gnd.n4319 gnd.n4318 19.3944
R9399 gnd.n4318 gnd.n4317 19.3944
R9400 gnd.n4317 gnd.n2579 19.3944
R9401 gnd.n6158 gnd.n2579 19.3944
R9402 gnd.n6158 gnd.n2580 19.3944
R9403 gnd.n4126 gnd.n3840 19.3944
R9404 gnd.n4127 gnd.n4126 19.3944
R9405 gnd.n4158 gnd.n4127 19.3944
R9406 gnd.n4158 gnd.n4157 19.3944
R9407 gnd.n4157 gnd.n4156 19.3944
R9408 gnd.n4156 gnd.n4129 19.3944
R9409 gnd.n4146 gnd.n4129 19.3944
R9410 gnd.n4146 gnd.n4145 19.3944
R9411 gnd.n4145 gnd.n4144 19.3944
R9412 gnd.n4144 gnd.n4137 19.3944
R9413 gnd.n4137 gnd.n4136 19.3944
R9414 gnd.n4136 gnd.n3813 19.3944
R9415 gnd.n4207 gnd.n3813 19.3944
R9416 gnd.n4208 gnd.n4207 19.3944
R9417 gnd.n4209 gnd.n4208 19.3944
R9418 gnd.n4209 gnd.n3808 19.3944
R9419 gnd.n4222 gnd.n3808 19.3944
R9420 gnd.n4223 gnd.n4222 19.3944
R9421 gnd.n4224 gnd.n4223 19.3944
R9422 gnd.n4225 gnd.n4224 19.3944
R9423 gnd.n4229 gnd.n4225 19.3944
R9424 gnd.n4230 gnd.n4229 19.3944
R9425 gnd.n4244 gnd.n4230 19.3944
R9426 gnd.n4245 gnd.n4244 19.3944
R9427 gnd.n4249 gnd.n4245 19.3944
R9428 gnd.n4249 gnd.n4248 19.3944
R9429 gnd.n4248 gnd.n4247 19.3944
R9430 gnd.n4247 gnd.n3779 19.3944
R9431 gnd.n4293 gnd.n3779 19.3944
R9432 gnd.n4294 gnd.n4293 19.3944
R9433 gnd.n4295 gnd.n4294 19.3944
R9434 gnd.n4296 gnd.n4295 19.3944
R9435 gnd.n4300 gnd.n4296 19.3944
R9436 gnd.n4301 gnd.n4300 19.3944
R9437 gnd.n4305 gnd.n4301 19.3944
R9438 gnd.n4306 gnd.n4305 19.3944
R9439 gnd.n4310 gnd.n4306 19.3944
R9440 gnd.n4311 gnd.n4310 19.3944
R9441 gnd.n4312 gnd.n4311 19.3944
R9442 gnd.n4312 gnd.n2578 19.3944
R9443 gnd.n6162 gnd.n2578 19.3944
R9444 gnd.n6163 gnd.n6162 19.3944
R9445 gnd.n4123 gnd.n2380 19.3944
R9446 gnd.n6288 gnd.n2380 19.3944
R9447 gnd.n6288 gnd.n6287 19.3944
R9448 gnd.n6287 gnd.n6286 19.3944
R9449 gnd.n6286 gnd.n2384 19.3944
R9450 gnd.n6276 gnd.n2384 19.3944
R9451 gnd.n6276 gnd.n6275 19.3944
R9452 gnd.n6275 gnd.n6274 19.3944
R9453 gnd.n6274 gnd.n2405 19.3944
R9454 gnd.n6264 gnd.n2405 19.3944
R9455 gnd.n6264 gnd.n6263 19.3944
R9456 gnd.n6263 gnd.n6262 19.3944
R9457 gnd.n6262 gnd.n2426 19.3944
R9458 gnd.n6252 gnd.n2426 19.3944
R9459 gnd.n6252 gnd.n6251 19.3944
R9460 gnd.n6251 gnd.n6250 19.3944
R9461 gnd.n6250 gnd.n2446 19.3944
R9462 gnd.n6239 gnd.n2446 19.3944
R9463 gnd.n6239 gnd.n6238 19.3944
R9464 gnd.n6238 gnd.n6237 19.3944
R9465 gnd.n6237 gnd.n2465 19.3944
R9466 gnd.n6226 gnd.n2465 19.3944
R9467 gnd.n6226 gnd.n6225 19.3944
R9468 gnd.n6225 gnd.n6224 19.3944
R9469 gnd.n6224 gnd.n2481 19.3944
R9470 gnd.n6213 gnd.n2481 19.3944
R9471 gnd.n6213 gnd.n6212 19.3944
R9472 gnd.n6212 gnd.n6211 19.3944
R9473 gnd.n6211 gnd.n2499 19.3944
R9474 gnd.n6201 gnd.n2499 19.3944
R9475 gnd.n6201 gnd.n6200 19.3944
R9476 gnd.n6200 gnd.n6199 19.3944
R9477 gnd.n6199 gnd.n2518 19.3944
R9478 gnd.n6189 gnd.n2518 19.3944
R9479 gnd.n6189 gnd.n6188 19.3944
R9480 gnd.n6188 gnd.n6187 19.3944
R9481 gnd.n6187 gnd.n2539 19.3944
R9482 gnd.n6177 gnd.n2539 19.3944
R9483 gnd.n6177 gnd.n6176 19.3944
R9484 gnd.n6176 gnd.n6175 19.3944
R9485 gnd.n6175 gnd.n2559 19.3944
R9486 gnd.n6165 gnd.n2559 19.3944
R9487 gnd.n2722 gnd.n2721 19.3944
R9488 gnd.n6081 gnd.n2721 19.3944
R9489 gnd.n6081 gnd.n6080 19.3944
R9490 gnd.n6080 gnd.n6079 19.3944
R9491 gnd.n6079 gnd.n6076 19.3944
R9492 gnd.n6076 gnd.n6075 19.3944
R9493 gnd.n6075 gnd.n6072 19.3944
R9494 gnd.n6072 gnd.n6071 19.3944
R9495 gnd.n6071 gnd.n6068 19.3944
R9496 gnd.n6068 gnd.n6067 19.3944
R9497 gnd.n6067 gnd.n6064 19.3944
R9498 gnd.n6064 gnd.n6063 19.3944
R9499 gnd.n6063 gnd.n6060 19.3944
R9500 gnd.n6060 gnd.n6059 19.3944
R9501 gnd.n6059 gnd.n6056 19.3944
R9502 gnd.n6056 gnd.n6055 19.3944
R9503 gnd.n6055 gnd.n6052 19.3944
R9504 gnd.n2824 gnd.n2760 19.3944
R9505 gnd.n2824 gnd.n2821 19.3944
R9506 gnd.n2821 gnd.n2818 19.3944
R9507 gnd.n2818 gnd.n2817 19.3944
R9508 gnd.n2817 gnd.n2814 19.3944
R9509 gnd.n2814 gnd.n2813 19.3944
R9510 gnd.n2813 gnd.n2810 19.3944
R9511 gnd.n2810 gnd.n2809 19.3944
R9512 gnd.n2809 gnd.n2806 19.3944
R9513 gnd.n2806 gnd.n2805 19.3944
R9514 gnd.n2805 gnd.n2802 19.3944
R9515 gnd.n2802 gnd.n2801 19.3944
R9516 gnd.n2801 gnd.n2798 19.3944
R9517 gnd.n2798 gnd.n2797 19.3944
R9518 gnd.n2797 gnd.n2794 19.3944
R9519 gnd.n2794 gnd.n2793 19.3944
R9520 gnd.n2793 gnd.n2790 19.3944
R9521 gnd.n2790 gnd.n2789 19.3944
R9522 gnd.n2846 gnd.n2751 19.3944
R9523 gnd.n2846 gnd.n2843 19.3944
R9524 gnd.n2843 gnd.n2840 19.3944
R9525 gnd.n2840 gnd.n2839 19.3944
R9526 gnd.n2839 gnd.n2836 19.3944
R9527 gnd.n2836 gnd.n2835 19.3944
R9528 gnd.n2835 gnd.n2832 19.3944
R9529 gnd.n2832 gnd.n2831 19.3944
R9530 gnd.n6050 gnd.n6047 19.3944
R9531 gnd.n6047 gnd.n6046 19.3944
R9532 gnd.n6046 gnd.n6043 19.3944
R9533 gnd.n6043 gnd.n6042 19.3944
R9534 gnd.n6042 gnd.n6039 19.3944
R9535 gnd.n6039 gnd.n6038 19.3944
R9536 gnd.n6038 gnd.n6035 19.3944
R9537 gnd.n6294 gnd.n6293 19.3944
R9538 gnd.n6293 gnd.n6292 19.3944
R9539 gnd.n6292 gnd.n2373 19.3944
R9540 gnd.n6282 gnd.n2373 19.3944
R9541 gnd.n6282 gnd.n6281 19.3944
R9542 gnd.n6281 gnd.n6280 19.3944
R9543 gnd.n6280 gnd.n2395 19.3944
R9544 gnd.n6270 gnd.n2395 19.3944
R9545 gnd.n6270 gnd.n6269 19.3944
R9546 gnd.n6269 gnd.n6268 19.3944
R9547 gnd.n6268 gnd.n2416 19.3944
R9548 gnd.n6258 gnd.n2416 19.3944
R9549 gnd.n6258 gnd.n6257 19.3944
R9550 gnd.n6257 gnd.n6256 19.3944
R9551 gnd.n6256 gnd.n2436 19.3944
R9552 gnd.n6246 gnd.n2436 19.3944
R9553 gnd.n6244 gnd.n6243 19.3944
R9554 gnd.n6233 gnd.n2471 19.3944
R9555 gnd.n6231 gnd.n6230 19.3944
R9556 gnd.n6220 gnd.n2488 19.3944
R9557 gnd.n6218 gnd.n6217 19.3944
R9558 gnd.n6217 gnd.n2489 19.3944
R9559 gnd.n6207 gnd.n2489 19.3944
R9560 gnd.n6207 gnd.n6206 19.3944
R9561 gnd.n6206 gnd.n6205 19.3944
R9562 gnd.n6205 gnd.n2509 19.3944
R9563 gnd.n6195 gnd.n2509 19.3944
R9564 gnd.n6195 gnd.n6194 19.3944
R9565 gnd.n6194 gnd.n6193 19.3944
R9566 gnd.n6193 gnd.n2529 19.3944
R9567 gnd.n6183 gnd.n2529 19.3944
R9568 gnd.n6183 gnd.n6182 19.3944
R9569 gnd.n6182 gnd.n6181 19.3944
R9570 gnd.n6181 gnd.n2549 19.3944
R9571 gnd.n6171 gnd.n2549 19.3944
R9572 gnd.n6171 gnd.n6170 19.3944
R9573 gnd.n6170 gnd.n6169 19.3944
R9574 gnd.n6495 gnd.n6494 19.3944
R9575 gnd.n6494 gnd.n708 19.3944
R9576 gnd.n6488 gnd.n708 19.3944
R9577 gnd.n6488 gnd.n6487 19.3944
R9578 gnd.n6487 gnd.n6486 19.3944
R9579 gnd.n6486 gnd.n716 19.3944
R9580 gnd.n6480 gnd.n716 19.3944
R9581 gnd.n6480 gnd.n6479 19.3944
R9582 gnd.n6479 gnd.n6478 19.3944
R9583 gnd.n6478 gnd.n724 19.3944
R9584 gnd.n6472 gnd.n724 19.3944
R9585 gnd.n6472 gnd.n6471 19.3944
R9586 gnd.n6471 gnd.n6470 19.3944
R9587 gnd.n6470 gnd.n732 19.3944
R9588 gnd.n6464 gnd.n732 19.3944
R9589 gnd.n6464 gnd.n6463 19.3944
R9590 gnd.n6463 gnd.n6462 19.3944
R9591 gnd.n6462 gnd.n740 19.3944
R9592 gnd.n6456 gnd.n740 19.3944
R9593 gnd.n6456 gnd.n6455 19.3944
R9594 gnd.n6455 gnd.n6454 19.3944
R9595 gnd.n6454 gnd.n748 19.3944
R9596 gnd.n6448 gnd.n748 19.3944
R9597 gnd.n6448 gnd.n6447 19.3944
R9598 gnd.n6447 gnd.n6446 19.3944
R9599 gnd.n6446 gnd.n756 19.3944
R9600 gnd.n6440 gnd.n756 19.3944
R9601 gnd.n6440 gnd.n6439 19.3944
R9602 gnd.n6439 gnd.n6438 19.3944
R9603 gnd.n6438 gnd.n764 19.3944
R9604 gnd.n6432 gnd.n764 19.3944
R9605 gnd.n6432 gnd.n6431 19.3944
R9606 gnd.n6431 gnd.n6430 19.3944
R9607 gnd.n6430 gnd.n772 19.3944
R9608 gnd.n6424 gnd.n772 19.3944
R9609 gnd.n6424 gnd.n6423 19.3944
R9610 gnd.n6423 gnd.n6422 19.3944
R9611 gnd.n6422 gnd.n780 19.3944
R9612 gnd.n6416 gnd.n780 19.3944
R9613 gnd.n6416 gnd.n6415 19.3944
R9614 gnd.n6415 gnd.n6414 19.3944
R9615 gnd.n6414 gnd.n788 19.3944
R9616 gnd.n6408 gnd.n788 19.3944
R9617 gnd.n6408 gnd.n6407 19.3944
R9618 gnd.n6407 gnd.n6406 19.3944
R9619 gnd.n6406 gnd.n796 19.3944
R9620 gnd.n6400 gnd.n796 19.3944
R9621 gnd.n6400 gnd.n6399 19.3944
R9622 gnd.n6399 gnd.n6398 19.3944
R9623 gnd.n6398 gnd.n804 19.3944
R9624 gnd.n6392 gnd.n804 19.3944
R9625 gnd.n6392 gnd.n6391 19.3944
R9626 gnd.n6391 gnd.n6390 19.3944
R9627 gnd.n6390 gnd.n812 19.3944
R9628 gnd.n6384 gnd.n812 19.3944
R9629 gnd.n6384 gnd.n6383 19.3944
R9630 gnd.n6383 gnd.n6382 19.3944
R9631 gnd.n6382 gnd.n820 19.3944
R9632 gnd.n6376 gnd.n820 19.3944
R9633 gnd.n6376 gnd.n6375 19.3944
R9634 gnd.n6375 gnd.n6374 19.3944
R9635 gnd.n6374 gnd.n828 19.3944
R9636 gnd.n6368 gnd.n828 19.3944
R9637 gnd.n6368 gnd.n6367 19.3944
R9638 gnd.n6367 gnd.n6366 19.3944
R9639 gnd.n6366 gnd.n836 19.3944
R9640 gnd.n6360 gnd.n836 19.3944
R9641 gnd.n6360 gnd.n6359 19.3944
R9642 gnd.n6359 gnd.n6358 19.3944
R9643 gnd.n6358 gnd.n844 19.3944
R9644 gnd.n6352 gnd.n844 19.3944
R9645 gnd.n6352 gnd.n6351 19.3944
R9646 gnd.n6351 gnd.n6350 19.3944
R9647 gnd.n6350 gnd.n852 19.3944
R9648 gnd.n6344 gnd.n852 19.3944
R9649 gnd.n6344 gnd.n6343 19.3944
R9650 gnd.n6343 gnd.n6342 19.3944
R9651 gnd.n6342 gnd.n860 19.3944
R9652 gnd.n6336 gnd.n860 19.3944
R9653 gnd.n6336 gnd.n6335 19.3944
R9654 gnd.n6335 gnd.n6334 19.3944
R9655 gnd.n6334 gnd.n868 19.3944
R9656 gnd.n6328 gnd.n868 19.3944
R9657 gnd.n6328 gnd.n6327 19.3944
R9658 gnd.n4379 gnd.n4376 19.3944
R9659 gnd.n4379 gnd.n3737 19.3944
R9660 gnd.n4406 gnd.n3737 19.3944
R9661 gnd.n4406 gnd.n3734 19.3944
R9662 gnd.n4411 gnd.n3734 19.3944
R9663 gnd.n4411 gnd.n3735 19.3944
R9664 gnd.n3735 gnd.n3712 19.3944
R9665 gnd.n4436 gnd.n3712 19.3944
R9666 gnd.n4436 gnd.n3709 19.3944
R9667 gnd.n4441 gnd.n3709 19.3944
R9668 gnd.n4441 gnd.n3710 19.3944
R9669 gnd.n3710 gnd.n3687 19.3944
R9670 gnd.n4476 gnd.n3687 19.3944
R9671 gnd.n4476 gnd.n3684 19.3944
R9672 gnd.n4481 gnd.n3684 19.3944
R9673 gnd.n4481 gnd.n3685 19.3944
R9674 gnd.n3685 gnd.n2917 19.3944
R9675 gnd.n5957 gnd.n2917 19.3944
R9676 gnd.n5957 gnd.n2918 19.3944
R9677 gnd.n5953 gnd.n2918 19.3944
R9678 gnd.n5953 gnd.n5952 19.3944
R9679 gnd.n5952 gnd.n5951 19.3944
R9680 gnd.n5951 gnd.n2924 19.3944
R9681 gnd.n5947 gnd.n2924 19.3944
R9682 gnd.n5947 gnd.n5946 19.3944
R9683 gnd.n5946 gnd.n5945 19.3944
R9684 gnd.n5945 gnd.n2929 19.3944
R9685 gnd.n5941 gnd.n2929 19.3944
R9686 gnd.n5941 gnd.n5940 19.3944
R9687 gnd.n5940 gnd.n5939 19.3944
R9688 gnd.n5939 gnd.n2934 19.3944
R9689 gnd.n5935 gnd.n2934 19.3944
R9690 gnd.n5935 gnd.n5934 19.3944
R9691 gnd.n5934 gnd.n5933 19.3944
R9692 gnd.n5933 gnd.n2939 19.3944
R9693 gnd.n5929 gnd.n2939 19.3944
R9694 gnd.n5929 gnd.n5928 19.3944
R9695 gnd.n5928 gnd.n5927 19.3944
R9696 gnd.n5927 gnd.n2944 19.3944
R9697 gnd.n5923 gnd.n2944 19.3944
R9698 gnd.n5923 gnd.n5922 19.3944
R9699 gnd.n5922 gnd.n5921 19.3944
R9700 gnd.n5921 gnd.n2949 19.3944
R9701 gnd.n5917 gnd.n2949 19.3944
R9702 gnd.n5917 gnd.n5916 19.3944
R9703 gnd.n5916 gnd.n5915 19.3944
R9704 gnd.n5915 gnd.n2954 19.3944
R9705 gnd.n5911 gnd.n2954 19.3944
R9706 gnd.n5911 gnd.n5910 19.3944
R9707 gnd.n5910 gnd.n5909 19.3944
R9708 gnd.n5909 gnd.n2959 19.3944
R9709 gnd.n5905 gnd.n2959 19.3944
R9710 gnd.n5905 gnd.n5904 19.3944
R9711 gnd.n5904 gnd.n5903 19.3944
R9712 gnd.n5903 gnd.n2964 19.3944
R9713 gnd.n5899 gnd.n2964 19.3944
R9714 gnd.n5899 gnd.n5898 19.3944
R9715 gnd.n5898 gnd.n5897 19.3944
R9716 gnd.n5897 gnd.n2969 19.3944
R9717 gnd.n5893 gnd.n2969 19.3944
R9718 gnd.n5893 gnd.n5892 19.3944
R9719 gnd.n5892 gnd.n5891 19.3944
R9720 gnd.n5891 gnd.n2974 19.3944
R9721 gnd.n5887 gnd.n2974 19.3944
R9722 gnd.n5887 gnd.n5886 19.3944
R9723 gnd.n5886 gnd.n5885 19.3944
R9724 gnd.n5885 gnd.n2979 19.3944
R9725 gnd.n5881 gnd.n2979 19.3944
R9726 gnd.n5881 gnd.n5880 19.3944
R9727 gnd.n5880 gnd.n5879 19.3944
R9728 gnd.n5879 gnd.n2984 19.3944
R9729 gnd.n5875 gnd.n2984 19.3944
R9730 gnd.n5875 gnd.n5874 19.3944
R9731 gnd.n5874 gnd.n5873 19.3944
R9732 gnd.n5873 gnd.n2989 19.3944
R9733 gnd.n5869 gnd.n2989 19.3944
R9734 gnd.n5869 gnd.n5868 19.3944
R9735 gnd.n5868 gnd.n5867 19.3944
R9736 gnd.n5867 gnd.n2994 19.3944
R9737 gnd.n5863 gnd.n2994 19.3944
R9738 gnd.n5863 gnd.n5862 19.3944
R9739 gnd.n5862 gnd.n5861 19.3944
R9740 gnd.n5058 gnd.n5055 19.3944
R9741 gnd.n5058 gnd.n5053 19.3944
R9742 gnd.n5064 gnd.n5053 19.3944
R9743 gnd.n5064 gnd.n5051 19.3944
R9744 gnd.n5069 gnd.n5051 19.3944
R9745 gnd.n5069 gnd.n5049 19.3944
R9746 gnd.n5075 gnd.n5049 19.3944
R9747 gnd.n5075 gnd.n5048 19.3944
R9748 gnd.n5084 gnd.n5048 19.3944
R9749 gnd.n5084 gnd.n5046 19.3944
R9750 gnd.n5090 gnd.n5046 19.3944
R9751 gnd.n5090 gnd.n5039 19.3944
R9752 gnd.n5103 gnd.n5039 19.3944
R9753 gnd.n5103 gnd.n5037 19.3944
R9754 gnd.n5109 gnd.n5037 19.3944
R9755 gnd.n5109 gnd.n5030 19.3944
R9756 gnd.n5122 gnd.n5030 19.3944
R9757 gnd.n5122 gnd.n5028 19.3944
R9758 gnd.n5128 gnd.n5028 19.3944
R9759 gnd.n5128 gnd.n5021 19.3944
R9760 gnd.n5141 gnd.n5021 19.3944
R9761 gnd.n5141 gnd.n5019 19.3944
R9762 gnd.n5148 gnd.n5019 19.3944
R9763 gnd.n5148 gnd.n5147 19.3944
R9764 gnd.n5161 gnd.n5000 19.3944
R9765 gnd.n5000 gnd.n4999 19.3944
R9766 gnd.n5168 gnd.n4999 19.3944
R9767 gnd.n1723 gnd.t156 18.8012
R9768 gnd.n1708 gnd.t8 18.8012
R9769 gnd.n1567 gnd.n1566 18.4825
R9770 gnd.n5480 gnd.n5388 18.4247
R9771 gnd.n6035 gnd.n6034 18.4247
R9772 gnd.n5158 gnd.n5157 18.2308
R9773 gnd.n6089 gnd.n6088 18.2308
R9774 gnd.n240 gnd.n182 18.2308
R9775 gnd.n3873 gnd.n3864 18.2308
R9776 gnd.t298 gnd.n1247 18.1639
R9777 gnd.n1853 gnd.n870 18.1639
R9778 gnd.n5964 gnd.n5963 17.9517
R9779 gnd.n5315 gnd.n5314 17.9517
R9780 gnd.n1275 gnd.t66 17.5266
R9781 gnd.n1674 gnd.t20 16.8893
R9782 gnd.n6160 gnd.t211 16.8893
R9783 gnd.n4993 gnd.t194 16.8893
R9784 gnd.n5510 gnd.n3254 16.6793
R9785 gnd.n7397 gnd.n7394 16.6793
R9786 gnd.n4068 gnd.n3934 16.6793
R9787 gnd.n2831 gnd.n2828 16.6793
R9788 gnd.n1502 gnd.t183 16.2519
R9789 gnd.n1202 gnd.t47 16.2519
R9790 gnd.n6149 gnd.n2587 15.9333
R9791 gnd.n6149 gnd.n2601 15.9333
R9792 gnd.n4374 gnd.n4373 15.9333
R9793 gnd.n4375 gnd.n4374 15.9333
R9794 gnd.n4381 gnd.n4375 15.9333
R9795 gnd.n4393 gnd.n4381 15.9333
R9796 gnd.n4392 gnd.n3739 15.9333
R9797 gnd.n4404 gnd.n3739 15.9333
R9798 gnd.n4404 gnd.n4403 15.9333
R9799 gnd.n4403 gnd.n3741 15.9333
R9800 gnd.n3741 gnd.n3729 15.9333
R9801 gnd.n4413 gnd.n3729 15.9333
R9802 gnd.n4413 gnd.n3730 15.9333
R9803 gnd.n3732 gnd.n3730 15.9333
R9804 gnd.n4423 gnd.n4422 15.9333
R9805 gnd.n4422 gnd.n3714 15.9333
R9806 gnd.n4434 gnd.n3714 15.9333
R9807 gnd.n4434 gnd.n4433 15.9333
R9808 gnd.n4433 gnd.n3716 15.9333
R9809 gnd.n3716 gnd.n3705 15.9333
R9810 gnd.n4443 gnd.n3705 15.9333
R9811 gnd.n4443 gnd.n3706 15.9333
R9812 gnd.n4453 gnd.n3698 15.9333
R9813 gnd.n4453 gnd.n4452 15.9333
R9814 gnd.n4452 gnd.n3689 15.9333
R9815 gnd.n4474 gnd.n3689 15.9333
R9816 gnd.n4474 gnd.n4473 15.9333
R9817 gnd.n4473 gnd.n3691 15.9333
R9818 gnd.n3691 gnd.n3680 15.9333
R9819 gnd.n4483 gnd.n3680 15.9333
R9820 gnd.n4483 gnd.n3681 15.9333
R9821 gnd.n4466 gnd.n2885 15.9333
R9822 gnd.n4495 gnd.n2911 15.9333
R9823 gnd.n4528 gnd.n3604 15.9333
R9824 gnd.n4539 gnd.n4538 15.9333
R9825 gnd.n4658 gnd.n3534 15.9333
R9826 gnd.n4677 gnd.n3511 15.9333
R9827 gnd.n3518 gnd.n3506 15.9333
R9828 gnd.n4717 gnd.n3489 15.9333
R9829 gnd.n4764 gnd.n4763 15.9333
R9830 gnd.n4772 gnd.n3476 15.9333
R9831 gnd.n4789 gnd.n4788 15.9333
R9832 gnd.n4849 gnd.n3444 15.9333
R9833 gnd.n4923 gnd.n4922 15.9333
R9834 gnd.n4937 gnd.n3386 15.9333
R9835 gnd.n4955 gnd.n3372 15.9333
R9836 gnd.n3305 gnd.n3267 15.9333
R9837 gnd.n5218 gnd.n5217 15.9333
R9838 gnd.n5217 gnd.n5215 15.9333
R9839 gnd.n5215 gnd.n5214 15.9333
R9840 gnd.n5214 gnd.n5213 15.9333
R9841 gnd.n5213 gnd.n3323 15.9333
R9842 gnd.n3331 gnd.n3323 15.9333
R9843 gnd.n3332 gnd.n3331 15.9333
R9844 gnd.n5207 gnd.n3332 15.9333
R9845 gnd.n5207 gnd.n5206 15.9333
R9846 gnd.n5204 gnd.n5203 15.9333
R9847 gnd.n5203 gnd.n5202 15.9333
R9848 gnd.n5202 gnd.n3335 15.9333
R9849 gnd.n3343 gnd.n3335 15.9333
R9850 gnd.n3344 gnd.n3343 15.9333
R9851 gnd.n5196 gnd.n3344 15.9333
R9852 gnd.n5196 gnd.n5195 15.9333
R9853 gnd.n5195 gnd.n5193 15.9333
R9854 gnd.n5192 gnd.n5191 15.9333
R9855 gnd.n5191 gnd.n3347 15.9333
R9856 gnd.n3355 gnd.n3347 15.9333
R9857 gnd.n3356 gnd.n3355 15.9333
R9858 gnd.n5185 gnd.n3356 15.9333
R9859 gnd.n5185 gnd.n5184 15.9333
R9860 gnd.n5184 gnd.n5182 15.9333
R9861 gnd.n5182 gnd.n5181 15.9333
R9862 gnd.n5180 gnd.n5174 15.9333
R9863 gnd.n5174 gnd.n3000 15.9333
R9864 gnd.n5859 gnd.n3000 15.9333
R9865 gnd.n5859 gnd.n5858 15.9333
R9866 gnd.n3011 gnd.n3002 15.9333
R9867 gnd.n5852 gnd.n3011 15.9333
R9868 gnd.n2191 gnd.n2189 15.6674
R9869 gnd.n2159 gnd.n2157 15.6674
R9870 gnd.n2127 gnd.n2125 15.6674
R9871 gnd.n2096 gnd.n2094 15.6674
R9872 gnd.n2064 gnd.n2062 15.6674
R9873 gnd.n2032 gnd.n2030 15.6674
R9874 gnd.n2000 gnd.n1998 15.6674
R9875 gnd.n1969 gnd.n1967 15.6674
R9876 gnd.n1493 gnd.t183 15.6146
R9877 gnd.t179 gnd.n958 15.6146
R9878 gnd.t273 gnd.n959 15.6146
R9879 gnd.t238 gnd.n4392 15.6146
R9880 gnd.n5181 gnd.t218 15.6146
R9881 gnd.n5562 gnd.n3233 15.3217
R9882 gnd.n7352 gnd.n7347 15.3217
R9883 gnd.n4120 gnd.n3913 15.3217
R9884 gnd.n2786 gnd.n2781 15.3217
R9885 gnd.n4569 gnd.n3589 15.296
R9886 gnd.n4588 gnd.n3580 15.296
R9887 gnd.n4548 gnd.t143 15.296
R9888 gnd.n4718 gnd.n4716 15.296
R9889 gnd.n4762 gnd.n3485 15.296
R9890 gnd.n4890 gnd.t125 15.296
R9891 gnd.n4829 gnd.n3409 15.296
R9892 gnd.n4920 gnd.n3396 15.296
R9893 gnd.n5235 gnd.n5234 15.0827
R9894 gnd.n2897 gnd.n2892 15.0481
R9895 gnd.n5245 gnd.n5244 15.0481
R9896 gnd.n1863 gnd.t153 14.9773
R9897 gnd.n6290 gnd.t187 14.9773
R9898 gnd.n3706 gnd.t134 14.9773
R9899 gnd.t316 gnd.n5204 14.9773
R9900 gnd.n7491 gnd.t175 14.9773
R9901 gnd.n5960 gnd.n5959 14.6587
R9902 gnd.n4629 gnd.n4628 14.6587
R9903 gnd.n3437 gnd.n3426 14.6587
R9904 gnd.n5226 gnd.n5225 14.6587
R9905 gnd.t137 gnd.n1001 14.34
R9906 gnd.n1941 gnd.t68 14.34
R9907 gnd.n4512 gnd.n3596 14.0214
R9908 gnd.n4546 gnd.n3565 14.0214
R9909 gnd.n4708 gnd.n4707 14.0214
R9910 gnd.n3475 gnd.n3468 14.0214
R9911 gnd.n4891 gnd.n3413 14.0214
R9912 gnd.n1649 gnd.t39 13.7027
R9913 gnd.n3538 gnd.t105 13.7027
R9914 gnd.n4797 gnd.t77 13.7027
R9915 gnd.n1359 gnd.n1358 13.5763
R9916 gnd.n2305 gnd.n915 13.5763
R9917 gnd.n1567 gnd.n1305 13.384
R9918 gnd.n4527 gnd.n3606 13.384
R9919 gnd.n3566 gnd.n3560 13.384
R9920 gnd.t144 gnd.n4616 13.384
R9921 gnd.n4868 gnd.t10 13.384
R9922 gnd.n4877 gnd.n3422 13.384
R9923 gnd.n3379 gnd.n3378 13.384
R9924 gnd.n2908 gnd.n2889 13.1884
R9925 gnd.n2903 gnd.n2902 13.1884
R9926 gnd.n2902 gnd.n2901 13.1884
R9927 gnd.n5238 gnd.n5233 13.1884
R9928 gnd.n5239 gnd.n5238 13.1884
R9929 gnd.n2904 gnd.n2891 13.146
R9930 gnd.n2900 gnd.n2891 13.146
R9931 gnd.n5237 gnd.n5236 13.146
R9932 gnd.n5237 gnd.n5232 13.146
R9933 gnd.n2192 gnd.n2188 12.8005
R9934 gnd.n2160 gnd.n2156 12.8005
R9935 gnd.n2128 gnd.n2124 12.8005
R9936 gnd.n2097 gnd.n2093 12.8005
R9937 gnd.n2065 gnd.n2061 12.8005
R9938 gnd.n2033 gnd.n2029 12.8005
R9939 gnd.n2001 gnd.n1997 12.8005
R9940 gnd.n1970 gnd.n1966 12.8005
R9941 gnd.n4503 gnd.n4502 12.7467
R9942 gnd.n4678 gnd.n4676 12.7467
R9943 gnd.n4787 gnd.n3455 12.7467
R9944 gnd.n3385 gnd.t198 12.7467
R9945 gnd.n1358 gnd.n1353 12.4126
R9946 gnd.n2308 gnd.n2305 12.4126
R9947 gnd.n6027 gnd.n5964 12.1761
R9948 gnd.n5314 gnd.n5313 12.1761
R9949 gnd.n4599 gnd.n3571 12.1094
R9950 gnd.n4898 gnd.n3407 12.1094
R9951 gnd.n4938 gnd.n3383 12.1094
R9952 gnd.t267 gnd.n3310 12.1094
R9953 gnd.n2196 gnd.n2195 12.0247
R9954 gnd.n2164 gnd.n2163 12.0247
R9955 gnd.n2132 gnd.n2131 12.0247
R9956 gnd.n2101 gnd.n2100 12.0247
R9957 gnd.n2069 gnd.n2068 12.0247
R9958 gnd.n2037 gnd.n2036 12.0247
R9959 gnd.n2005 gnd.n2004 12.0247
R9960 gnd.n1974 gnd.n1973 12.0247
R9961 gnd.n6185 gnd.t54 11.7908
R9962 gnd.n5825 gnd.t81 11.7908
R9963 gnd.n6084 gnd.n2690 11.4721
R9964 gnd.n4638 gnd.t291 11.4721
R9965 gnd.n4636 gnd.n3547 11.4721
R9966 gnd.n4668 gnd.n4667 11.4721
R9967 gnd.n4815 gnd.n3450 11.4721
R9968 gnd.n4807 gnd.n3436 11.4721
R9969 gnd.n4859 gnd.t92 11.4721
R9970 gnd.n5317 gnd.n3305 11.4721
R9971 gnd.n5850 gnd.n3012 11.4721
R9972 gnd.n2199 gnd.n2186 11.249
R9973 gnd.n2167 gnd.n2154 11.249
R9974 gnd.n2135 gnd.n2122 11.249
R9975 gnd.n2104 gnd.n2091 11.249
R9976 gnd.n2072 gnd.n2059 11.249
R9977 gnd.n2040 gnd.n2027 11.249
R9978 gnd.n2008 gnd.n1995 11.249
R9979 gnd.n1977 gnd.n1964 11.249
R9980 gnd.n1637 gnd.t39 11.1535
R9981 gnd.n4196 gnd.t41 11.1535
R9982 gnd.n6209 gnd.t56 11.1535
R9983 gnd.n3732 gnd.t304 11.1535
R9984 gnd.n4615 gnd.t89 11.1535
R9985 gnd.t102 gnd.n4869 11.1535
R9986 gnd.t312 gnd.n5192 11.1535
R9987 gnd.n5801 gnd.t6 11.1535
R9988 gnd.n5756 gnd.t109 11.1535
R9989 gnd.n6296 gnd.n2366 10.8348
R9990 gnd.n4167 gnd.n4166 10.8348
R9991 gnd.n6290 gnd.n2377 10.8348
R9992 gnd.n4160 gnd.n2386 10.8348
R9993 gnd.n6284 gnd.n2389 10.8348
R9994 gnd.n4154 gnd.n2397 10.8348
R9995 gnd.n6278 gnd.n2400 10.8348
R9996 gnd.n4148 gnd.n2407 10.8348
R9997 gnd.n6272 gnd.n2410 10.8348
R9998 gnd.n6266 gnd.n2421 10.8348
R9999 gnd.n4197 gnd.n4196 10.8348
R10000 gnd.n6260 gnd.n2430 10.8348
R10001 gnd.n4205 gnd.n2438 10.8348
R10002 gnd.n6254 gnd.n2441 10.8348
R10003 gnd.n4211 gnd.n2448 10.8348
R10004 gnd.n6248 gnd.n2451 10.8348
R10005 gnd.n6241 gnd.n2460 10.8348
R10006 gnd.n4265 gnd.n4264 10.8348
R10007 gnd.n6235 gnd.n2469 10.8348
R10008 gnd.n4227 gnd.n2474 10.8348
R10009 gnd.n4242 gnd.n2483 10.8348
R10010 gnd.n6222 gnd.n2486 10.8348
R10011 gnd.n4251 gnd.n2491 10.8348
R10012 gnd.n6215 gnd.n2494 10.8348
R10013 gnd.n4283 gnd.n4282 10.8348
R10014 gnd.n6209 gnd.n2503 10.8348
R10015 gnd.n4291 gnd.n2511 10.8348
R10016 gnd.n4331 gnd.n2520 10.8348
R10017 gnd.n6197 gnd.n2523 10.8348
R10018 gnd.n4298 gnd.n2531 10.8348
R10019 gnd.n6191 gnd.n2534 10.8348
R10020 gnd.n4303 gnd.n4302 10.8348
R10021 gnd.n6185 gnd.n2543 10.8348
R10022 gnd.n4308 gnd.n2551 10.8348
R10023 gnd.n6179 gnd.n2554 10.8348
R10024 gnd.n4314 gnd.n2561 10.8348
R10025 gnd.n6173 gnd.n2564 10.8348
R10026 gnd.n6160 gnd.n2571 10.8348
R10027 gnd.n6167 gnd.n2574 10.8348
R10028 gnd.n4568 gnd.t252 10.8348
R10029 gnd.n4582 gnd.n4581 10.8348
R10030 gnd.n4581 gnd.n4580 10.8348
R10031 gnd.n4756 gnd.n4755 10.8348
R10032 gnd.n4755 gnd.n3482 10.8348
R10033 gnd.n4914 gnd.n4913 10.8348
R10034 gnd.n4913 gnd.n3393 10.8348
R10035 gnd.n5844 gnd.n5843 10.8348
R10036 gnd.n4993 gnd.n3023 10.8348
R10037 gnd.n5837 gnd.n3032 10.8348
R10038 gnd.n5572 gnd.n3035 10.8348
R10039 gnd.n5831 gnd.n3044 10.8348
R10040 gnd.n5580 gnd.n3047 10.8348
R10041 gnd.n5825 gnd.n3055 10.8348
R10042 gnd.n5601 gnd.n5600 10.8348
R10043 gnd.n5819 gnd.n3064 10.8348
R10044 gnd.n5589 gnd.n3067 10.8348
R10045 gnd.n5813 gnd.n3075 10.8348
R10046 gnd.n5645 gnd.n3078 10.8348
R10047 gnd.n5652 gnd.n3087 10.8348
R10048 gnd.n5801 gnd.n3095 10.8348
R10049 gnd.n5670 gnd.n3205 10.8348
R10050 gnd.n5795 gnd.n3104 10.8348
R10051 gnd.n5791 gnd.n3107 10.8348
R10052 gnd.n5790 gnd.n3113 10.8348
R10053 gnd.n3120 gnd.n3119 10.8348
R10054 gnd.n5777 gnd.n3123 10.8348
R10055 gnd.n5687 gnd.n3130 10.8348
R10056 gnd.n7541 gnd.n69 10.8348
R10057 gnd.n5770 gnd.n71 10.8348
R10058 gnd.n7533 gnd.n86 10.8348
R10059 gnd.n5703 gnd.n89 10.8348
R10060 gnd.n7527 gnd.n98 10.8348
R10061 gnd.n5712 gnd.n101 10.8348
R10062 gnd.n7521 gnd.n108 10.8348
R10063 gnd.n5756 gnd.n5755 10.8348
R10064 gnd.n7515 gnd.n117 10.8348
R10065 gnd.n7509 gnd.n128 10.8348
R10066 gnd.n5743 gnd.n131 10.8348
R10067 gnd.n7503 gnd.n138 10.8348
R10068 gnd.n5737 gnd.n141 10.8348
R10069 gnd.n7497 gnd.n149 10.8348
R10070 gnd.n5731 gnd.n152 10.8348
R10071 gnd.n7491 gnd.n159 10.8348
R10072 gnd.n7478 gnd.n176 10.8348
R10073 gnd.n7485 gnd.n168 10.8348
R10074 gnd.n3234 gnd.n3233 10.6672
R10075 gnd.n7355 gnd.n7352 10.6672
R10076 gnd.n3914 gnd.n3913 10.6672
R10077 gnd.n2789 gnd.n2786 10.6672
R10078 gnd.n5379 gnd.n3263 10.6151
R10079 gnd.n5379 gnd.n5378 10.6151
R10080 gnd.n5376 gnd.n5373 10.6151
R10081 gnd.n5373 gnd.n5372 10.6151
R10082 gnd.n5372 gnd.n5369 10.6151
R10083 gnd.n5369 gnd.n5368 10.6151
R10084 gnd.n5368 gnd.n5365 10.6151
R10085 gnd.n5365 gnd.n5364 10.6151
R10086 gnd.n5364 gnd.n5361 10.6151
R10087 gnd.n5361 gnd.n5360 10.6151
R10088 gnd.n5360 gnd.n5357 10.6151
R10089 gnd.n5357 gnd.n5356 10.6151
R10090 gnd.n5356 gnd.n5353 10.6151
R10091 gnd.n5353 gnd.n5352 10.6151
R10092 gnd.n5352 gnd.n5349 10.6151
R10093 gnd.n5349 gnd.n5348 10.6151
R10094 gnd.n5348 gnd.n5345 10.6151
R10095 gnd.n5345 gnd.n5344 10.6151
R10096 gnd.n5344 gnd.n5341 10.6151
R10097 gnd.n5341 gnd.n5340 10.6151
R10098 gnd.n5340 gnd.n5337 10.6151
R10099 gnd.n5337 gnd.n5336 10.6151
R10100 gnd.n5336 gnd.n5333 10.6151
R10101 gnd.n5333 gnd.n5332 10.6151
R10102 gnd.n5332 gnd.n5329 10.6151
R10103 gnd.n5329 gnd.n5328 10.6151
R10104 gnd.n5328 gnd.n5325 10.6151
R10105 gnd.n5325 gnd.n5324 10.6151
R10106 gnd.n5324 gnd.n5321 10.6151
R10107 gnd.n5321 gnd.n5320 10.6151
R10108 gnd.n4499 gnd.n4498 10.6151
R10109 gnd.n4500 gnd.n4499 10.6151
R10110 gnd.n4505 gnd.n4500 10.6151
R10111 gnd.n4506 gnd.n4505 10.6151
R10112 gnd.n4510 gnd.n4506 10.6151
R10113 gnd.n4510 gnd.n4509 10.6151
R10114 gnd.n4509 gnd.n4508 10.6151
R10115 gnd.n4508 gnd.n3587 10.6151
R10116 gnd.n4571 gnd.n3587 10.6151
R10117 gnd.n4572 gnd.n4571 10.6151
R10118 gnd.n4578 gnd.n4572 10.6151
R10119 gnd.n4578 gnd.n4577 10.6151
R10120 gnd.n4577 gnd.n4576 10.6151
R10121 gnd.n4576 gnd.n4573 10.6151
R10122 gnd.n4573 gnd.n3563 10.6151
R10123 gnd.n4608 gnd.n3563 10.6151
R10124 gnd.n4609 gnd.n4608 10.6151
R10125 gnd.n4613 gnd.n4609 10.6151
R10126 gnd.n4613 gnd.n4612 10.6151
R10127 gnd.n4612 gnd.n4611 10.6151
R10128 gnd.n4611 gnd.n4610 10.6151
R10129 gnd.n4610 gnd.n3537 10.6151
R10130 gnd.n4656 gnd.n3537 10.6151
R10131 gnd.n4656 gnd.n4655 10.6151
R10132 gnd.n4655 gnd.n4654 10.6151
R10133 gnd.n4654 gnd.n4653 10.6151
R10134 gnd.n4653 gnd.n3519 10.6151
R10135 gnd.n4680 gnd.n3519 10.6151
R10136 gnd.n4681 gnd.n4680 10.6151
R10137 gnd.n4683 gnd.n4681 10.6151
R10138 gnd.n4684 gnd.n4683 10.6151
R10139 gnd.n4685 gnd.n4684 10.6151
R10140 gnd.n4685 gnd.n3496 10.6151
R10141 gnd.n4720 gnd.n3496 10.6151
R10142 gnd.n4721 gnd.n4720 10.6151
R10143 gnd.n4723 gnd.n4721 10.6151
R10144 gnd.n4724 gnd.n4723 10.6151
R10145 gnd.n4726 gnd.n4724 10.6151
R10146 gnd.n4726 gnd.n4725 10.6151
R10147 gnd.n4725 gnd.n3466 10.6151
R10148 gnd.n4782 gnd.n3466 10.6151
R10149 gnd.n4783 gnd.n4782 10.6151
R10150 gnd.n4785 gnd.n4783 10.6151
R10151 gnd.n4785 gnd.n4784 10.6151
R10152 gnd.n4784 gnd.n3447 10.6151
R10153 gnd.n4817 gnd.n3447 10.6151
R10154 gnd.n4818 gnd.n4817 10.6151
R10155 gnd.n4847 gnd.n4818 10.6151
R10156 gnd.n4847 gnd.n4846 10.6151
R10157 gnd.n4846 gnd.n4845 10.6151
R10158 gnd.n4845 gnd.n4842 10.6151
R10159 gnd.n4842 gnd.n4841 10.6151
R10160 gnd.n4841 gnd.n4840 10.6151
R10161 gnd.n4840 gnd.n4839 10.6151
R10162 gnd.n4839 gnd.n4838 10.6151
R10163 gnd.n4838 gnd.n4835 10.6151
R10164 gnd.n4835 gnd.n4834 10.6151
R10165 gnd.n4834 gnd.n4832 10.6151
R10166 gnd.n4832 gnd.n4831 10.6151
R10167 gnd.n4831 gnd.n4826 10.6151
R10168 gnd.n4826 gnd.n4825 10.6151
R10169 gnd.n4825 gnd.n4823 10.6151
R10170 gnd.n4823 gnd.n4822 10.6151
R10171 gnd.n4822 gnd.n4819 10.6151
R10172 gnd.n4819 gnd.n3374 10.6151
R10173 gnd.n4947 gnd.n3374 10.6151
R10174 gnd.n4948 gnd.n4947 10.6151
R10175 gnd.n4951 gnd.n4948 10.6151
R10176 gnd.n4951 gnd.n4950 10.6151
R10177 gnd.n4950 gnd.n4949 10.6151
R10178 gnd.n4949 gnd.n3302 10.6151
R10179 gnd.n3611 gnd.n2850 10.6151
R10180 gnd.n3614 gnd.n3611 10.6151
R10181 gnd.n3619 gnd.n3616 10.6151
R10182 gnd.n3620 gnd.n3619 10.6151
R10183 gnd.n3623 gnd.n3620 10.6151
R10184 gnd.n3624 gnd.n3623 10.6151
R10185 gnd.n3627 gnd.n3624 10.6151
R10186 gnd.n3628 gnd.n3627 10.6151
R10187 gnd.n3631 gnd.n3628 10.6151
R10188 gnd.n3632 gnd.n3631 10.6151
R10189 gnd.n3635 gnd.n3632 10.6151
R10190 gnd.n3636 gnd.n3635 10.6151
R10191 gnd.n3639 gnd.n3636 10.6151
R10192 gnd.n3640 gnd.n3639 10.6151
R10193 gnd.n3643 gnd.n3640 10.6151
R10194 gnd.n3644 gnd.n3643 10.6151
R10195 gnd.n3647 gnd.n3644 10.6151
R10196 gnd.n3648 gnd.n3647 10.6151
R10197 gnd.n3651 gnd.n3648 10.6151
R10198 gnd.n3652 gnd.n3651 10.6151
R10199 gnd.n3655 gnd.n3652 10.6151
R10200 gnd.n3656 gnd.n3655 10.6151
R10201 gnd.n3659 gnd.n3656 10.6151
R10202 gnd.n3660 gnd.n3659 10.6151
R10203 gnd.n3663 gnd.n3660 10.6151
R10204 gnd.n3664 gnd.n3663 10.6151
R10205 gnd.n3667 gnd.n3664 10.6151
R10206 gnd.n3668 gnd.n3667 10.6151
R10207 gnd.n3671 gnd.n3668 10.6151
R10208 gnd.n3672 gnd.n3671 10.6151
R10209 gnd.n6027 gnd.n6026 10.6151
R10210 gnd.n6026 gnd.n6025 10.6151
R10211 gnd.n6025 gnd.n6024 10.6151
R10212 gnd.n6024 gnd.n6022 10.6151
R10213 gnd.n6022 gnd.n6019 10.6151
R10214 gnd.n6019 gnd.n6018 10.6151
R10215 gnd.n6018 gnd.n6015 10.6151
R10216 gnd.n6015 gnd.n6014 10.6151
R10217 gnd.n6014 gnd.n6011 10.6151
R10218 gnd.n6011 gnd.n6010 10.6151
R10219 gnd.n6010 gnd.n6007 10.6151
R10220 gnd.n6007 gnd.n6006 10.6151
R10221 gnd.n6006 gnd.n6003 10.6151
R10222 gnd.n6003 gnd.n6002 10.6151
R10223 gnd.n6002 gnd.n5999 10.6151
R10224 gnd.n5999 gnd.n5998 10.6151
R10225 gnd.n5998 gnd.n5995 10.6151
R10226 gnd.n5995 gnd.n5994 10.6151
R10227 gnd.n5994 gnd.n5991 10.6151
R10228 gnd.n5991 gnd.n5990 10.6151
R10229 gnd.n5990 gnd.n5987 10.6151
R10230 gnd.n5987 gnd.n5986 10.6151
R10231 gnd.n5986 gnd.n5983 10.6151
R10232 gnd.n5983 gnd.n5982 10.6151
R10233 gnd.n5982 gnd.n5979 10.6151
R10234 gnd.n5979 gnd.n5978 10.6151
R10235 gnd.n5978 gnd.n5975 10.6151
R10236 gnd.n5975 gnd.n5974 10.6151
R10237 gnd.n5971 gnd.n5970 10.6151
R10238 gnd.n5970 gnd.n2851 10.6151
R10239 gnd.n5313 gnd.n5312 10.6151
R10240 gnd.n5312 gnd.n5309 10.6151
R10241 gnd.n5309 gnd.n5308 10.6151
R10242 gnd.n5308 gnd.n5305 10.6151
R10243 gnd.n5305 gnd.n5304 10.6151
R10244 gnd.n5304 gnd.n5301 10.6151
R10245 gnd.n5301 gnd.n5300 10.6151
R10246 gnd.n5300 gnd.n5297 10.6151
R10247 gnd.n5297 gnd.n5296 10.6151
R10248 gnd.n5296 gnd.n5293 10.6151
R10249 gnd.n5293 gnd.n5292 10.6151
R10250 gnd.n5292 gnd.n5289 10.6151
R10251 gnd.n5289 gnd.n5288 10.6151
R10252 gnd.n5288 gnd.n5285 10.6151
R10253 gnd.n5285 gnd.n5284 10.6151
R10254 gnd.n5284 gnd.n5281 10.6151
R10255 gnd.n5281 gnd.n5280 10.6151
R10256 gnd.n5280 gnd.n5277 10.6151
R10257 gnd.n5277 gnd.n5276 10.6151
R10258 gnd.n5276 gnd.n5273 10.6151
R10259 gnd.n5273 gnd.n5272 10.6151
R10260 gnd.n5272 gnd.n5269 10.6151
R10261 gnd.n5269 gnd.n5268 10.6151
R10262 gnd.n5268 gnd.n5265 10.6151
R10263 gnd.n5265 gnd.n5264 10.6151
R10264 gnd.n5264 gnd.n5261 10.6151
R10265 gnd.n5261 gnd.n5260 10.6151
R10266 gnd.n5260 gnd.n5257 10.6151
R10267 gnd.n5255 gnd.n5252 10.6151
R10268 gnd.n5252 gnd.n3264 10.6151
R10269 gnd.n5963 gnd.n5962 10.6151
R10270 gnd.n5962 gnd.n2909 10.6151
R10271 gnd.n4515 gnd.n2909 10.6151
R10272 gnd.n4525 gnd.n4515 10.6151
R10273 gnd.n4525 gnd.n4524 10.6151
R10274 gnd.n4524 gnd.n4523 10.6151
R10275 gnd.n4523 gnd.n4516 10.6151
R10276 gnd.n4517 gnd.n4516 10.6151
R10277 gnd.n4517 gnd.n3582 10.6151
R10278 gnd.n4584 gnd.n3582 10.6151
R10279 gnd.n4585 gnd.n4584 10.6151
R10280 gnd.n4586 gnd.n4585 10.6151
R10281 gnd.n4586 gnd.n3569 10.6151
R10282 gnd.n4601 gnd.n3569 10.6151
R10283 gnd.n4602 gnd.n4601 10.6151
R10284 gnd.n4604 gnd.n4602 10.6151
R10285 gnd.n4604 gnd.n4603 10.6151
R10286 gnd.n4603 gnd.n3549 10.6151
R10287 gnd.n4632 gnd.n3549 10.6151
R10288 gnd.n4633 gnd.n4632 10.6151
R10289 gnd.n4634 gnd.n4633 10.6151
R10290 gnd.n4634 gnd.n3532 10.6151
R10291 gnd.n4660 gnd.n3532 10.6151
R10292 gnd.n4661 gnd.n4660 10.6151
R10293 gnd.n4665 gnd.n4661 10.6151
R10294 gnd.n4665 gnd.n4664 10.6151
R10295 gnd.n4664 gnd.n4663 10.6151
R10296 gnd.n4663 gnd.n3509 10.6151
R10297 gnd.n4700 gnd.n3509 10.6151
R10298 gnd.n4701 gnd.n4700 10.6151
R10299 gnd.n4705 gnd.n4701 10.6151
R10300 gnd.n4705 gnd.n4704 10.6151
R10301 gnd.n4704 gnd.n4703 10.6151
R10302 gnd.n4703 gnd.n3487 10.6151
R10303 gnd.n4758 gnd.n3487 10.6151
R10304 gnd.n4759 gnd.n4758 10.6151
R10305 gnd.n4760 gnd.n4759 10.6151
R10306 gnd.n4760 gnd.n3472 10.6151
R10307 gnd.n4775 gnd.n3472 10.6151
R10308 gnd.n4776 gnd.n4775 10.6151
R10309 gnd.n4778 gnd.n4776 10.6151
R10310 gnd.n4778 gnd.n4777 10.6151
R10311 gnd.n4777 gnd.n3453 10.6151
R10312 gnd.n4803 gnd.n3453 10.6151
R10313 gnd.n4804 gnd.n4803 10.6151
R10314 gnd.n4813 gnd.n4804 10.6151
R10315 gnd.n4813 gnd.n4812 10.6151
R10316 gnd.n4812 gnd.n4811 10.6151
R10317 gnd.n4811 gnd.n4810 10.6151
R10318 gnd.n4810 gnd.n4805 10.6151
R10319 gnd.n4805 gnd.n3424 10.6151
R10320 gnd.n4873 gnd.n3424 10.6151
R10321 gnd.n4874 gnd.n4873 10.6151
R10322 gnd.n4875 gnd.n4874 10.6151
R10323 gnd.n4875 gnd.n3411 10.6151
R10324 gnd.n4893 gnd.n3411 10.6151
R10325 gnd.n4894 gnd.n4893 10.6151
R10326 gnd.n4895 gnd.n4894 10.6151
R10327 gnd.n4895 gnd.n3398 10.6151
R10328 gnd.n4916 gnd.n3398 10.6151
R10329 gnd.n4917 gnd.n4916 10.6151
R10330 gnd.n4918 gnd.n4917 10.6151
R10331 gnd.n4918 gnd.n3381 10.6151
R10332 gnd.n4940 gnd.n3381 10.6151
R10333 gnd.n4941 gnd.n4940 10.6151
R10334 gnd.n4943 gnd.n4941 10.6151
R10335 gnd.n4943 gnd.n4942 10.6151
R10336 gnd.n4942 gnd.n3308 10.6151
R10337 gnd.n5229 gnd.n3308 10.6151
R10338 gnd.n5230 gnd.n5229 10.6151
R10339 gnd.n5315 gnd.n5230 10.6151
R10340 gnd.n1556 gnd.t141 10.5161
R10341 gnd.n1003 gnd.t137 10.5161
R10342 gnd.n1924 gnd.t68 10.5161
R10343 gnd.t95 gnd.n2457 10.5161
R10344 gnd.n4265 gnd.t43 10.5161
R10345 gnd.n6235 gnd.t43 10.5161
R10346 gnd.n6228 gnd.t17 10.5161
R10347 gnd.n4590 gnd.t87 10.5161
R10348 gnd.t115 gnd.n4827 10.5161
R10349 gnd.t61 gnd.n5782 10.5161
R10350 gnd.n5687 gnd.t33 10.5161
R10351 gnd.t33 gnd.n69 10.5161
R10352 gnd.n5769 gnd.t35 10.5161
R10353 gnd.n2200 gnd.n2184 10.4732
R10354 gnd.n2168 gnd.n2152 10.4732
R10355 gnd.n2136 gnd.n2120 10.4732
R10356 gnd.n2105 gnd.n2089 10.4732
R10357 gnd.n2073 gnd.n2057 10.4732
R10358 gnd.n2041 gnd.n2025 10.4732
R10359 gnd.n2009 gnd.n1993 10.4732
R10360 gnd.n1978 gnd.n1962 10.4732
R10361 gnd.n6298 gnd.n2363 10.1975
R10362 gnd.n4518 gnd.t289 10.1975
R10363 gnd.n3547 gnd.n3546 10.1975
R10364 gnd.n4668 gnd.n3527 10.1975
R10365 gnd.n4737 gnd.n3450 10.1975
R10366 gnd.n4808 gnd.n4807 10.1975
R10367 gnd.n7469 gnd.n184 10.1975
R10368 gnd.t153 gnd.n1020 9.87883
R10369 gnd.t73 gnd.n2418 9.87883
R10370 gnd.n6260 gnd.t41 9.87883
R10371 gnd.n4282 gnd.t56 9.87883
R10372 gnd.n6203 gnd.t69 9.87883
R10373 gnd.n5807 gnd.t13 9.87883
R10374 gnd.n3205 gnd.t6 9.87883
R10375 gnd.n7521 gnd.t109 9.87883
R10376 gnd.t25 gnd.n120 9.87883
R10377 gnd.n2204 gnd.n2203 9.69747
R10378 gnd.n2172 gnd.n2171 9.69747
R10379 gnd.n2140 gnd.n2139 9.69747
R10380 gnd.n2109 gnd.n2108 9.69747
R10381 gnd.n2077 gnd.n2076 9.69747
R10382 gnd.n2045 gnd.n2044 9.69747
R10383 gnd.n2013 gnd.n2012 9.69747
R10384 gnd.n1982 gnd.n1981 9.69747
R10385 gnd.n4519 gnd.n4518 9.56018
R10386 gnd.n4574 gnd.n3571 9.56018
R10387 gnd.n4641 gnd.t31 9.56018
R10388 gnd.n4689 gnd.n3498 9.56018
R10389 gnd.n4730 gnd.n4728 9.56018
R10390 gnd.n4738 gnd.t30 9.56018
R10391 gnd.n4898 gnd.n4897 9.56018
R10392 gnd.n2210 gnd.n2209 9.45567
R10393 gnd.n2178 gnd.n2177 9.45567
R10394 gnd.n2146 gnd.n2145 9.45567
R10395 gnd.n2115 gnd.n2114 9.45567
R10396 gnd.n2083 gnd.n2082 9.45567
R10397 gnd.n2051 gnd.n2050 9.45567
R10398 gnd.n2019 gnd.n2018 9.45567
R10399 gnd.n1988 gnd.n1987 9.45567
R10400 gnd.n5510 gnd.n3252 9.30959
R10401 gnd.n7394 gnd.n7326 9.30959
R10402 gnd.n4068 gnd.n3932 9.30959
R10403 gnd.n2828 gnd.n2760 9.30959
R10404 gnd.n2209 gnd.n2208 9.3005
R10405 gnd.n2182 gnd.n2181 9.3005
R10406 gnd.n2203 gnd.n2202 9.3005
R10407 gnd.n2201 gnd.n2200 9.3005
R10408 gnd.n2186 gnd.n2185 9.3005
R10409 gnd.n2195 gnd.n2194 9.3005
R10410 gnd.n2193 gnd.n2192 9.3005
R10411 gnd.n2177 gnd.n2176 9.3005
R10412 gnd.n2150 gnd.n2149 9.3005
R10413 gnd.n2171 gnd.n2170 9.3005
R10414 gnd.n2169 gnd.n2168 9.3005
R10415 gnd.n2154 gnd.n2153 9.3005
R10416 gnd.n2163 gnd.n2162 9.3005
R10417 gnd.n2161 gnd.n2160 9.3005
R10418 gnd.n2145 gnd.n2144 9.3005
R10419 gnd.n2118 gnd.n2117 9.3005
R10420 gnd.n2139 gnd.n2138 9.3005
R10421 gnd.n2137 gnd.n2136 9.3005
R10422 gnd.n2122 gnd.n2121 9.3005
R10423 gnd.n2131 gnd.n2130 9.3005
R10424 gnd.n2129 gnd.n2128 9.3005
R10425 gnd.n2114 gnd.n2113 9.3005
R10426 gnd.n2087 gnd.n2086 9.3005
R10427 gnd.n2108 gnd.n2107 9.3005
R10428 gnd.n2106 gnd.n2105 9.3005
R10429 gnd.n2091 gnd.n2090 9.3005
R10430 gnd.n2100 gnd.n2099 9.3005
R10431 gnd.n2098 gnd.n2097 9.3005
R10432 gnd.n2082 gnd.n2081 9.3005
R10433 gnd.n2055 gnd.n2054 9.3005
R10434 gnd.n2076 gnd.n2075 9.3005
R10435 gnd.n2074 gnd.n2073 9.3005
R10436 gnd.n2059 gnd.n2058 9.3005
R10437 gnd.n2068 gnd.n2067 9.3005
R10438 gnd.n2066 gnd.n2065 9.3005
R10439 gnd.n2050 gnd.n2049 9.3005
R10440 gnd.n2023 gnd.n2022 9.3005
R10441 gnd.n2044 gnd.n2043 9.3005
R10442 gnd.n2042 gnd.n2041 9.3005
R10443 gnd.n2027 gnd.n2026 9.3005
R10444 gnd.n2036 gnd.n2035 9.3005
R10445 gnd.n2034 gnd.n2033 9.3005
R10446 gnd.n2018 gnd.n2017 9.3005
R10447 gnd.n1991 gnd.n1990 9.3005
R10448 gnd.n2012 gnd.n2011 9.3005
R10449 gnd.n2010 gnd.n2009 9.3005
R10450 gnd.n1995 gnd.n1994 9.3005
R10451 gnd.n2004 gnd.n2003 9.3005
R10452 gnd.n2002 gnd.n2001 9.3005
R10453 gnd.n1987 gnd.n1986 9.3005
R10454 gnd.n1960 gnd.n1959 9.3005
R10455 gnd.n1981 gnd.n1980 9.3005
R10456 gnd.n1979 gnd.n1978 9.3005
R10457 gnd.n1964 gnd.n1963 9.3005
R10458 gnd.n1973 gnd.n1972 9.3005
R10459 gnd.n1971 gnd.n1970 9.3005
R10460 gnd.n2335 gnd.n2334 9.3005
R10461 gnd.n2333 gnd.n903 9.3005
R10462 gnd.n2332 gnd.n2331 9.3005
R10463 gnd.n2328 gnd.n904 9.3005
R10464 gnd.n2325 gnd.n905 9.3005
R10465 gnd.n2324 gnd.n906 9.3005
R10466 gnd.n2321 gnd.n907 9.3005
R10467 gnd.n2320 gnd.n908 9.3005
R10468 gnd.n2317 gnd.n909 9.3005
R10469 gnd.n2316 gnd.n910 9.3005
R10470 gnd.n2313 gnd.n911 9.3005
R10471 gnd.n2312 gnd.n912 9.3005
R10472 gnd.n2309 gnd.n913 9.3005
R10473 gnd.n2308 gnd.n914 9.3005
R10474 gnd.n2305 gnd.n2304 9.3005
R10475 gnd.n2303 gnd.n915 9.3005
R10476 gnd.n2336 gnd.n902 9.3005
R10477 gnd.n1575 gnd.n1574 9.3005
R10478 gnd.n1279 gnd.n1278 9.3005
R10479 gnd.n1602 gnd.n1601 9.3005
R10480 gnd.n1603 gnd.n1277 9.3005
R10481 gnd.n1607 gnd.n1604 9.3005
R10482 gnd.n1606 gnd.n1605 9.3005
R10483 gnd.n1251 gnd.n1250 9.3005
R10484 gnd.n1632 gnd.n1631 9.3005
R10485 gnd.n1633 gnd.n1249 9.3005
R10486 gnd.n1635 gnd.n1634 9.3005
R10487 gnd.n1229 gnd.n1228 9.3005
R10488 gnd.n1663 gnd.n1662 9.3005
R10489 gnd.n1664 gnd.n1227 9.3005
R10490 gnd.n1672 gnd.n1665 9.3005
R10491 gnd.n1671 gnd.n1666 9.3005
R10492 gnd.n1670 gnd.n1668 9.3005
R10493 gnd.n1667 gnd.n1176 9.3005
R10494 gnd.n1720 gnd.n1177 9.3005
R10495 gnd.n1719 gnd.n1178 9.3005
R10496 gnd.n1718 gnd.n1179 9.3005
R10497 gnd.n1198 gnd.n1180 9.3005
R10498 gnd.n1200 gnd.n1199 9.3005
R10499 gnd.n1098 gnd.n1097 9.3005
R10500 gnd.n1758 gnd.n1757 9.3005
R10501 gnd.n1759 gnd.n1096 9.3005
R10502 gnd.n1763 gnd.n1760 9.3005
R10503 gnd.n1762 gnd.n1761 9.3005
R10504 gnd.n1071 gnd.n1070 9.3005
R10505 gnd.n1798 gnd.n1797 9.3005
R10506 gnd.n1799 gnd.n1069 9.3005
R10507 gnd.n1803 gnd.n1800 9.3005
R10508 gnd.n1802 gnd.n1801 9.3005
R10509 gnd.n1045 gnd.n1044 9.3005
R10510 gnd.n1845 gnd.n1844 9.3005
R10511 gnd.n1846 gnd.n1043 9.3005
R10512 gnd.n1850 gnd.n1847 9.3005
R10513 gnd.n1849 gnd.n1848 9.3005
R10514 gnd.n1018 gnd.n1017 9.3005
R10515 gnd.n1885 gnd.n1884 9.3005
R10516 gnd.n1886 gnd.n1016 9.3005
R10517 gnd.n1890 gnd.n1887 9.3005
R10518 gnd.n1889 gnd.n1888 9.3005
R10519 gnd.n991 gnd.n990 9.3005
R10520 gnd.n1934 gnd.n1933 9.3005
R10521 gnd.n1935 gnd.n989 9.3005
R10522 gnd.n1939 gnd.n1936 9.3005
R10523 gnd.n1938 gnd.n1937 9.3005
R10524 gnd.n964 gnd.n963 9.3005
R10525 gnd.n2228 gnd.n2227 9.3005
R10526 gnd.n2229 gnd.n962 9.3005
R10527 gnd.n2235 gnd.n2230 9.3005
R10528 gnd.n2234 gnd.n2231 9.3005
R10529 gnd.n2233 gnd.n2232 9.3005
R10530 gnd.n1576 gnd.n1573 9.3005
R10531 gnd.n1358 gnd.n1317 9.3005
R10532 gnd.n1353 gnd.n1352 9.3005
R10533 gnd.n1351 gnd.n1318 9.3005
R10534 gnd.n1350 gnd.n1349 9.3005
R10535 gnd.n1346 gnd.n1319 9.3005
R10536 gnd.n1343 gnd.n1342 9.3005
R10537 gnd.n1341 gnd.n1320 9.3005
R10538 gnd.n1340 gnd.n1339 9.3005
R10539 gnd.n1336 gnd.n1321 9.3005
R10540 gnd.n1333 gnd.n1332 9.3005
R10541 gnd.n1331 gnd.n1322 9.3005
R10542 gnd.n1330 gnd.n1329 9.3005
R10543 gnd.n1326 gnd.n1324 9.3005
R10544 gnd.n1323 gnd.n1303 9.3005
R10545 gnd.n1570 gnd.n1302 9.3005
R10546 gnd.n1572 gnd.n1571 9.3005
R10547 gnd.n1360 gnd.n1359 9.3005
R10548 gnd.n1583 gnd.n1289 9.3005
R10549 gnd.n1590 gnd.n1290 9.3005
R10550 gnd.n1592 gnd.n1591 9.3005
R10551 gnd.n1593 gnd.n1270 9.3005
R10552 gnd.n1612 gnd.n1611 9.3005
R10553 gnd.n1614 gnd.n1262 9.3005
R10554 gnd.n1621 gnd.n1264 9.3005
R10555 gnd.n1622 gnd.n1259 9.3005
R10556 gnd.n1624 gnd.n1623 9.3005
R10557 gnd.n1260 gnd.n1245 9.3005
R10558 gnd.n1640 gnd.n1243 9.3005
R10559 gnd.n1644 gnd.n1643 9.3005
R10560 gnd.n1642 gnd.n1219 9.3005
R10561 gnd.n1679 gnd.n1218 9.3005
R10562 gnd.n1682 gnd.n1681 9.3005
R10563 gnd.n1215 gnd.n1214 9.3005
R10564 gnd.n1688 gnd.n1216 9.3005
R10565 gnd.n1690 gnd.n1689 9.3005
R10566 gnd.n1692 gnd.n1213 9.3005
R10567 gnd.n1695 gnd.n1694 9.3005
R10568 gnd.n1698 gnd.n1696 9.3005
R10569 gnd.n1700 gnd.n1699 9.3005
R10570 gnd.n1706 gnd.n1701 9.3005
R10571 gnd.n1705 gnd.n1704 9.3005
R10572 gnd.n1089 gnd.n1088 9.3005
R10573 gnd.n1772 gnd.n1771 9.3005
R10574 gnd.n1773 gnd.n1082 9.3005
R10575 gnd.n1781 gnd.n1081 9.3005
R10576 gnd.n1784 gnd.n1783 9.3005
R10577 gnd.n1786 gnd.n1785 9.3005
R10578 gnd.n1789 gnd.n1064 9.3005
R10579 gnd.n1787 gnd.n1062 9.3005
R10580 gnd.n1809 gnd.n1060 9.3005
R10581 gnd.n1811 gnd.n1810 9.3005
R10582 gnd.n1036 gnd.n1035 9.3005
R10583 gnd.n1859 gnd.n1858 9.3005
R10584 gnd.n1860 gnd.n1029 9.3005
R10585 gnd.n1868 gnd.n1028 9.3005
R10586 gnd.n1871 gnd.n1870 9.3005
R10587 gnd.n1873 gnd.n1872 9.3005
R10588 gnd.n1876 gnd.n1011 9.3005
R10589 gnd.n1874 gnd.n1009 9.3005
R10590 gnd.n1896 gnd.n1007 9.3005
R10591 gnd.n1898 gnd.n1897 9.3005
R10592 gnd.n982 gnd.n981 9.3005
R10593 gnd.n1948 gnd.n1947 9.3005
R10594 gnd.n1949 gnd.n975 9.3005
R10595 gnd.n1957 gnd.n974 9.3005
R10596 gnd.n2216 gnd.n2215 9.3005
R10597 gnd.n2218 gnd.n2217 9.3005
R10598 gnd.n2219 gnd.n955 9.3005
R10599 gnd.n2243 gnd.n2242 9.3005
R10600 gnd.n956 gnd.n918 9.3005
R10601 gnd.n1581 gnd.n1580 9.3005
R10602 gnd.n2299 gnd.n919 9.3005
R10603 gnd.n2298 gnd.n921 9.3005
R10604 gnd.n2295 gnd.n922 9.3005
R10605 gnd.n2294 gnd.n923 9.3005
R10606 gnd.n2291 gnd.n924 9.3005
R10607 gnd.n2290 gnd.n925 9.3005
R10608 gnd.n2287 gnd.n926 9.3005
R10609 gnd.n2286 gnd.n927 9.3005
R10610 gnd.n2283 gnd.n928 9.3005
R10611 gnd.n2282 gnd.n929 9.3005
R10612 gnd.n2279 gnd.n930 9.3005
R10613 gnd.n2278 gnd.n931 9.3005
R10614 gnd.n2275 gnd.n932 9.3005
R10615 gnd.n2274 gnd.n933 9.3005
R10616 gnd.n2271 gnd.n934 9.3005
R10617 gnd.n2270 gnd.n935 9.3005
R10618 gnd.n2267 gnd.n936 9.3005
R10619 gnd.n2266 gnd.n937 9.3005
R10620 gnd.n2263 gnd.n938 9.3005
R10621 gnd.n2262 gnd.n939 9.3005
R10622 gnd.n2259 gnd.n940 9.3005
R10623 gnd.n2258 gnd.n941 9.3005
R10624 gnd.n2255 gnd.n945 9.3005
R10625 gnd.n2254 gnd.n946 9.3005
R10626 gnd.n2251 gnd.n947 9.3005
R10627 gnd.n2250 gnd.n948 9.3005
R10628 gnd.n2301 gnd.n2300 9.3005
R10629 gnd.n1750 gnd.n1734 9.3005
R10630 gnd.n1749 gnd.n1735 9.3005
R10631 gnd.n1748 gnd.n1736 9.3005
R10632 gnd.n1746 gnd.n1737 9.3005
R10633 gnd.n1745 gnd.n1738 9.3005
R10634 gnd.n1743 gnd.n1739 9.3005
R10635 gnd.n1742 gnd.n1740 9.3005
R10636 gnd.n1052 gnd.n1051 9.3005
R10637 gnd.n1819 gnd.n1818 9.3005
R10638 gnd.n1820 gnd.n1050 9.3005
R10639 gnd.n1837 gnd.n1821 9.3005
R10640 gnd.n1836 gnd.n1822 9.3005
R10641 gnd.n1835 gnd.n1823 9.3005
R10642 gnd.n1833 gnd.n1824 9.3005
R10643 gnd.n1832 gnd.n1825 9.3005
R10644 gnd.n1830 gnd.n1826 9.3005
R10645 gnd.n1829 gnd.n1827 9.3005
R10646 gnd.n998 gnd.n997 9.3005
R10647 gnd.n1906 gnd.n1905 9.3005
R10648 gnd.n1907 gnd.n996 9.3005
R10649 gnd.n1928 gnd.n1908 9.3005
R10650 gnd.n1927 gnd.n1909 9.3005
R10651 gnd.n1926 gnd.n1910 9.3005
R10652 gnd.n1923 gnd.n1911 9.3005
R10653 gnd.n1922 gnd.n1912 9.3005
R10654 gnd.n1920 gnd.n1913 9.3005
R10655 gnd.n1919 gnd.n1914 9.3005
R10656 gnd.n1917 gnd.n1916 9.3005
R10657 gnd.n1915 gnd.n950 9.3005
R10658 gnd.n1491 gnd.n1490 9.3005
R10659 gnd.n1381 gnd.n1380 9.3005
R10660 gnd.n1505 gnd.n1504 9.3005
R10661 gnd.n1506 gnd.n1379 9.3005
R10662 gnd.n1508 gnd.n1507 9.3005
R10663 gnd.n1369 gnd.n1368 9.3005
R10664 gnd.n1521 gnd.n1520 9.3005
R10665 gnd.n1522 gnd.n1367 9.3005
R10666 gnd.n1554 gnd.n1523 9.3005
R10667 gnd.n1553 gnd.n1524 9.3005
R10668 gnd.n1552 gnd.n1525 9.3005
R10669 gnd.n1551 gnd.n1526 9.3005
R10670 gnd.n1548 gnd.n1527 9.3005
R10671 gnd.n1547 gnd.n1528 9.3005
R10672 gnd.n1546 gnd.n1529 9.3005
R10673 gnd.n1544 gnd.n1530 9.3005
R10674 gnd.n1543 gnd.n1531 9.3005
R10675 gnd.n1540 gnd.n1532 9.3005
R10676 gnd.n1539 gnd.n1533 9.3005
R10677 gnd.n1538 gnd.n1534 9.3005
R10678 gnd.n1536 gnd.n1535 9.3005
R10679 gnd.n1235 gnd.n1234 9.3005
R10680 gnd.n1652 gnd.n1651 9.3005
R10681 gnd.n1653 gnd.n1233 9.3005
R10682 gnd.n1657 gnd.n1654 9.3005
R10683 gnd.n1656 gnd.n1655 9.3005
R10684 gnd.n1157 gnd.n1156 9.3005
R10685 gnd.n1732 gnd.n1731 9.3005
R10686 gnd.n1489 gnd.n1390 9.3005
R10687 gnd.n1392 gnd.n1391 9.3005
R10688 gnd.n1436 gnd.n1434 9.3005
R10689 gnd.n1437 gnd.n1433 9.3005
R10690 gnd.n1440 gnd.n1429 9.3005
R10691 gnd.n1441 gnd.n1428 9.3005
R10692 gnd.n1444 gnd.n1427 9.3005
R10693 gnd.n1445 gnd.n1426 9.3005
R10694 gnd.n1448 gnd.n1425 9.3005
R10695 gnd.n1449 gnd.n1424 9.3005
R10696 gnd.n1452 gnd.n1423 9.3005
R10697 gnd.n1453 gnd.n1422 9.3005
R10698 gnd.n1456 gnd.n1421 9.3005
R10699 gnd.n1457 gnd.n1420 9.3005
R10700 gnd.n1460 gnd.n1419 9.3005
R10701 gnd.n1461 gnd.n1418 9.3005
R10702 gnd.n1464 gnd.n1417 9.3005
R10703 gnd.n1465 gnd.n1416 9.3005
R10704 gnd.n1468 gnd.n1415 9.3005
R10705 gnd.n1469 gnd.n1414 9.3005
R10706 gnd.n1472 gnd.n1413 9.3005
R10707 gnd.n1473 gnd.n1412 9.3005
R10708 gnd.n1476 gnd.n1411 9.3005
R10709 gnd.n1478 gnd.n1410 9.3005
R10710 gnd.n1479 gnd.n1409 9.3005
R10711 gnd.n1480 gnd.n1408 9.3005
R10712 gnd.n1481 gnd.n1407 9.3005
R10713 gnd.n1488 gnd.n1487 9.3005
R10714 gnd.n1497 gnd.n1496 9.3005
R10715 gnd.n1498 gnd.n1384 9.3005
R10716 gnd.n1500 gnd.n1499 9.3005
R10717 gnd.n1375 gnd.n1374 9.3005
R10718 gnd.n1513 gnd.n1512 9.3005
R10719 gnd.n1514 gnd.n1373 9.3005
R10720 gnd.n1516 gnd.n1515 9.3005
R10721 gnd.n1362 gnd.n1361 9.3005
R10722 gnd.n1559 gnd.n1558 9.3005
R10723 gnd.n1560 gnd.n1316 9.3005
R10724 gnd.n1564 gnd.n1562 9.3005
R10725 gnd.n1563 gnd.n1295 9.3005
R10726 gnd.n1582 gnd.n1294 9.3005
R10727 gnd.n1585 gnd.n1584 9.3005
R10728 gnd.n1288 gnd.n1287 9.3005
R10729 gnd.n1596 gnd.n1594 9.3005
R10730 gnd.n1595 gnd.n1269 9.3005
R10731 gnd.n1613 gnd.n1268 9.3005
R10732 gnd.n1616 gnd.n1615 9.3005
R10733 gnd.n1263 gnd.n1258 9.3005
R10734 gnd.n1626 gnd.n1625 9.3005
R10735 gnd.n1261 gnd.n1241 9.3005
R10736 gnd.n1647 gnd.n1242 9.3005
R10737 gnd.n1646 gnd.n1645 9.3005
R10738 gnd.n1244 gnd.n1220 9.3005
R10739 gnd.n1678 gnd.n1677 9.3005
R10740 gnd.n1680 gnd.n1165 9.3005
R10741 gnd.n1727 gnd.n1166 9.3005
R10742 gnd.n1726 gnd.n1167 9.3005
R10743 gnd.n1725 gnd.n1168 9.3005
R10744 gnd.n1691 gnd.n1169 9.3005
R10745 gnd.n1693 gnd.n1187 9.3005
R10746 gnd.n1713 gnd.n1188 9.3005
R10747 gnd.n1712 gnd.n1189 9.3005
R10748 gnd.n1711 gnd.n1190 9.3005
R10749 gnd.n1702 gnd.n1191 9.3005
R10750 gnd.n1703 gnd.n1090 9.3005
R10751 gnd.n1769 gnd.n1768 9.3005
R10752 gnd.n1770 gnd.n1083 9.3005
R10753 gnd.n1780 gnd.n1779 9.3005
R10754 gnd.n1782 gnd.n1079 9.3005
R10755 gnd.n1792 gnd.n1080 9.3005
R10756 gnd.n1791 gnd.n1790 9.3005
R10757 gnd.n1788 gnd.n1058 9.3005
R10758 gnd.n1814 gnd.n1059 9.3005
R10759 gnd.n1813 gnd.n1812 9.3005
R10760 gnd.n1061 gnd.n1037 9.3005
R10761 gnd.n1856 gnd.n1855 9.3005
R10762 gnd.n1857 gnd.n1030 9.3005
R10763 gnd.n1867 gnd.n1866 9.3005
R10764 gnd.n1869 gnd.n1026 9.3005
R10765 gnd.n1879 gnd.n1027 9.3005
R10766 gnd.n1878 gnd.n1877 9.3005
R10767 gnd.n1875 gnd.n1005 9.3005
R10768 gnd.n1901 gnd.n1006 9.3005
R10769 gnd.n1900 gnd.n1899 9.3005
R10770 gnd.n1008 gnd.n983 9.3005
R10771 gnd.n1945 gnd.n1944 9.3005
R10772 gnd.n1946 gnd.n976 9.3005
R10773 gnd.n1956 gnd.n1955 9.3005
R10774 gnd.n2214 gnd.n972 9.3005
R10775 gnd.n2222 gnd.n973 9.3005
R10776 gnd.n2221 gnd.n2220 9.3005
R10777 gnd.n954 gnd.n953 9.3005
R10778 gnd.n2245 gnd.n2244 9.3005
R10779 gnd.n1386 gnd.n1385 9.3005
R10780 gnd.n6498 gnd.n6497 9.3005
R10781 gnd.n703 gnd.n702 9.3005
R10782 gnd.n6505 gnd.n6504 9.3005
R10783 gnd.n6506 gnd.n701 9.3005
R10784 gnd.n6508 gnd.n6507 9.3005
R10785 gnd.n697 gnd.n696 9.3005
R10786 gnd.n6515 gnd.n6514 9.3005
R10787 gnd.n6516 gnd.n695 9.3005
R10788 gnd.n6518 gnd.n6517 9.3005
R10789 gnd.n691 gnd.n690 9.3005
R10790 gnd.n6525 gnd.n6524 9.3005
R10791 gnd.n6526 gnd.n689 9.3005
R10792 gnd.n6528 gnd.n6527 9.3005
R10793 gnd.n685 gnd.n684 9.3005
R10794 gnd.n6535 gnd.n6534 9.3005
R10795 gnd.n6536 gnd.n683 9.3005
R10796 gnd.n6538 gnd.n6537 9.3005
R10797 gnd.n679 gnd.n678 9.3005
R10798 gnd.n6545 gnd.n6544 9.3005
R10799 gnd.n6546 gnd.n677 9.3005
R10800 gnd.n6548 gnd.n6547 9.3005
R10801 gnd.n673 gnd.n672 9.3005
R10802 gnd.n6555 gnd.n6554 9.3005
R10803 gnd.n6556 gnd.n671 9.3005
R10804 gnd.n6558 gnd.n6557 9.3005
R10805 gnd.n667 gnd.n666 9.3005
R10806 gnd.n6565 gnd.n6564 9.3005
R10807 gnd.n6566 gnd.n665 9.3005
R10808 gnd.n6568 gnd.n6567 9.3005
R10809 gnd.n661 gnd.n660 9.3005
R10810 gnd.n6575 gnd.n6574 9.3005
R10811 gnd.n6576 gnd.n659 9.3005
R10812 gnd.n6578 gnd.n6577 9.3005
R10813 gnd.n655 gnd.n654 9.3005
R10814 gnd.n6585 gnd.n6584 9.3005
R10815 gnd.n6586 gnd.n653 9.3005
R10816 gnd.n6588 gnd.n6587 9.3005
R10817 gnd.n649 gnd.n648 9.3005
R10818 gnd.n6595 gnd.n6594 9.3005
R10819 gnd.n6596 gnd.n647 9.3005
R10820 gnd.n6598 gnd.n6597 9.3005
R10821 gnd.n643 gnd.n642 9.3005
R10822 gnd.n6605 gnd.n6604 9.3005
R10823 gnd.n6606 gnd.n641 9.3005
R10824 gnd.n6608 gnd.n6607 9.3005
R10825 gnd.n637 gnd.n636 9.3005
R10826 gnd.n6615 gnd.n6614 9.3005
R10827 gnd.n6616 gnd.n635 9.3005
R10828 gnd.n6618 gnd.n6617 9.3005
R10829 gnd.n631 gnd.n630 9.3005
R10830 gnd.n6625 gnd.n6624 9.3005
R10831 gnd.n6626 gnd.n629 9.3005
R10832 gnd.n6628 gnd.n6627 9.3005
R10833 gnd.n625 gnd.n624 9.3005
R10834 gnd.n6635 gnd.n6634 9.3005
R10835 gnd.n6636 gnd.n623 9.3005
R10836 gnd.n6638 gnd.n6637 9.3005
R10837 gnd.n619 gnd.n618 9.3005
R10838 gnd.n6645 gnd.n6644 9.3005
R10839 gnd.n6646 gnd.n617 9.3005
R10840 gnd.n6648 gnd.n6647 9.3005
R10841 gnd.n613 gnd.n612 9.3005
R10842 gnd.n6655 gnd.n6654 9.3005
R10843 gnd.n6656 gnd.n611 9.3005
R10844 gnd.n6658 gnd.n6657 9.3005
R10845 gnd.n607 gnd.n606 9.3005
R10846 gnd.n6665 gnd.n6664 9.3005
R10847 gnd.n6666 gnd.n605 9.3005
R10848 gnd.n6668 gnd.n6667 9.3005
R10849 gnd.n601 gnd.n600 9.3005
R10850 gnd.n6675 gnd.n6674 9.3005
R10851 gnd.n6676 gnd.n599 9.3005
R10852 gnd.n6678 gnd.n6677 9.3005
R10853 gnd.n595 gnd.n594 9.3005
R10854 gnd.n6685 gnd.n6684 9.3005
R10855 gnd.n6686 gnd.n593 9.3005
R10856 gnd.n6688 gnd.n6687 9.3005
R10857 gnd.n589 gnd.n588 9.3005
R10858 gnd.n6695 gnd.n6694 9.3005
R10859 gnd.n6696 gnd.n587 9.3005
R10860 gnd.n6698 gnd.n6697 9.3005
R10861 gnd.n583 gnd.n582 9.3005
R10862 gnd.n6705 gnd.n6704 9.3005
R10863 gnd.n6706 gnd.n581 9.3005
R10864 gnd.n6708 gnd.n6707 9.3005
R10865 gnd.n577 gnd.n576 9.3005
R10866 gnd.n6715 gnd.n6714 9.3005
R10867 gnd.n6716 gnd.n575 9.3005
R10868 gnd.n6718 gnd.n6717 9.3005
R10869 gnd.n571 gnd.n570 9.3005
R10870 gnd.n6725 gnd.n6724 9.3005
R10871 gnd.n6726 gnd.n569 9.3005
R10872 gnd.n6728 gnd.n6727 9.3005
R10873 gnd.n565 gnd.n564 9.3005
R10874 gnd.n6735 gnd.n6734 9.3005
R10875 gnd.n6736 gnd.n563 9.3005
R10876 gnd.n6738 gnd.n6737 9.3005
R10877 gnd.n559 gnd.n558 9.3005
R10878 gnd.n6745 gnd.n6744 9.3005
R10879 gnd.n6746 gnd.n557 9.3005
R10880 gnd.n6748 gnd.n6747 9.3005
R10881 gnd.n553 gnd.n552 9.3005
R10882 gnd.n6755 gnd.n6754 9.3005
R10883 gnd.n6756 gnd.n551 9.3005
R10884 gnd.n6758 gnd.n6757 9.3005
R10885 gnd.n547 gnd.n546 9.3005
R10886 gnd.n6765 gnd.n6764 9.3005
R10887 gnd.n6766 gnd.n545 9.3005
R10888 gnd.n6768 gnd.n6767 9.3005
R10889 gnd.n541 gnd.n540 9.3005
R10890 gnd.n6775 gnd.n6774 9.3005
R10891 gnd.n6776 gnd.n539 9.3005
R10892 gnd.n6778 gnd.n6777 9.3005
R10893 gnd.n535 gnd.n534 9.3005
R10894 gnd.n6785 gnd.n6784 9.3005
R10895 gnd.n6786 gnd.n533 9.3005
R10896 gnd.n6788 gnd.n6787 9.3005
R10897 gnd.n529 gnd.n528 9.3005
R10898 gnd.n6795 gnd.n6794 9.3005
R10899 gnd.n6796 gnd.n527 9.3005
R10900 gnd.n6798 gnd.n6797 9.3005
R10901 gnd.n523 gnd.n522 9.3005
R10902 gnd.n6805 gnd.n6804 9.3005
R10903 gnd.n6806 gnd.n521 9.3005
R10904 gnd.n6808 gnd.n6807 9.3005
R10905 gnd.n517 gnd.n516 9.3005
R10906 gnd.n6815 gnd.n6814 9.3005
R10907 gnd.n6816 gnd.n515 9.3005
R10908 gnd.n6818 gnd.n6817 9.3005
R10909 gnd.n511 gnd.n510 9.3005
R10910 gnd.n6825 gnd.n6824 9.3005
R10911 gnd.n6826 gnd.n509 9.3005
R10912 gnd.n6828 gnd.n6827 9.3005
R10913 gnd.n505 gnd.n504 9.3005
R10914 gnd.n6835 gnd.n6834 9.3005
R10915 gnd.n6836 gnd.n503 9.3005
R10916 gnd.n6838 gnd.n6837 9.3005
R10917 gnd.n499 gnd.n498 9.3005
R10918 gnd.n6845 gnd.n6844 9.3005
R10919 gnd.n6846 gnd.n497 9.3005
R10920 gnd.n6848 gnd.n6847 9.3005
R10921 gnd.n493 gnd.n492 9.3005
R10922 gnd.n6855 gnd.n6854 9.3005
R10923 gnd.n6856 gnd.n491 9.3005
R10924 gnd.n6858 gnd.n6857 9.3005
R10925 gnd.n487 gnd.n486 9.3005
R10926 gnd.n6865 gnd.n6864 9.3005
R10927 gnd.n6866 gnd.n485 9.3005
R10928 gnd.n6868 gnd.n6867 9.3005
R10929 gnd.n481 gnd.n480 9.3005
R10930 gnd.n6875 gnd.n6874 9.3005
R10931 gnd.n6876 gnd.n479 9.3005
R10932 gnd.n6878 gnd.n6877 9.3005
R10933 gnd.n475 gnd.n474 9.3005
R10934 gnd.n6885 gnd.n6884 9.3005
R10935 gnd.n6886 gnd.n473 9.3005
R10936 gnd.n6888 gnd.n6887 9.3005
R10937 gnd.n469 gnd.n468 9.3005
R10938 gnd.n6895 gnd.n6894 9.3005
R10939 gnd.n6896 gnd.n467 9.3005
R10940 gnd.n6898 gnd.n6897 9.3005
R10941 gnd.n463 gnd.n462 9.3005
R10942 gnd.n6905 gnd.n6904 9.3005
R10943 gnd.n6906 gnd.n461 9.3005
R10944 gnd.n6908 gnd.n6907 9.3005
R10945 gnd.n457 gnd.n456 9.3005
R10946 gnd.n6915 gnd.n6914 9.3005
R10947 gnd.n6916 gnd.n455 9.3005
R10948 gnd.n6918 gnd.n6917 9.3005
R10949 gnd.n451 gnd.n450 9.3005
R10950 gnd.n6925 gnd.n6924 9.3005
R10951 gnd.n6926 gnd.n449 9.3005
R10952 gnd.n6928 gnd.n6927 9.3005
R10953 gnd.n445 gnd.n444 9.3005
R10954 gnd.n6935 gnd.n6934 9.3005
R10955 gnd.n6936 gnd.n443 9.3005
R10956 gnd.n6938 gnd.n6937 9.3005
R10957 gnd.n439 gnd.n438 9.3005
R10958 gnd.n6945 gnd.n6944 9.3005
R10959 gnd.n6946 gnd.n437 9.3005
R10960 gnd.n6948 gnd.n6947 9.3005
R10961 gnd.n433 gnd.n432 9.3005
R10962 gnd.n6955 gnd.n6954 9.3005
R10963 gnd.n6956 gnd.n431 9.3005
R10964 gnd.n6958 gnd.n6957 9.3005
R10965 gnd.n427 gnd.n426 9.3005
R10966 gnd.n6965 gnd.n6964 9.3005
R10967 gnd.n6966 gnd.n425 9.3005
R10968 gnd.n6968 gnd.n6967 9.3005
R10969 gnd.n421 gnd.n420 9.3005
R10970 gnd.n6975 gnd.n6974 9.3005
R10971 gnd.n6976 gnd.n419 9.3005
R10972 gnd.n6978 gnd.n6977 9.3005
R10973 gnd.n415 gnd.n414 9.3005
R10974 gnd.n6985 gnd.n6984 9.3005
R10975 gnd.n6986 gnd.n413 9.3005
R10976 gnd.n6988 gnd.n6987 9.3005
R10977 gnd.n409 gnd.n408 9.3005
R10978 gnd.n6995 gnd.n6994 9.3005
R10979 gnd.n6996 gnd.n407 9.3005
R10980 gnd.n6998 gnd.n6997 9.3005
R10981 gnd.n403 gnd.n402 9.3005
R10982 gnd.n7005 gnd.n7004 9.3005
R10983 gnd.n7006 gnd.n401 9.3005
R10984 gnd.n7009 gnd.n7008 9.3005
R10985 gnd.n7007 gnd.n397 9.3005
R10986 gnd.n7015 gnd.n396 9.3005
R10987 gnd.n7017 gnd.n7016 9.3005
R10988 gnd.n392 gnd.n391 9.3005
R10989 gnd.n7026 gnd.n7025 9.3005
R10990 gnd.n7027 gnd.n390 9.3005
R10991 gnd.n7029 gnd.n7028 9.3005
R10992 gnd.n386 gnd.n385 9.3005
R10993 gnd.n7036 gnd.n7035 9.3005
R10994 gnd.n7037 gnd.n384 9.3005
R10995 gnd.n7039 gnd.n7038 9.3005
R10996 gnd.n380 gnd.n379 9.3005
R10997 gnd.n7046 gnd.n7045 9.3005
R10998 gnd.n7047 gnd.n378 9.3005
R10999 gnd.n7049 gnd.n7048 9.3005
R11000 gnd.n374 gnd.n373 9.3005
R11001 gnd.n7056 gnd.n7055 9.3005
R11002 gnd.n7057 gnd.n372 9.3005
R11003 gnd.n7059 gnd.n7058 9.3005
R11004 gnd.n368 gnd.n367 9.3005
R11005 gnd.n7066 gnd.n7065 9.3005
R11006 gnd.n7067 gnd.n366 9.3005
R11007 gnd.n7069 gnd.n7068 9.3005
R11008 gnd.n362 gnd.n361 9.3005
R11009 gnd.n7076 gnd.n7075 9.3005
R11010 gnd.n7077 gnd.n360 9.3005
R11011 gnd.n7079 gnd.n7078 9.3005
R11012 gnd.n356 gnd.n355 9.3005
R11013 gnd.n7086 gnd.n7085 9.3005
R11014 gnd.n7087 gnd.n354 9.3005
R11015 gnd.n7089 gnd.n7088 9.3005
R11016 gnd.n350 gnd.n349 9.3005
R11017 gnd.n7096 gnd.n7095 9.3005
R11018 gnd.n7097 gnd.n348 9.3005
R11019 gnd.n7099 gnd.n7098 9.3005
R11020 gnd.n344 gnd.n343 9.3005
R11021 gnd.n7106 gnd.n7105 9.3005
R11022 gnd.n7107 gnd.n342 9.3005
R11023 gnd.n7109 gnd.n7108 9.3005
R11024 gnd.n338 gnd.n337 9.3005
R11025 gnd.n7116 gnd.n7115 9.3005
R11026 gnd.n7117 gnd.n336 9.3005
R11027 gnd.n7119 gnd.n7118 9.3005
R11028 gnd.n332 gnd.n331 9.3005
R11029 gnd.n7126 gnd.n7125 9.3005
R11030 gnd.n7127 gnd.n330 9.3005
R11031 gnd.n7129 gnd.n7128 9.3005
R11032 gnd.n326 gnd.n325 9.3005
R11033 gnd.n7136 gnd.n7135 9.3005
R11034 gnd.n7137 gnd.n324 9.3005
R11035 gnd.n7139 gnd.n7138 9.3005
R11036 gnd.n320 gnd.n319 9.3005
R11037 gnd.n7146 gnd.n7145 9.3005
R11038 gnd.n7147 gnd.n318 9.3005
R11039 gnd.n7149 gnd.n7148 9.3005
R11040 gnd.n314 gnd.n313 9.3005
R11041 gnd.n7156 gnd.n7155 9.3005
R11042 gnd.n7157 gnd.n312 9.3005
R11043 gnd.n7159 gnd.n7158 9.3005
R11044 gnd.n308 gnd.n307 9.3005
R11045 gnd.n7166 gnd.n7165 9.3005
R11046 gnd.n7167 gnd.n306 9.3005
R11047 gnd.n7169 gnd.n7168 9.3005
R11048 gnd.n302 gnd.n301 9.3005
R11049 gnd.n7176 gnd.n7175 9.3005
R11050 gnd.n7177 gnd.n300 9.3005
R11051 gnd.n7179 gnd.n7178 9.3005
R11052 gnd.n296 gnd.n295 9.3005
R11053 gnd.n7186 gnd.n7185 9.3005
R11054 gnd.n7187 gnd.n294 9.3005
R11055 gnd.n7189 gnd.n7188 9.3005
R11056 gnd.n290 gnd.n289 9.3005
R11057 gnd.n7196 gnd.n7195 9.3005
R11058 gnd.n7197 gnd.n288 9.3005
R11059 gnd.n7199 gnd.n7198 9.3005
R11060 gnd.n284 gnd.n283 9.3005
R11061 gnd.n7206 gnd.n7205 9.3005
R11062 gnd.n7207 gnd.n282 9.3005
R11063 gnd.n7209 gnd.n7208 9.3005
R11064 gnd.n278 gnd.n277 9.3005
R11065 gnd.n7216 gnd.n7215 9.3005
R11066 gnd.n7217 gnd.n276 9.3005
R11067 gnd.n7219 gnd.n7218 9.3005
R11068 gnd.n272 gnd.n271 9.3005
R11069 gnd.n7226 gnd.n7225 9.3005
R11070 gnd.n7227 gnd.n270 9.3005
R11071 gnd.n7230 gnd.n7229 9.3005
R11072 gnd.n7019 gnd.n7018 9.3005
R11073 gnd.n7545 gnd.n7544 9.3005
R11074 gnd.n7543 gnd.n65 9.3005
R11075 gnd.n5693 gnd.n67 9.3005
R11076 gnd.n5695 gnd.n5694 9.3005
R11077 gnd.n3201 gnd.n3200 9.3005
R11078 gnd.n5706 gnd.n5705 9.3005
R11079 gnd.n5707 gnd.n3199 9.3005
R11080 gnd.n5710 gnd.n5709 9.3005
R11081 gnd.n5708 gnd.n3192 9.3005
R11082 gnd.n5753 gnd.n3193 9.3005
R11083 gnd.n5752 gnd.n3194 9.3005
R11084 gnd.n5751 gnd.n3195 9.3005
R11085 gnd.n5720 gnd.n3196 9.3005
R11086 gnd.n5741 gnd.n5721 9.3005
R11087 gnd.n5740 gnd.n5722 9.3005
R11088 gnd.n5739 gnd.n5723 9.3005
R11089 gnd.n5726 gnd.n5724 9.3005
R11090 gnd.n5729 gnd.n5728 9.3005
R11091 gnd.n5727 gnd.n177 9.3005
R11092 gnd.n7476 gnd.n178 9.3005
R11093 gnd.n7475 gnd.n7474 9.3005
R11094 gnd.n204 gnd.n200 9.3005
R11095 gnd.n208 gnd.n207 9.3005
R11096 gnd.n209 gnd.n199 9.3005
R11097 gnd.n211 gnd.n210 9.3005
R11098 gnd.n214 gnd.n198 9.3005
R11099 gnd.n218 gnd.n217 9.3005
R11100 gnd.n219 gnd.n197 9.3005
R11101 gnd.n221 gnd.n220 9.3005
R11102 gnd.n224 gnd.n196 9.3005
R11103 gnd.n228 gnd.n227 9.3005
R11104 gnd.n229 gnd.n195 9.3005
R11105 gnd.n231 gnd.n230 9.3005
R11106 gnd.n234 gnd.n194 9.3005
R11107 gnd.n237 gnd.n236 9.3005
R11108 gnd.n238 gnd.n193 9.3005
R11109 gnd.n240 gnd.n239 9.3005
R11110 gnd.n182 gnd.n179 9.3005
R11111 gnd.n7473 gnd.n7472 9.3005
R11112 gnd.n202 gnd.n201 9.3005
R11113 gnd.n7290 gnd.n7287 9.3005
R11114 gnd.n7466 gnd.n7291 9.3005
R11115 gnd.n7465 gnd.n7292 9.3005
R11116 gnd.n7464 gnd.n7293 9.3005
R11117 gnd.n7461 gnd.n7294 9.3005
R11118 gnd.n7460 gnd.n7295 9.3005
R11119 gnd.n7457 gnd.n7296 9.3005
R11120 gnd.n7456 gnd.n7297 9.3005
R11121 gnd.n7453 gnd.n7298 9.3005
R11122 gnd.n7452 gnd.n7299 9.3005
R11123 gnd.n7449 gnd.n7300 9.3005
R11124 gnd.n7448 gnd.n7301 9.3005
R11125 gnd.n7445 gnd.n7302 9.3005
R11126 gnd.n7444 gnd.n7303 9.3005
R11127 gnd.n7441 gnd.n7304 9.3005
R11128 gnd.n7440 gnd.n7305 9.3005
R11129 gnd.n7437 gnd.n7306 9.3005
R11130 gnd.n7433 gnd.n7307 9.3005
R11131 gnd.n7430 gnd.n7308 9.3005
R11132 gnd.n7429 gnd.n7309 9.3005
R11133 gnd.n7426 gnd.n7310 9.3005
R11134 gnd.n7425 gnd.n7311 9.3005
R11135 gnd.n7422 gnd.n7312 9.3005
R11136 gnd.n7421 gnd.n7313 9.3005
R11137 gnd.n7418 gnd.n7314 9.3005
R11138 gnd.n7417 gnd.n7315 9.3005
R11139 gnd.n7414 gnd.n7316 9.3005
R11140 gnd.n7413 gnd.n7317 9.3005
R11141 gnd.n7410 gnd.n7318 9.3005
R11142 gnd.n7409 gnd.n7319 9.3005
R11143 gnd.n7406 gnd.n7320 9.3005
R11144 gnd.n7405 gnd.n7321 9.3005
R11145 gnd.n7402 gnd.n7322 9.3005
R11146 gnd.n7401 gnd.n7323 9.3005
R11147 gnd.n7398 gnd.n7324 9.3005
R11148 gnd.n7397 gnd.n7325 9.3005
R11149 gnd.n7394 gnd.n7393 9.3005
R11150 gnd.n7392 gnd.n7326 9.3005
R11151 gnd.n7391 gnd.n7390 9.3005
R11152 gnd.n7387 gnd.n7329 9.3005
R11153 gnd.n7384 gnd.n7330 9.3005
R11154 gnd.n7383 gnd.n7331 9.3005
R11155 gnd.n7380 gnd.n7332 9.3005
R11156 gnd.n7379 gnd.n7333 9.3005
R11157 gnd.n7376 gnd.n7334 9.3005
R11158 gnd.n7375 gnd.n7335 9.3005
R11159 gnd.n7372 gnd.n7336 9.3005
R11160 gnd.n7371 gnd.n7337 9.3005
R11161 gnd.n7368 gnd.n7338 9.3005
R11162 gnd.n7367 gnd.n7339 9.3005
R11163 gnd.n7364 gnd.n7340 9.3005
R11164 gnd.n7363 gnd.n7341 9.3005
R11165 gnd.n7360 gnd.n7342 9.3005
R11166 gnd.n7359 gnd.n7343 9.3005
R11167 gnd.n7356 gnd.n7344 9.3005
R11168 gnd.n7355 gnd.n7345 9.3005
R11169 gnd.n7352 gnd.n7351 9.3005
R11170 gnd.n7350 gnd.n7347 9.3005
R11171 gnd.n7289 gnd.n7288 9.3005
R11172 gnd.n5567 gnd.n3038 9.3005
R11173 gnd.n5835 gnd.n3039 9.3005
R11174 gnd.n5834 gnd.n3040 9.3005
R11175 gnd.n5833 gnd.n3041 9.3005
R11176 gnd.n3223 gnd.n3042 9.3005
R11177 gnd.n5823 gnd.n3059 9.3005
R11178 gnd.n5822 gnd.n3060 9.3005
R11179 gnd.n5821 gnd.n3061 9.3005
R11180 gnd.n5586 gnd.n3062 9.3005
R11181 gnd.n5811 gnd.n3080 9.3005
R11182 gnd.n5810 gnd.n3081 9.3005
R11183 gnd.n5809 gnd.n3082 9.3005
R11184 gnd.n5649 gnd.n3083 9.3005
R11185 gnd.n5799 gnd.n3099 9.3005
R11186 gnd.n5798 gnd.n3100 9.3005
R11187 gnd.n5797 gnd.n3101 9.3005
R11188 gnd.n3203 gnd.n3102 9.3005
R11189 gnd.n5679 gnd.n5678 9.3005
R11190 gnd.n5683 gnd.n5682 9.3005
R11191 gnd.n5684 gnd.n3132 9.3005
R11192 gnd.n5775 gnd.n3133 9.3005
R11193 gnd.n5774 gnd.n3134 9.3005
R11194 gnd.n5773 gnd.n3135 9.3005
R11195 gnd.n5772 gnd.n3136 9.3005
R11196 gnd.n5692 gnd.n92 9.3005
R11197 gnd.n7531 gnd.n93 9.3005
R11198 gnd.n7530 gnd.n94 9.3005
R11199 gnd.n7529 gnd.n95 9.3005
R11200 gnd.n3198 gnd.n96 9.3005
R11201 gnd.n7519 gnd.n112 9.3005
R11202 gnd.n7518 gnd.n113 9.3005
R11203 gnd.n7517 gnd.n114 9.3005
R11204 gnd.n5718 gnd.n115 9.3005
R11205 gnd.n7507 gnd.n133 9.3005
R11206 gnd.n7506 gnd.n134 9.3005
R11207 gnd.n7505 gnd.n135 9.3005
R11208 gnd.n5725 gnd.n136 9.3005
R11209 gnd.n7495 gnd.n154 9.3005
R11210 gnd.n7494 gnd.n155 9.3005
R11211 gnd.n7493 gnd.n156 9.3005
R11212 gnd.n173 gnd.n157 9.3005
R11213 gnd.n7483 gnd.n7482 9.3005
R11214 gnd.n5566 gnd.n5565 9.3005
R11215 gnd.n5568 gnd.n5567 9.3005
R11216 gnd.n5569 gnd.n3039 9.3005
R11217 gnd.n5570 gnd.n3040 9.3005
R11218 gnd.n3222 gnd.n3041 9.3005
R11219 gnd.n5582 gnd.n3223 9.3005
R11220 gnd.n5583 gnd.n3059 9.3005
R11221 gnd.n5584 gnd.n3060 9.3005
R11222 gnd.n5585 gnd.n3061 9.3005
R11223 gnd.n5587 gnd.n5586 9.3005
R11224 gnd.n3210 gnd.n3080 9.3005
R11225 gnd.n5647 gnd.n3081 9.3005
R11226 gnd.n5648 gnd.n3082 9.3005
R11227 gnd.n5650 gnd.n5649 9.3005
R11228 gnd.n3204 gnd.n3099 9.3005
R11229 gnd.n5672 gnd.n3100 9.3005
R11230 gnd.n5673 gnd.n3101 9.3005
R11231 gnd.n5674 gnd.n3203 9.3005
R11232 gnd.n5678 gnd.n5677 9.3005
R11233 gnd.n5683 gnd.n3202 9.3005
R11234 gnd.n5685 gnd.n5684 9.3005
R11235 gnd.n5686 gnd.n3133 9.3005
R11236 gnd.n5689 gnd.n3134 9.3005
R11237 gnd.n5690 gnd.n3135 9.3005
R11238 gnd.n5691 gnd.n3136 9.3005
R11239 gnd.n5699 gnd.n5692 9.3005
R11240 gnd.n5700 gnd.n93 9.3005
R11241 gnd.n5701 gnd.n94 9.3005
R11242 gnd.n3197 gnd.n95 9.3005
R11243 gnd.n5714 gnd.n3198 9.3005
R11244 gnd.n5715 gnd.n112 9.3005
R11245 gnd.n5716 gnd.n113 9.3005
R11246 gnd.n5717 gnd.n114 9.3005
R11247 gnd.n5747 gnd.n5718 9.3005
R11248 gnd.n5746 gnd.n133 9.3005
R11249 gnd.n5745 gnd.n134 9.3005
R11250 gnd.n5719 gnd.n135 9.3005
R11251 gnd.n5735 gnd.n5725 9.3005
R11252 gnd.n5734 gnd.n154 9.3005
R11253 gnd.n5733 gnd.n155 9.3005
R11254 gnd.n175 gnd.n156 9.3005
R11255 gnd.n7480 gnd.n173 9.3005
R11256 gnd.n7482 gnd.n7481 9.3005
R11257 gnd.n5566 gnd.n3227 9.3005
R11258 gnd.n3233 gnd.n3230 9.3005
R11259 gnd.n5553 gnd.n3234 9.3005
R11260 gnd.n5555 gnd.n5554 9.3005
R11261 gnd.n5552 gnd.n3236 9.3005
R11262 gnd.n5551 gnd.n5550 9.3005
R11263 gnd.n3238 gnd.n3237 9.3005
R11264 gnd.n5544 gnd.n5543 9.3005
R11265 gnd.n5542 gnd.n3240 9.3005
R11266 gnd.n5541 gnd.n5540 9.3005
R11267 gnd.n3242 gnd.n3241 9.3005
R11268 gnd.n5534 gnd.n5533 9.3005
R11269 gnd.n5532 gnd.n3244 9.3005
R11270 gnd.n5531 gnd.n5530 9.3005
R11271 gnd.n3246 gnd.n3245 9.3005
R11272 gnd.n5524 gnd.n5523 9.3005
R11273 gnd.n5522 gnd.n3248 9.3005
R11274 gnd.n5521 gnd.n5520 9.3005
R11275 gnd.n3250 gnd.n3249 9.3005
R11276 gnd.n5514 gnd.n5513 9.3005
R11277 gnd.n5512 gnd.n3252 9.3005
R11278 gnd.n3254 gnd.n3253 9.3005
R11279 gnd.n5502 gnd.n5501 9.3005
R11280 gnd.n5500 gnd.n3256 9.3005
R11281 gnd.n5499 gnd.n5498 9.3005
R11282 gnd.n3258 gnd.n3257 9.3005
R11283 gnd.n5492 gnd.n5491 9.3005
R11284 gnd.n5490 gnd.n3260 9.3005
R11285 gnd.n5489 gnd.n5488 9.3005
R11286 gnd.n3262 gnd.n3261 9.3005
R11287 gnd.n5480 gnd.n5479 9.3005
R11288 gnd.n5477 gnd.n5390 9.3005
R11289 gnd.n5476 gnd.n5475 9.3005
R11290 gnd.n5392 gnd.n5391 9.3005
R11291 gnd.n5469 gnd.n5468 9.3005
R11292 gnd.n5467 gnd.n5394 9.3005
R11293 gnd.n5466 gnd.n5465 9.3005
R11294 gnd.n5396 gnd.n5395 9.3005
R11295 gnd.n5459 gnd.n5455 9.3005
R11296 gnd.n5454 gnd.n5398 9.3005
R11297 gnd.n5453 gnd.n5452 9.3005
R11298 gnd.n5400 gnd.n5399 9.3005
R11299 gnd.n5446 gnd.n5445 9.3005
R11300 gnd.n5444 gnd.n5402 9.3005
R11301 gnd.n5443 gnd.n5442 9.3005
R11302 gnd.n5404 gnd.n5403 9.3005
R11303 gnd.n5436 gnd.n5435 9.3005
R11304 gnd.n5434 gnd.n5406 9.3005
R11305 gnd.n5433 gnd.n5432 9.3005
R11306 gnd.n5408 gnd.n5407 9.3005
R11307 gnd.n5426 gnd.n5425 9.3005
R11308 gnd.n5424 gnd.n5410 9.3005
R11309 gnd.n5423 gnd.n5422 9.3005
R11310 gnd.n5412 gnd.n5411 9.3005
R11311 gnd.n5416 gnd.n5415 9.3005
R11312 gnd.n5414 gnd.n5413 9.3005
R11313 gnd.n5511 gnd.n5510 9.3005
R11314 gnd.n5563 gnd.n5562 9.3005
R11315 gnd.n5840 gnd.n3028 9.3005
R11316 gnd.n5839 gnd.n3029 9.3005
R11317 gnd.n3049 gnd.n3030 9.3005
R11318 gnd.n5829 gnd.n3050 9.3005
R11319 gnd.n5828 gnd.n3051 9.3005
R11320 gnd.n5827 gnd.n3052 9.3005
R11321 gnd.n3069 gnd.n3053 9.3005
R11322 gnd.n5817 gnd.n3070 9.3005
R11323 gnd.n5816 gnd.n3071 9.3005
R11324 gnd.n5815 gnd.n3072 9.3005
R11325 gnd.n3089 gnd.n3073 9.3005
R11326 gnd.n5805 gnd.n3090 9.3005
R11327 gnd.n5804 gnd.n3091 9.3005
R11328 gnd.n5803 gnd.n3092 9.3005
R11329 gnd.n3093 gnd.n78 9.3005
R11330 gnd.n83 gnd.n77 9.3005
R11331 gnd.n7525 gnd.n103 9.3005
R11332 gnd.n7524 gnd.n104 9.3005
R11333 gnd.n7523 gnd.n105 9.3005
R11334 gnd.n122 gnd.n106 9.3005
R11335 gnd.n7513 gnd.n123 9.3005
R11336 gnd.n7512 gnd.n124 9.3005
R11337 gnd.n7511 gnd.n125 9.3005
R11338 gnd.n143 gnd.n126 9.3005
R11339 gnd.n7501 gnd.n144 9.3005
R11340 gnd.n7500 gnd.n145 9.3005
R11341 gnd.n7499 gnd.n146 9.3005
R11342 gnd.n163 gnd.n147 9.3005
R11343 gnd.n7489 gnd.n164 9.3005
R11344 gnd.n7488 gnd.n165 9.3005
R11345 gnd.n7487 gnd.n166 9.3005
R11346 gnd.n5841 gnd.n3027 9.3005
R11347 gnd.n7536 gnd.n7535 9.3005
R11348 gnd.n4276 gnd.n3787 9.3005
R11349 gnd.n4280 gnd.n4277 9.3005
R11350 gnd.n4279 gnd.n4278 9.3005
R11351 gnd.n3767 gnd.n3766 9.3005
R11352 gnd.n4335 gnd.n4334 9.3005
R11353 gnd.n4336 gnd.n3765 9.3005
R11354 gnd.n4338 gnd.n4337 9.3005
R11355 gnd.n3763 gnd.n3762 9.3005
R11356 gnd.n4343 gnd.n4342 9.3005
R11357 gnd.n4344 gnd.n3761 9.3005
R11358 gnd.n4346 gnd.n4345 9.3005
R11359 gnd.n3759 gnd.n3758 9.3005
R11360 gnd.n4351 gnd.n4350 9.3005
R11361 gnd.n4352 gnd.n3757 9.3005
R11362 gnd.n4354 gnd.n4353 9.3005
R11363 gnd.n3755 gnd.n3754 9.3005
R11364 gnd.n4359 gnd.n4358 9.3005
R11365 gnd.n4360 gnd.n3753 9.3005
R11366 gnd.n4362 gnd.n4361 9.3005
R11367 gnd.n3751 gnd.n3750 9.3005
R11368 gnd.n4368 gnd.n4367 9.3005
R11369 gnd.n4369 gnd.n3749 9.3005
R11370 gnd.n4371 gnd.n4370 9.3005
R11371 gnd.n3746 gnd.n3745 9.3005
R11372 gnd.n4396 gnd.n4395 9.3005
R11373 gnd.n4397 gnd.n3744 9.3005
R11374 gnd.n4401 gnd.n4398 9.3005
R11375 gnd.n4400 gnd.n4399 9.3005
R11376 gnd.n3721 gnd.n3720 9.3005
R11377 gnd.n4426 gnd.n4425 9.3005
R11378 gnd.n4427 gnd.n3719 9.3005
R11379 gnd.n4431 gnd.n4428 9.3005
R11380 gnd.n4430 gnd.n4429 9.3005
R11381 gnd.n3696 gnd.n3695 9.3005
R11382 gnd.n4456 gnd.n4455 9.3005
R11383 gnd.n4457 gnd.n3694 9.3005
R11384 gnd.n4471 gnd.n4458 9.3005
R11385 gnd.n4470 gnd.n4459 9.3005
R11386 gnd.n4469 gnd.n4460 9.3005
R11387 gnd.n4462 gnd.n4461 9.3005
R11388 gnd.n4464 gnd.n4463 9.3005
R11389 gnd.n3602 gnd.n3601 9.3005
R11390 gnd.n4531 gnd.n4530 9.3005
R11391 gnd.n4532 gnd.n3600 9.3005
R11392 gnd.n4536 gnd.n4533 9.3005
R11393 gnd.n4535 gnd.n4534 9.3005
R11394 gnd.n3576 gnd.n3575 9.3005
R11395 gnd.n4593 gnd.n4592 9.3005
R11396 gnd.n4594 gnd.n3574 9.3005
R11397 gnd.n4596 gnd.n4595 9.3005
R11398 gnd.n3558 gnd.n3557 9.3005
R11399 gnd.n4620 gnd.n4619 9.3005
R11400 gnd.n4621 gnd.n3556 9.3005
R11401 gnd.n4625 gnd.n4622 9.3005
R11402 gnd.n4624 gnd.n4623 9.3005
R11403 gnd.n3525 gnd.n3524 9.3005
R11404 gnd.n4671 gnd.n4670 9.3005
R11405 gnd.n4672 gnd.n3523 9.3005
R11406 gnd.n4674 gnd.n4673 9.3005
R11407 gnd.n3502 gnd.n3501 9.3005
R11408 gnd.n4711 gnd.n4710 9.3005
R11409 gnd.n4712 gnd.n3500 9.3005
R11410 gnd.n4714 gnd.n4713 9.3005
R11411 gnd.n3480 gnd.n3479 9.3005
R11412 gnd.n4767 gnd.n4766 9.3005
R11413 gnd.n4768 gnd.n3478 9.3005
R11414 gnd.n4770 gnd.n4769 9.3005
R11415 gnd.n3461 gnd.n3460 9.3005
R11416 gnd.n4792 gnd.n4791 9.3005
R11417 gnd.n4793 gnd.n3459 9.3005
R11418 gnd.n4795 gnd.n4794 9.3005
R11419 gnd.n3441 gnd.n3440 9.3005
R11420 gnd.n4852 gnd.n4851 9.3005
R11421 gnd.n4853 gnd.n3439 9.3005
R11422 gnd.n4855 gnd.n4854 9.3005
R11423 gnd.n3419 gnd.n3418 9.3005
R11424 gnd.n4881 gnd.n4880 9.3005
R11425 gnd.n4882 gnd.n3417 9.3005
R11426 gnd.n4886 gnd.n4883 9.3005
R11427 gnd.n4885 gnd.n4884 9.3005
R11428 gnd.n3391 gnd.n3390 9.3005
R11429 gnd.n4926 gnd.n4925 9.3005
R11430 gnd.n4927 gnd.n3389 9.3005
R11431 gnd.n4935 gnd.n4928 9.3005
R11432 gnd.n4934 gnd.n4929 9.3005
R11433 gnd.n4933 gnd.n4931 9.3005
R11434 gnd.n4930 gnd.n3315 9.3005
R11435 gnd.n5222 gnd.n3316 9.3005
R11436 gnd.n5221 gnd.n3317 9.3005
R11437 gnd.n5220 gnd.n3318 9.3005
R11438 gnd.n3325 gnd.n3319 9.3005
R11439 gnd.n5211 gnd.n3326 9.3005
R11440 gnd.n5210 gnd.n3327 9.3005
R11441 gnd.n5209 gnd.n3328 9.3005
R11442 gnd.n3337 gnd.n3329 9.3005
R11443 gnd.n5200 gnd.n3338 9.3005
R11444 gnd.n5199 gnd.n3339 9.3005
R11445 gnd.n5198 gnd.n3340 9.3005
R11446 gnd.n3349 gnd.n3341 9.3005
R11447 gnd.n5189 gnd.n3350 9.3005
R11448 gnd.n5188 gnd.n3351 9.3005
R11449 gnd.n5187 gnd.n3352 9.3005
R11450 gnd.n5175 gnd.n3353 9.3005
R11451 gnd.n5178 gnd.n5177 9.3005
R11452 gnd.n5176 gnd.n3005 9.3005
R11453 gnd.n5856 gnd.n3006 9.3005
R11454 gnd.n5855 gnd.n3007 9.3005
R11455 gnd.n5854 gnd.n3008 9.3005
R11456 gnd.n3014 gnd.n3009 9.3005
R11457 gnd.n5848 gnd.n3015 9.3005
R11458 gnd.n5847 gnd.n3016 9.3005
R11459 gnd.n5846 gnd.n3017 9.3005
R11460 gnd.n5608 gnd.n3018 9.3005
R11461 gnd.n5611 gnd.n5610 9.3005
R11462 gnd.n5612 gnd.n5607 9.3005
R11463 gnd.n5614 gnd.n5613 9.3005
R11464 gnd.n5605 gnd.n5604 9.3005
R11465 gnd.n5619 gnd.n5618 9.3005
R11466 gnd.n5620 gnd.n5603 9.3005
R11467 gnd.n5622 gnd.n5621 9.3005
R11468 gnd.n3216 gnd.n3215 9.3005
R11469 gnd.n5627 gnd.n5626 9.3005
R11470 gnd.n5628 gnd.n3214 9.3005
R11471 gnd.n5642 gnd.n5629 9.3005
R11472 gnd.n5641 gnd.n5630 9.3005
R11473 gnd.n5640 gnd.n5631 9.3005
R11474 gnd.n5633 gnd.n5632 9.3005
R11475 gnd.n5636 gnd.n5634 9.3005
R11476 gnd.n5764 gnd.n3147 9.3005
R11477 gnd.n3150 gnd.n3148 9.3005
R11478 gnd.n5760 gnd.n3151 9.3005
R11479 gnd.n5759 gnd.n3152 9.3005
R11480 gnd.n5758 gnd.n3153 9.3005
R11481 gnd.n3156 gnd.n3154 9.3005
R11482 gnd.n3188 gnd.n3157 9.3005
R11483 gnd.n3187 gnd.n3158 9.3005
R11484 gnd.n3186 gnd.n3159 9.3005
R11485 gnd.n3162 gnd.n3160 9.3005
R11486 gnd.n3182 gnd.n3163 9.3005
R11487 gnd.n3181 gnd.n3164 9.3005
R11488 gnd.n3180 gnd.n3165 9.3005
R11489 gnd.n3168 gnd.n3166 9.3005
R11490 gnd.n3176 gnd.n3169 9.3005
R11491 gnd.n3175 gnd.n3170 9.3005
R11492 gnd.n3174 gnd.n3172 9.3005
R11493 gnd.n3171 gnd.n246 9.3005
R11494 gnd.n7254 gnd.n247 9.3005
R11495 gnd.n7253 gnd.n248 9.3005
R11496 gnd.n7252 gnd.n249 9.3005
R11497 gnd.n254 gnd.n250 9.3005
R11498 gnd.n7246 gnd.n255 9.3005
R11499 gnd.n7245 gnd.n256 9.3005
R11500 gnd.n7244 gnd.n257 9.3005
R11501 gnd.n262 gnd.n258 9.3005
R11502 gnd.n7238 gnd.n263 9.3005
R11503 gnd.n7237 gnd.n264 9.3005
R11504 gnd.n7236 gnd.n265 9.3005
R11505 gnd.n7228 gnd.n266 9.3005
R11506 gnd.n4260 gnd.n4259 9.3005
R11507 gnd.n4164 gnd.n3836 9.3005
R11508 gnd.n4163 gnd.n3837 9.3005
R11509 gnd.n4162 gnd.n3838 9.3005
R11510 gnd.n4130 gnd.n3839 9.3005
R11511 gnd.n4152 gnd.n4131 9.3005
R11512 gnd.n4151 gnd.n4132 9.3005
R11513 gnd.n4150 gnd.n4133 9.3005
R11514 gnd.n4138 gnd.n4134 9.3005
R11515 gnd.n4140 gnd.n4139 9.3005
R11516 gnd.n3817 gnd.n3816 9.3005
R11517 gnd.n4200 gnd.n4199 9.3005
R11518 gnd.n4201 gnd.n3815 9.3005
R11519 gnd.n4203 gnd.n4202 9.3005
R11520 gnd.n3812 gnd.n3811 9.3005
R11521 gnd.n4214 gnd.n4213 9.3005
R11522 gnd.n4215 gnd.n3810 9.3005
R11523 gnd.n4218 gnd.n4217 9.3005
R11524 gnd.n4216 gnd.n3801 9.3005
R11525 gnd.n4262 gnd.n3802 9.3005
R11526 gnd.n4261 gnd.n3803 9.3005
R11527 gnd.n3868 gnd.n3835 9.3005
R11528 gnd.n3867 gnd.n3864 9.3005
R11529 gnd.n3879 gnd.n3863 9.3005
R11530 gnd.n3880 gnd.n3862 9.3005
R11531 gnd.n3881 gnd.n3861 9.3005
R11532 gnd.n3860 gnd.n3858 9.3005
R11533 gnd.n3887 gnd.n3857 9.3005
R11534 gnd.n3888 gnd.n3856 9.3005
R11535 gnd.n3889 gnd.n3855 9.3005
R11536 gnd.n3854 gnd.n3852 9.3005
R11537 gnd.n3895 gnd.n3851 9.3005
R11538 gnd.n3896 gnd.n3850 9.3005
R11539 gnd.n3897 gnd.n3849 9.3005
R11540 gnd.n3848 gnd.n3846 9.3005
R11541 gnd.n3902 gnd.n3845 9.3005
R11542 gnd.n3903 gnd.n3844 9.3005
R11543 gnd.n3842 gnd.n3841 9.3005
R11544 gnd.n3909 gnd.n3908 9.3005
R11545 gnd.n3873 gnd.n3870 9.3005
R11546 gnd.n3869 gnd.n3866 9.3005
R11547 gnd.n6035 gnd.n2750 9.3005
R11548 gnd.n6038 gnd.n2749 9.3005
R11549 gnd.n6039 gnd.n2748 9.3005
R11550 gnd.n6042 gnd.n2747 9.3005
R11551 gnd.n6043 gnd.n2746 9.3005
R11552 gnd.n6046 gnd.n2745 9.3005
R11553 gnd.n6047 gnd.n2744 9.3005
R11554 gnd.n6050 gnd.n2743 9.3005
R11555 gnd.n6052 gnd.n2740 9.3005
R11556 gnd.n6055 gnd.n2739 9.3005
R11557 gnd.n6056 gnd.n2738 9.3005
R11558 gnd.n6059 gnd.n2737 9.3005
R11559 gnd.n6060 gnd.n2736 9.3005
R11560 gnd.n6063 gnd.n2735 9.3005
R11561 gnd.n6064 gnd.n2734 9.3005
R11562 gnd.n6067 gnd.n2733 9.3005
R11563 gnd.n6068 gnd.n2732 9.3005
R11564 gnd.n6071 gnd.n2731 9.3005
R11565 gnd.n6072 gnd.n2730 9.3005
R11566 gnd.n6075 gnd.n2729 9.3005
R11567 gnd.n6076 gnd.n2728 9.3005
R11568 gnd.n6079 gnd.n2727 9.3005
R11569 gnd.n6080 gnd.n2726 9.3005
R11570 gnd.n6081 gnd.n2725 9.3005
R11571 gnd.n2724 gnd.n2721 9.3005
R11572 gnd.n2723 gnd.n2722 9.3005
R11573 gnd.n2847 gnd.n2846 9.3005
R11574 gnd.n2843 gnd.n2753 9.3005
R11575 gnd.n2840 gnd.n2754 9.3005
R11576 gnd.n2839 gnd.n2755 9.3005
R11577 gnd.n2836 gnd.n2756 9.3005
R11578 gnd.n2835 gnd.n2757 9.3005
R11579 gnd.n2832 gnd.n2758 9.3005
R11580 gnd.n2831 gnd.n2759 9.3005
R11581 gnd.n2828 gnd.n2827 9.3005
R11582 gnd.n2826 gnd.n2760 9.3005
R11583 gnd.n2825 gnd.n2824 9.3005
R11584 gnd.n2821 gnd.n2763 9.3005
R11585 gnd.n2818 gnd.n2764 9.3005
R11586 gnd.n2817 gnd.n2765 9.3005
R11587 gnd.n2814 gnd.n2766 9.3005
R11588 gnd.n2813 gnd.n2767 9.3005
R11589 gnd.n2810 gnd.n2768 9.3005
R11590 gnd.n2809 gnd.n2769 9.3005
R11591 gnd.n2806 gnd.n2770 9.3005
R11592 gnd.n2805 gnd.n2771 9.3005
R11593 gnd.n2802 gnd.n2772 9.3005
R11594 gnd.n2801 gnd.n2773 9.3005
R11595 gnd.n2798 gnd.n2774 9.3005
R11596 gnd.n2797 gnd.n2775 9.3005
R11597 gnd.n2794 gnd.n2776 9.3005
R11598 gnd.n2793 gnd.n2777 9.3005
R11599 gnd.n2790 gnd.n2778 9.3005
R11600 gnd.n2789 gnd.n2779 9.3005
R11601 gnd.n2786 gnd.n2785 9.3005
R11602 gnd.n2784 gnd.n2781 9.3005
R11603 gnd.n2848 gnd.n2751 9.3005
R11604 gnd.n4125 gnd.n2380 9.3005
R11605 gnd.n6288 gnd.n2381 9.3005
R11606 gnd.n6287 gnd.n2382 9.3005
R11607 gnd.n6286 gnd.n2383 9.3005
R11608 gnd.n4128 gnd.n2384 9.3005
R11609 gnd.n6276 gnd.n2402 9.3005
R11610 gnd.n6275 gnd.n2403 9.3005
R11611 gnd.n6274 gnd.n2404 9.3005
R11612 gnd.n4135 gnd.n2405 9.3005
R11613 gnd.n6264 gnd.n2423 9.3005
R11614 gnd.n6263 gnd.n2424 9.3005
R11615 gnd.n6262 gnd.n2425 9.3005
R11616 gnd.n3814 gnd.n2426 9.3005
R11617 gnd.n6252 gnd.n2443 9.3005
R11618 gnd.n6251 gnd.n2444 9.3005
R11619 gnd.n6250 gnd.n2445 9.3005
R11620 gnd.n3809 gnd.n2446 9.3005
R11621 gnd.n6239 gnd.n2462 9.3005
R11622 gnd.n6238 gnd.n2463 9.3005
R11623 gnd.n6237 gnd.n2464 9.3005
R11624 gnd.n4226 gnd.n2465 9.3005
R11625 gnd.n6226 gnd.n2478 9.3005
R11626 gnd.n6225 gnd.n2479 9.3005
R11627 gnd.n6224 gnd.n2480 9.3005
R11628 gnd.n4246 gnd.n2481 9.3005
R11629 gnd.n6213 gnd.n2496 9.3005
R11630 gnd.n6212 gnd.n2497 9.3005
R11631 gnd.n6211 gnd.n2498 9.3005
R11632 gnd.n3780 gnd.n2499 9.3005
R11633 gnd.n6201 gnd.n2515 9.3005
R11634 gnd.n6200 gnd.n2516 9.3005
R11635 gnd.n6199 gnd.n2517 9.3005
R11636 gnd.n4297 gnd.n2518 9.3005
R11637 gnd.n6189 gnd.n2536 9.3005
R11638 gnd.n6188 gnd.n2537 9.3005
R11639 gnd.n6187 gnd.n2538 9.3005
R11640 gnd.n4307 gnd.n2539 9.3005
R11641 gnd.n6177 gnd.n2556 9.3005
R11642 gnd.n6176 gnd.n2557 9.3005
R11643 gnd.n6175 gnd.n2558 9.3005
R11644 gnd.n2576 gnd.n2559 9.3005
R11645 gnd.n6165 gnd.n6164 9.3005
R11646 gnd.n4124 gnd.n4123 9.3005
R11647 gnd.n4126 gnd.n4125 9.3005
R11648 gnd.n4127 gnd.n2381 9.3005
R11649 gnd.n4158 gnd.n2382 9.3005
R11650 gnd.n4157 gnd.n2383 9.3005
R11651 gnd.n4156 gnd.n4128 9.3005
R11652 gnd.n4129 gnd.n2402 9.3005
R11653 gnd.n4146 gnd.n2403 9.3005
R11654 gnd.n4145 gnd.n2404 9.3005
R11655 gnd.n4144 gnd.n4135 9.3005
R11656 gnd.n4137 gnd.n2423 9.3005
R11657 gnd.n4136 gnd.n2424 9.3005
R11658 gnd.n3813 gnd.n2425 9.3005
R11659 gnd.n4207 gnd.n3814 9.3005
R11660 gnd.n4208 gnd.n2443 9.3005
R11661 gnd.n4209 gnd.n2444 9.3005
R11662 gnd.n3808 gnd.n2445 9.3005
R11663 gnd.n4222 gnd.n3809 9.3005
R11664 gnd.n4223 gnd.n2462 9.3005
R11665 gnd.n4224 gnd.n2463 9.3005
R11666 gnd.n4225 gnd.n2464 9.3005
R11667 gnd.n4229 gnd.n4226 9.3005
R11668 gnd.n4230 gnd.n2478 9.3005
R11669 gnd.n4244 gnd.n2479 9.3005
R11670 gnd.n4245 gnd.n2480 9.3005
R11671 gnd.n4249 gnd.n4246 9.3005
R11672 gnd.n4248 gnd.n2496 9.3005
R11673 gnd.n4247 gnd.n2497 9.3005
R11674 gnd.n3779 gnd.n2498 9.3005
R11675 gnd.n4293 gnd.n3780 9.3005
R11676 gnd.n4294 gnd.n2515 9.3005
R11677 gnd.n4295 gnd.n2516 9.3005
R11678 gnd.n4296 gnd.n2517 9.3005
R11679 gnd.n4300 gnd.n4297 9.3005
R11680 gnd.n4301 gnd.n2536 9.3005
R11681 gnd.n4305 gnd.n2537 9.3005
R11682 gnd.n4306 gnd.n2538 9.3005
R11683 gnd.n4310 gnd.n4307 9.3005
R11684 gnd.n4311 gnd.n2556 9.3005
R11685 gnd.n4312 gnd.n2557 9.3005
R11686 gnd.n2578 gnd.n2558 9.3005
R11687 gnd.n6162 gnd.n2576 9.3005
R11688 gnd.n6164 gnd.n6163 9.3005
R11689 gnd.n4124 gnd.n3840 9.3005
R11690 gnd.n3913 gnd.n3910 9.3005
R11691 gnd.n4111 gnd.n3914 9.3005
R11692 gnd.n4113 gnd.n4112 9.3005
R11693 gnd.n4110 gnd.n3916 9.3005
R11694 gnd.n4109 gnd.n4108 9.3005
R11695 gnd.n3918 gnd.n3917 9.3005
R11696 gnd.n4102 gnd.n4101 9.3005
R11697 gnd.n4100 gnd.n3920 9.3005
R11698 gnd.n4099 gnd.n4098 9.3005
R11699 gnd.n3922 gnd.n3921 9.3005
R11700 gnd.n4092 gnd.n4091 9.3005
R11701 gnd.n4090 gnd.n3924 9.3005
R11702 gnd.n4089 gnd.n4088 9.3005
R11703 gnd.n3926 gnd.n3925 9.3005
R11704 gnd.n4082 gnd.n4081 9.3005
R11705 gnd.n4080 gnd.n3928 9.3005
R11706 gnd.n4079 gnd.n4078 9.3005
R11707 gnd.n3930 gnd.n3929 9.3005
R11708 gnd.n4072 gnd.n4071 9.3005
R11709 gnd.n4070 gnd.n3932 9.3005
R11710 gnd.n3934 gnd.n3933 9.3005
R11711 gnd.n4060 gnd.n4059 9.3005
R11712 gnd.n4058 gnd.n3936 9.3005
R11713 gnd.n4057 gnd.n4056 9.3005
R11714 gnd.n3938 gnd.n3937 9.3005
R11715 gnd.n4050 gnd.n4049 9.3005
R11716 gnd.n4048 gnd.n3940 9.3005
R11717 gnd.n4047 gnd.n4046 9.3005
R11718 gnd.n3942 gnd.n3941 9.3005
R11719 gnd.n4040 gnd.n4039 9.3005
R11720 gnd.n4038 gnd.n3944 9.3005
R11721 gnd.n4037 gnd.n4036 9.3005
R11722 gnd.n3946 gnd.n3945 9.3005
R11723 gnd.n4030 gnd.n4029 9.3005
R11724 gnd.n4028 gnd.n3948 9.3005
R11725 gnd.n4027 gnd.n4026 9.3005
R11726 gnd.n3950 gnd.n3949 9.3005
R11727 gnd.n4020 gnd.n4019 9.3005
R11728 gnd.n4018 gnd.n3952 9.3005
R11729 gnd.n4017 gnd.n4016 9.3005
R11730 gnd.n3954 gnd.n3953 9.3005
R11731 gnd.n4010 gnd.n4009 9.3005
R11732 gnd.n4008 gnd.n3959 9.3005
R11733 gnd.n4007 gnd.n4006 9.3005
R11734 gnd.n3961 gnd.n3960 9.3005
R11735 gnd.n4000 gnd.n3999 9.3005
R11736 gnd.n3998 gnd.n3963 9.3005
R11737 gnd.n3997 gnd.n3996 9.3005
R11738 gnd.n3965 gnd.n3964 9.3005
R11739 gnd.n3990 gnd.n3989 9.3005
R11740 gnd.n3988 gnd.n3967 9.3005
R11741 gnd.n3987 gnd.n3986 9.3005
R11742 gnd.n3969 gnd.n3968 9.3005
R11743 gnd.n3980 gnd.n3979 9.3005
R11744 gnd.n3978 gnd.n3971 9.3005
R11745 gnd.n3977 gnd.n3976 9.3005
R11746 gnd.n3973 gnd.n3972 9.3005
R11747 gnd.n4069 gnd.n4068 9.3005
R11748 gnd.n4121 gnd.n4120 9.3005
R11749 gnd.n6293 gnd.n2371 9.3005
R11750 gnd.n6292 gnd.n2372 9.3005
R11751 gnd.n2391 gnd.n2373 9.3005
R11752 gnd.n6282 gnd.n2392 9.3005
R11753 gnd.n6281 gnd.n2393 9.3005
R11754 gnd.n6280 gnd.n2394 9.3005
R11755 gnd.n2412 gnd.n2395 9.3005
R11756 gnd.n6270 gnd.n2413 9.3005
R11757 gnd.n6269 gnd.n2414 9.3005
R11758 gnd.n6268 gnd.n2415 9.3005
R11759 gnd.n2432 gnd.n2416 9.3005
R11760 gnd.n6258 gnd.n2433 9.3005
R11761 gnd.n6257 gnd.n2434 9.3005
R11762 gnd.n6256 gnd.n2435 9.3005
R11763 gnd.n2453 gnd.n2436 9.3005
R11764 gnd.n2505 gnd.n2489 9.3005
R11765 gnd.n6207 gnd.n2506 9.3005
R11766 gnd.n6206 gnd.n2507 9.3005
R11767 gnd.n6205 gnd.n2508 9.3005
R11768 gnd.n2525 gnd.n2509 9.3005
R11769 gnd.n6195 gnd.n2526 9.3005
R11770 gnd.n6194 gnd.n2527 9.3005
R11771 gnd.n6193 gnd.n2528 9.3005
R11772 gnd.n2545 gnd.n2529 9.3005
R11773 gnd.n6183 gnd.n2546 9.3005
R11774 gnd.n6182 gnd.n2547 9.3005
R11775 gnd.n6181 gnd.n2548 9.3005
R11776 gnd.n2566 gnd.n2549 9.3005
R11777 gnd.n6171 gnd.n2567 9.3005
R11778 gnd.n6170 gnd.n2568 9.3005
R11779 gnd.n6169 gnd.n2569 9.3005
R11780 gnd.n6294 gnd.n2370 9.3005
R11781 gnd.n6217 gnd.n2454 9.3005
R11782 gnd.n875 gnd.n874 9.3005
R11783 gnd.n6318 gnd.n2342 9.3005
R11784 gnd.n6317 gnd.n2343 9.3005
R11785 gnd.n6316 gnd.n2344 9.3005
R11786 gnd.n2349 gnd.n2345 9.3005
R11787 gnd.n6310 gnd.n2350 9.3005
R11788 gnd.n6309 gnd.n2351 9.3005
R11789 gnd.n6308 gnd.n2352 9.3005
R11790 gnd.n2357 gnd.n2353 9.3005
R11791 gnd.n6302 gnd.n2358 9.3005
R11792 gnd.n6301 gnd.n2359 9.3005
R11793 gnd.n6300 gnd.n2360 9.3005
R11794 gnd.n3830 gnd.n2361 9.3005
R11795 gnd.n3832 gnd.n3831 9.3005
R11796 gnd.n4170 gnd.n4169 9.3005
R11797 gnd.n4171 gnd.n3829 9.3005
R11798 gnd.n4173 gnd.n4172 9.3005
R11799 gnd.n3827 gnd.n3826 9.3005
R11800 gnd.n4178 gnd.n4177 9.3005
R11801 gnd.n4179 gnd.n3825 9.3005
R11802 gnd.n4181 gnd.n4180 9.3005
R11803 gnd.n3823 gnd.n3822 9.3005
R11804 gnd.n4186 gnd.n4185 9.3005
R11805 gnd.n4187 gnd.n3821 9.3005
R11806 gnd.n4194 gnd.n4188 9.3005
R11807 gnd.n4193 gnd.n4189 9.3005
R11808 gnd.n4192 gnd.n4190 9.3005
R11809 gnd.n3794 gnd.n3793 9.3005
R11810 gnd.n4274 gnd.n4273 9.3005
R11811 gnd.n6325 gnd.n6324 9.3005
R11812 gnd.n6328 gnd.n873 9.3005
R11813 gnd.n872 gnd.n868 9.3005
R11814 gnd.n6334 gnd.n867 9.3005
R11815 gnd.n6335 gnd.n866 9.3005
R11816 gnd.n6336 gnd.n865 9.3005
R11817 gnd.n864 gnd.n860 9.3005
R11818 gnd.n6342 gnd.n859 9.3005
R11819 gnd.n6343 gnd.n858 9.3005
R11820 gnd.n6344 gnd.n857 9.3005
R11821 gnd.n856 gnd.n852 9.3005
R11822 gnd.n6350 gnd.n851 9.3005
R11823 gnd.n6351 gnd.n850 9.3005
R11824 gnd.n6352 gnd.n849 9.3005
R11825 gnd.n848 gnd.n844 9.3005
R11826 gnd.n6358 gnd.n843 9.3005
R11827 gnd.n6359 gnd.n842 9.3005
R11828 gnd.n6360 gnd.n841 9.3005
R11829 gnd.n840 gnd.n836 9.3005
R11830 gnd.n6366 gnd.n835 9.3005
R11831 gnd.n6367 gnd.n834 9.3005
R11832 gnd.n6368 gnd.n833 9.3005
R11833 gnd.n832 gnd.n828 9.3005
R11834 gnd.n6374 gnd.n827 9.3005
R11835 gnd.n6375 gnd.n826 9.3005
R11836 gnd.n6376 gnd.n825 9.3005
R11837 gnd.n824 gnd.n820 9.3005
R11838 gnd.n6382 gnd.n819 9.3005
R11839 gnd.n6383 gnd.n818 9.3005
R11840 gnd.n6384 gnd.n817 9.3005
R11841 gnd.n816 gnd.n812 9.3005
R11842 gnd.n6390 gnd.n811 9.3005
R11843 gnd.n6391 gnd.n810 9.3005
R11844 gnd.n6392 gnd.n809 9.3005
R11845 gnd.n808 gnd.n804 9.3005
R11846 gnd.n6398 gnd.n803 9.3005
R11847 gnd.n6399 gnd.n802 9.3005
R11848 gnd.n6400 gnd.n801 9.3005
R11849 gnd.n800 gnd.n796 9.3005
R11850 gnd.n6406 gnd.n795 9.3005
R11851 gnd.n6407 gnd.n794 9.3005
R11852 gnd.n6408 gnd.n793 9.3005
R11853 gnd.n792 gnd.n788 9.3005
R11854 gnd.n6414 gnd.n787 9.3005
R11855 gnd.n6415 gnd.n786 9.3005
R11856 gnd.n6416 gnd.n785 9.3005
R11857 gnd.n784 gnd.n780 9.3005
R11858 gnd.n6422 gnd.n779 9.3005
R11859 gnd.n6423 gnd.n778 9.3005
R11860 gnd.n6424 gnd.n777 9.3005
R11861 gnd.n776 gnd.n772 9.3005
R11862 gnd.n6430 gnd.n771 9.3005
R11863 gnd.n6431 gnd.n770 9.3005
R11864 gnd.n6432 gnd.n769 9.3005
R11865 gnd.n768 gnd.n764 9.3005
R11866 gnd.n6438 gnd.n763 9.3005
R11867 gnd.n6439 gnd.n762 9.3005
R11868 gnd.n6440 gnd.n761 9.3005
R11869 gnd.n760 gnd.n756 9.3005
R11870 gnd.n6446 gnd.n755 9.3005
R11871 gnd.n6447 gnd.n754 9.3005
R11872 gnd.n6448 gnd.n753 9.3005
R11873 gnd.n752 gnd.n748 9.3005
R11874 gnd.n6454 gnd.n747 9.3005
R11875 gnd.n6455 gnd.n746 9.3005
R11876 gnd.n6456 gnd.n745 9.3005
R11877 gnd.n744 gnd.n740 9.3005
R11878 gnd.n6462 gnd.n739 9.3005
R11879 gnd.n6463 gnd.n738 9.3005
R11880 gnd.n6464 gnd.n737 9.3005
R11881 gnd.n736 gnd.n732 9.3005
R11882 gnd.n6470 gnd.n731 9.3005
R11883 gnd.n6471 gnd.n730 9.3005
R11884 gnd.n6472 gnd.n729 9.3005
R11885 gnd.n728 gnd.n724 9.3005
R11886 gnd.n6478 gnd.n723 9.3005
R11887 gnd.n6479 gnd.n722 9.3005
R11888 gnd.n6480 gnd.n721 9.3005
R11889 gnd.n720 gnd.n716 9.3005
R11890 gnd.n6486 gnd.n715 9.3005
R11891 gnd.n6487 gnd.n714 9.3005
R11892 gnd.n6488 gnd.n713 9.3005
R11893 gnd.n712 gnd.n708 9.3005
R11894 gnd.n6494 gnd.n707 9.3005
R11895 gnd.n6496 gnd.n6495 9.3005
R11896 gnd.n6327 gnd.n6326 9.3005
R11897 gnd.n5169 gnd.n5168 9.3005
R11898 gnd.n4387 gnd.n4383 9.3005
R11899 gnd.n4390 gnd.n4389 9.3005
R11900 gnd.n4388 gnd.n4384 9.3005
R11901 gnd.n3727 gnd.n3726 9.3005
R11902 gnd.n4416 gnd.n4415 9.3005
R11903 gnd.n4417 gnd.n3724 9.3005
R11904 gnd.n4420 gnd.n4419 9.3005
R11905 gnd.n4418 gnd.n3725 9.3005
R11906 gnd.n3703 gnd.n3702 9.3005
R11907 gnd.n4446 gnd.n4445 9.3005
R11908 gnd.n4447 gnd.n3700 9.3005
R11909 gnd.n4450 gnd.n4449 9.3005
R11910 gnd.n4448 gnd.n3701 9.3005
R11911 gnd.n3678 gnd.n3677 9.3005
R11912 gnd.n4486 gnd.n4485 9.3005
R11913 gnd.n4487 gnd.n3675 9.3005
R11914 gnd.n4493 gnd.n4492 9.3005
R11915 gnd.n4491 gnd.n3676 9.3005
R11916 gnd.n4490 gnd.n4489 9.3005
R11917 gnd.n3594 gnd.n3593 9.3005
R11918 gnd.n4542 gnd.n4541 9.3005
R11919 gnd.n4543 gnd.n3591 9.3005
R11920 gnd.n4565 gnd.n4564 9.3005
R11921 gnd.n4563 gnd.n3592 9.3005
R11922 gnd.n4562 gnd.n4561 9.3005
R11923 gnd.n4560 gnd.n4544 9.3005
R11924 gnd.n4559 gnd.n4558 9.3005
R11925 gnd.n4557 gnd.n4551 9.3005
R11926 gnd.n4556 gnd.n4555 9.3005
R11927 gnd.n4554 gnd.n4553 9.3005
R11928 gnd.n4552 gnd.n3544 9.3005
R11929 gnd.n3542 gnd.n3541 9.3005
R11930 gnd.n4644 gnd.n4643 9.3005
R11931 gnd.n4645 gnd.n3540 9.3005
R11932 gnd.n4647 gnd.n4646 9.3005
R11933 gnd.n3517 gnd.n3515 9.3005
R11934 gnd.n4695 gnd.n4694 9.3005
R11935 gnd.n4693 gnd.n3516 9.3005
R11936 gnd.n4692 gnd.n4691 9.3005
R11937 gnd.n3494 gnd.n3492 9.3005
R11938 gnd.n4753 gnd.n4752 9.3005
R11939 gnd.n4751 gnd.n3493 9.3005
R11940 gnd.n4750 gnd.n4749 9.3005
R11941 gnd.n4748 gnd.n3495 9.3005
R11942 gnd.n4747 gnd.n4746 9.3005
R11943 gnd.n4745 gnd.n4734 9.3005
R11944 gnd.n4744 gnd.n4743 9.3005
R11945 gnd.n4742 gnd.n4735 9.3005
R11946 gnd.n4741 gnd.n4740 9.3005
R11947 gnd.n3434 gnd.n3433 9.3005
R11948 gnd.n4862 gnd.n4861 9.3005
R11949 gnd.n4863 gnd.n3431 9.3005
R11950 gnd.n4866 gnd.n4865 9.3005
R11951 gnd.n4864 gnd.n3432 9.3005
R11952 gnd.n3405 gnd.n3404 9.3005
R11953 gnd.n4901 gnd.n4900 9.3005
R11954 gnd.n4902 gnd.n3402 9.3005
R11955 gnd.n4911 gnd.n4910 9.3005
R11956 gnd.n4909 gnd.n3403 9.3005
R11957 gnd.n4908 gnd.n4907 9.3005
R11958 gnd.n4906 gnd.n4903 9.3005
R11959 gnd.n3370 gnd.n3369 9.3005
R11960 gnd.n4958 gnd.n4957 9.3005
R11961 gnd.n4959 gnd.n3368 9.3005
R11962 gnd.n4961 gnd.n4960 9.3005
R11963 gnd.n4964 gnd.n3367 9.3005
R11964 gnd.n4966 gnd.n4965 9.3005
R11965 gnd.n4967 gnd.n3366 9.3005
R11966 gnd.n4969 gnd.n4968 9.3005
R11967 gnd.n4972 gnd.n3365 9.3005
R11968 gnd.n4974 gnd.n4973 9.3005
R11969 gnd.n4975 gnd.n3364 9.3005
R11970 gnd.n4977 gnd.n4976 9.3005
R11971 gnd.n4980 gnd.n3363 9.3005
R11972 gnd.n4982 gnd.n4981 9.3005
R11973 gnd.n4983 gnd.n3362 9.3005
R11974 gnd.n4985 gnd.n4984 9.3005
R11975 gnd.n4988 gnd.n3361 9.3005
R11976 gnd.n4990 gnd.n4989 9.3005
R11977 gnd.n4991 gnd.n3359 9.3005
R11978 gnd.n5172 gnd.n5171 9.3005
R11979 gnd.n5170 gnd.n3360 9.3005
R11980 gnd.n4386 gnd.n4385 9.3005
R11981 gnd.n6152 gnd.n2582 9.3005
R11982 gnd.n4258 gnd.n3805 9.3005
R11983 gnd.n4257 gnd.n4256 9.3005
R11984 gnd.n4255 gnd.n3806 9.3005
R11985 gnd.n4254 gnd.n4253 9.3005
R11986 gnd.n3783 gnd.n3782 9.3005
R11987 gnd.n4286 gnd.n4285 9.3005
R11988 gnd.n4287 gnd.n3781 9.3005
R11989 gnd.n4289 gnd.n4288 9.3005
R11990 gnd.n3772 gnd.n3770 9.3005
R11991 gnd.n4329 gnd.n4328 9.3005
R11992 gnd.n4327 gnd.n3771 9.3005
R11993 gnd.n4326 gnd.n4325 9.3005
R11994 gnd.n4324 gnd.n3773 9.3005
R11995 gnd.n4323 gnd.n4322 9.3005
R11996 gnd.n4321 gnd.n3776 9.3005
R11997 gnd.n4320 gnd.n4319 9.3005
R11998 gnd.n4318 gnd.n3777 9.3005
R11999 gnd.n4317 gnd.n4316 9.3005
R12000 gnd.n2581 gnd.n2579 9.3005
R12001 gnd.n6158 gnd.n6157 9.3005
R12002 gnd.n6156 gnd.n2580 9.3005
R12003 gnd.n6130 gnd.n6129 9.3005
R12004 gnd.n6128 gnd.n6127 9.3005
R12005 gnd.n2624 gnd.n2623 9.3005
R12006 gnd.n6122 gnd.n6121 9.3005
R12007 gnd.n6120 gnd.n6119 9.3005
R12008 gnd.n2634 gnd.n2633 9.3005
R12009 gnd.n6114 gnd.n6113 9.3005
R12010 gnd.n6112 gnd.n6111 9.3005
R12011 gnd.n2642 gnd.n2641 9.3005
R12012 gnd.n6106 gnd.n6105 9.3005
R12013 gnd.n6104 gnd.n6103 9.3005
R12014 gnd.n2652 gnd.n2651 9.3005
R12015 gnd.n6098 gnd.n6097 9.3005
R12016 gnd.n6096 gnd.n6095 9.3005
R12017 gnd.n2660 gnd.n2659 9.3005
R12018 gnd.n6090 gnd.n6089 9.3005
R12019 gnd.n6088 gnd.n2674 9.3005
R12020 gnd.n6087 gnd.n2583 9.3005
R12021 gnd.n2620 gnd.n2618 9.3005
R12022 gnd.n6154 gnd.n6153 9.3005
R12023 gnd.n2673 gnd.n2584 9.3005
R12024 gnd.n2669 gnd.n2668 9.3005
R12025 gnd.n6092 gnd.n6091 9.3005
R12026 gnd.n6094 gnd.n6093 9.3005
R12027 gnd.n2656 gnd.n2655 9.3005
R12028 gnd.n6100 gnd.n6099 9.3005
R12029 gnd.n6102 gnd.n6101 9.3005
R12030 gnd.n2648 gnd.n2647 9.3005
R12031 gnd.n6108 gnd.n6107 9.3005
R12032 gnd.n6110 gnd.n6109 9.3005
R12033 gnd.n2638 gnd.n2637 9.3005
R12034 gnd.n6116 gnd.n6115 9.3005
R12035 gnd.n6118 gnd.n6117 9.3005
R12036 gnd.n2630 gnd.n2629 9.3005
R12037 gnd.n6124 gnd.n6123 9.3005
R12038 gnd.n6126 gnd.n6125 9.3005
R12039 gnd.n2619 gnd.n2617 9.3005
R12040 gnd.n6132 gnd.n6131 9.3005
R12041 gnd.n6133 gnd.n2612 9.3005
R12042 gnd.n6135 gnd.n6134 9.3005
R12043 gnd.n6137 gnd.n2611 9.3005
R12044 gnd.n6139 gnd.n6138 9.3005
R12045 gnd.n6140 gnd.n2607 9.3005
R12046 gnd.n6142 gnd.n6141 9.3005
R12047 gnd.n6143 gnd.n2606 9.3005
R12048 gnd.n6145 gnd.n6144 9.3005
R12049 gnd.n6146 gnd.n2605 9.3005
R12050 gnd.n4379 gnd.n4378 9.3005
R12051 gnd.n3737 gnd.n3736 9.3005
R12052 gnd.n4407 gnd.n4406 9.3005
R12053 gnd.n4408 gnd.n3734 9.3005
R12054 gnd.n4411 gnd.n4410 9.3005
R12055 gnd.n4409 gnd.n3735 9.3005
R12056 gnd.n3712 gnd.n3711 9.3005
R12057 gnd.n4437 gnd.n4436 9.3005
R12058 gnd.n4438 gnd.n3709 9.3005
R12059 gnd.n4441 gnd.n4440 9.3005
R12060 gnd.n4439 gnd.n3710 9.3005
R12061 gnd.n3687 gnd.n3686 9.3005
R12062 gnd.n4477 gnd.n4476 9.3005
R12063 gnd.n4478 gnd.n3684 9.3005
R12064 gnd.n4481 gnd.n4480 9.3005
R12065 gnd.n4479 gnd.n3685 9.3005
R12066 gnd.n2919 gnd.n2917 9.3005
R12067 gnd.n5957 gnd.n5956 9.3005
R12068 gnd.n5955 gnd.n2918 9.3005
R12069 gnd.n5954 gnd.n5953 9.3005
R12070 gnd.n5952 gnd.n2920 9.3005
R12071 gnd.n5951 gnd.n5950 9.3005
R12072 gnd.n5949 gnd.n2924 9.3005
R12073 gnd.n5948 gnd.n5947 9.3005
R12074 gnd.n5946 gnd.n2925 9.3005
R12075 gnd.n5945 gnd.n5944 9.3005
R12076 gnd.n5943 gnd.n2929 9.3005
R12077 gnd.n5942 gnd.n5941 9.3005
R12078 gnd.n5940 gnd.n2930 9.3005
R12079 gnd.n5939 gnd.n5938 9.3005
R12080 gnd.n5937 gnd.n2934 9.3005
R12081 gnd.n5936 gnd.n5935 9.3005
R12082 gnd.n5934 gnd.n2935 9.3005
R12083 gnd.n5933 gnd.n5932 9.3005
R12084 gnd.n5931 gnd.n2939 9.3005
R12085 gnd.n5930 gnd.n5929 9.3005
R12086 gnd.n5928 gnd.n2940 9.3005
R12087 gnd.n5927 gnd.n5926 9.3005
R12088 gnd.n5925 gnd.n2944 9.3005
R12089 gnd.n5924 gnd.n5923 9.3005
R12090 gnd.n5922 gnd.n2945 9.3005
R12091 gnd.n5921 gnd.n5920 9.3005
R12092 gnd.n5919 gnd.n2949 9.3005
R12093 gnd.n5918 gnd.n5917 9.3005
R12094 gnd.n5916 gnd.n2950 9.3005
R12095 gnd.n5915 gnd.n5914 9.3005
R12096 gnd.n5913 gnd.n2954 9.3005
R12097 gnd.n5912 gnd.n5911 9.3005
R12098 gnd.n5910 gnd.n2955 9.3005
R12099 gnd.n5909 gnd.n5908 9.3005
R12100 gnd.n5907 gnd.n2959 9.3005
R12101 gnd.n5906 gnd.n5905 9.3005
R12102 gnd.n5904 gnd.n2960 9.3005
R12103 gnd.n5903 gnd.n5902 9.3005
R12104 gnd.n5901 gnd.n2964 9.3005
R12105 gnd.n5900 gnd.n5899 9.3005
R12106 gnd.n5898 gnd.n2965 9.3005
R12107 gnd.n5897 gnd.n5896 9.3005
R12108 gnd.n5895 gnd.n2969 9.3005
R12109 gnd.n5894 gnd.n5893 9.3005
R12110 gnd.n5892 gnd.n2970 9.3005
R12111 gnd.n5891 gnd.n5890 9.3005
R12112 gnd.n5889 gnd.n2974 9.3005
R12113 gnd.n5888 gnd.n5887 9.3005
R12114 gnd.n5886 gnd.n2975 9.3005
R12115 gnd.n5885 gnd.n5884 9.3005
R12116 gnd.n5883 gnd.n2979 9.3005
R12117 gnd.n5882 gnd.n5881 9.3005
R12118 gnd.n5880 gnd.n2980 9.3005
R12119 gnd.n5879 gnd.n5878 9.3005
R12120 gnd.n5877 gnd.n2984 9.3005
R12121 gnd.n5876 gnd.n5875 9.3005
R12122 gnd.n5874 gnd.n2985 9.3005
R12123 gnd.n5873 gnd.n5872 9.3005
R12124 gnd.n5871 gnd.n2989 9.3005
R12125 gnd.n5870 gnd.n5869 9.3005
R12126 gnd.n5868 gnd.n2990 9.3005
R12127 gnd.n5867 gnd.n5866 9.3005
R12128 gnd.n5865 gnd.n2994 9.3005
R12129 gnd.n5864 gnd.n5863 9.3005
R12130 gnd.n5862 gnd.n2995 9.3005
R12131 gnd.n5861 gnd.n2998 9.3005
R12132 gnd.n4377 gnd.n4376 9.3005
R12133 gnd.n5058 gnd.n5057 9.3005
R12134 gnd.n5053 gnd.n5052 9.3005
R12135 gnd.n5065 gnd.n5064 9.3005
R12136 gnd.n5066 gnd.n5051 9.3005
R12137 gnd.n5069 gnd.n5068 9.3005
R12138 gnd.n5067 gnd.n5049 9.3005
R12139 gnd.n5056 gnd.n5055 9.3005
R12140 gnd.n5157 gnd.n5005 9.3005
R12141 gnd.n5018 gnd.n5014 9.3005
R12142 gnd.n5151 gnd.n5150 9.3005
R12143 gnd.n5139 gnd.n5016 9.3005
R12144 gnd.n5138 gnd.n5137 9.3005
R12145 gnd.n5027 gnd.n5023 9.3005
R12146 gnd.n5131 gnd.n5130 9.3005
R12147 gnd.n5120 gnd.n5025 9.3005
R12148 gnd.n5119 gnd.n5118 9.3005
R12149 gnd.n5036 gnd.n5032 9.3005
R12150 gnd.n5112 gnd.n5111 9.3005
R12151 gnd.n5101 gnd.n5034 9.3005
R12152 gnd.n5100 gnd.n5099 9.3005
R12153 gnd.n5045 gnd.n5041 9.3005
R12154 gnd.n5093 gnd.n5092 9.3005
R12155 gnd.n5082 gnd.n5043 9.3005
R12156 gnd.n5081 gnd.n5080 9.3005
R12157 gnd.n5159 gnd.n5158 9.3005
R12158 gnd.n5009 gnd.n5008 9.3005
R12159 gnd.n5076 gnd.n5075 9.3005
R12160 gnd.n5077 gnd.n5048 9.3005
R12161 gnd.n5084 gnd.n5083 9.3005
R12162 gnd.n5046 gnd.n5044 9.3005
R12163 gnd.n5091 gnd.n5090 9.3005
R12164 gnd.n5040 gnd.n5039 9.3005
R12165 gnd.n5103 gnd.n5102 9.3005
R12166 gnd.n5037 gnd.n5035 9.3005
R12167 gnd.n5110 gnd.n5109 9.3005
R12168 gnd.n5031 gnd.n5030 9.3005
R12169 gnd.n5122 gnd.n5121 9.3005
R12170 gnd.n5028 gnd.n5026 9.3005
R12171 gnd.n5129 gnd.n5128 9.3005
R12172 gnd.n5022 gnd.n5021 9.3005
R12173 gnd.n5141 gnd.n5140 9.3005
R12174 gnd.n5019 gnd.n5017 9.3005
R12175 gnd.n5149 gnd.n5148 9.3005
R12176 gnd.n5147 gnd.n5146 9.3005
R12177 gnd.n5161 gnd.n5160 9.3005
R12178 gnd.n5006 gnd.n5000 9.3005
R12179 gnd.n5007 gnd.n4999 9.3005
R12180 gnd.n4995 gnd.n4992 9.3005
R12181 gnd.n3226 gnd.n3225 9.3005
R12182 gnd.n5575 gnd.n5574 9.3005
R12183 gnd.n5576 gnd.n3224 9.3005
R12184 gnd.n5578 gnd.n5577 9.3005
R12185 gnd.n3220 gnd.n3218 9.3005
R12186 gnd.n5598 gnd.n5597 9.3005
R12187 gnd.n5596 gnd.n3219 9.3005
R12188 gnd.n5595 gnd.n5594 9.3005
R12189 gnd.n5593 gnd.n3221 9.3005
R12190 gnd.n5592 gnd.n5591 9.3005
R12191 gnd.n3209 gnd.n3208 9.3005
R12192 gnd.n5655 gnd.n5654 9.3005
R12193 gnd.n5656 gnd.n3206 9.3005
R12194 gnd.n5668 gnd.n5667 9.3005
R12195 gnd.n5666 gnd.n3207 9.3005
R12196 gnd.n5665 gnd.n5664 9.3005
R12197 gnd.n5663 gnd.n5657 9.3005
R12198 gnd.n5662 gnd.n5661 9.3005
R12199 gnd.n5660 gnd.n63 9.3005
R12200 gnd.n4997 gnd.n4996 9.3005
R12201 gnd.n7546 gnd.n64 9.3005
R12202 gnd.t152 gnd.n1065 9.24152
R12203 gnd.n969 gnd.t179 9.24152
R12204 gnd.n2237 gnd.t273 9.24152
R12205 gnd.n4302 gnd.t54 9.24152
R12206 gnd.n6030 gnd.n2885 9.24152
R12207 gnd.n5384 gnd.n3267 9.24152
R12208 gnd.n5601 gnd.t81 9.24152
R12209 gnd.t120 gnd.t152 8.92286
R12210 gnd.n4630 gnd.n3551 8.92286
R12211 gnd.n4676 gnd.n3521 8.92286
R12212 gnd.n4801 gnd.n3455 8.92286
R12213 gnd.n4871 gnd.n4870 8.92286
R12214 gnd.n5227 gnd.n3310 8.92286
R12215 gnd.n5224 gnd.t242 8.92286
R12216 gnd.n2207 gnd.n2182 8.92171
R12217 gnd.n2175 gnd.n2150 8.92171
R12218 gnd.n2143 gnd.n2118 8.92171
R12219 gnd.n2112 gnd.n2087 8.92171
R12220 gnd.n2080 gnd.n2055 8.92171
R12221 gnd.n2048 gnd.n2023 8.92171
R12222 gnd.n2016 gnd.n1991 8.92171
R12223 gnd.n1985 gnd.n1960 8.92171
R12224 gnd.n5249 gnd.n5231 8.72777
R12225 gnd.n1709 gnd.t47 8.60421
R12226 gnd.n1129 gnd.n1117 8.43656
R12227 gnd.n38 gnd.n26 8.43656
R12228 gnd.n4606 gnd.n3566 8.28555
R12229 gnd.n4697 gnd.n3504 8.28555
R12230 gnd.n4780 gnd.n3469 8.28555
R12231 gnd.n4836 gnd.n3422 8.28555
R12232 gnd.n2208 gnd.n2180 8.14595
R12233 gnd.n2176 gnd.n2148 8.14595
R12234 gnd.n2144 gnd.n2116 8.14595
R12235 gnd.n2113 gnd.n2085 8.14595
R12236 gnd.n2081 gnd.n2053 8.14595
R12237 gnd.n2049 gnd.n2021 8.14595
R12238 gnd.n2017 gnd.n1989 8.14595
R12239 gnd.n1986 gnd.n1958 8.14595
R12240 gnd.n4259 gnd.n0 8.10675
R12241 gnd.n7547 gnd.n7546 8.10675
R12242 gnd.n2213 gnd.n2212 7.97301
R12243 gnd.t20 gnd.n1224 7.9669
R12244 gnd.n7547 gnd.n62 7.78567
R12245 gnd.n5158 gnd.n5009 7.75808
R12246 gnd.n6088 gnd.n6087 7.75808
R12247 gnd.n7472 gnd.n182 7.75808
R12248 gnd.n3873 gnd.n3866 7.75808
R12249 gnd.n4513 gnd.n4512 7.64824
R12250 gnd.n4606 gnd.n3565 7.64824
R12251 gnd.t149 gnd.n4650 7.64824
R12252 gnd.n4698 gnd.t151 7.64824
R12253 gnd.n4708 gnd.n3504 7.64824
R12254 gnd.n4780 gnd.n3468 7.64824
R12255 gnd.t32 gnd.n3463 7.64824
R12256 gnd.n4800 gnd.t93 7.64824
R12257 gnd.n4836 gnd.n3413 7.64824
R12258 gnd.n4945 gnd.n3376 7.64824
R12259 gnd.n1154 gnd.n1153 7.53171
R12260 gnd.n1618 gnd.t66 7.32958
R12261 gnd.n2907 gnd.n2906 7.30353
R12262 gnd.n5248 gnd.n5247 7.30353
R12263 gnd.n1578 gnd.n1297 7.01093
R12264 gnd.n1300 gnd.n1298 7.01093
R12265 gnd.n1588 gnd.n1587 7.01093
R12266 gnd.n1599 gnd.n1281 7.01093
R12267 gnd.n1598 gnd.n1284 7.01093
R12268 gnd.n1609 gnd.n1272 7.01093
R12269 gnd.n1275 gnd.n1273 7.01093
R12270 gnd.n1619 gnd.n1618 7.01093
R12271 gnd.n1629 gnd.n1253 7.01093
R12272 gnd.n1628 gnd.n1256 7.01093
R12273 gnd.n1637 gnd.n1247 7.01093
R12274 gnd.n1649 gnd.n1237 7.01093
R12275 gnd.n1659 gnd.n1222 7.01093
R12276 gnd.n1675 gnd.n1674 7.01093
R12277 gnd.n1224 gnd.n1161 7.01093
R12278 gnd.n1729 gnd.n1162 7.01093
R12279 gnd.n1723 gnd.n1722 7.01093
R12280 gnd.n1211 gnd.n1173 7.01093
R12281 gnd.n1715 gnd.n1184 7.01093
R12282 gnd.n1202 gnd.n1197 7.01093
R12283 gnd.n1709 gnd.n1708 7.01093
R12284 gnd.n1755 gnd.n1100 7.01093
R12285 gnd.n1754 gnd.n1753 7.01093
R12286 gnd.n1766 gnd.n1765 7.01093
R12287 gnd.n1093 gnd.n1085 7.01093
R12288 gnd.n1795 gnd.n1073 7.01093
R12289 gnd.n1794 gnd.n1076 7.01093
R12290 gnd.n1805 gnd.n1065 7.01093
R12291 gnd.n1066 gnd.n1054 7.01093
R12292 gnd.n1816 gnd.n1055 7.01093
R12293 gnd.n1842 gnd.n1047 7.01093
R12294 gnd.n1841 gnd.n1840 7.01093
R12295 gnd.n1864 gnd.n1863 7.01093
R12296 gnd.n1882 gnd.n1020 7.01093
R12297 gnd.n1881 gnd.n1023 7.01093
R12298 gnd.n1892 gnd.n1012 7.01093
R12299 gnd.n1013 gnd.n1000 7.01093
R12300 gnd.n1903 gnd.n1001 7.01093
R12301 gnd.n1930 gnd.n985 7.01093
R12302 gnd.n1942 gnd.n1941 7.01093
R12303 gnd.n1924 gnd.n978 7.01093
R12304 gnd.n1953 gnd.n1952 7.01093
R12305 gnd.n2225 gnd.n966 7.01093
R12306 gnd.n2224 gnd.n969 7.01093
R12307 gnd.n2237 gnd.n958 7.01093
R12308 gnd.n959 gnd.n951 7.01093
R12309 gnd.n2247 gnd.n877 7.01093
R12310 gnd.n5959 gnd.n2914 7.01093
R12311 gnd.n4630 gnd.n4629 7.01093
R12312 gnd.n4651 gnd.t149 7.01093
R12313 gnd.n4650 gnd.n3521 7.01093
R12314 gnd.n4801 gnd.n4800 7.01093
R12315 gnd.t93 gnd.n4798 7.01093
R12316 gnd.n4871 gnd.n3426 7.01093
R12317 gnd.n5227 gnd.n5226 7.01093
R12318 gnd.t242 gnd.n3304 7.01093
R12319 gnd.n1256 gnd.t298 6.69227
R12320 gnd.n1076 gnd.t120 6.69227
R12321 gnd.n1840 gnd.n870 6.69227
R12322 gnd.n1931 gnd.t299 6.69227
R12323 gnd.n3378 gnd.t308 6.69227
R12324 gnd.n5378 gnd.n5377 6.5566
R12325 gnd.n3615 gnd.n3614 6.5566
R12326 gnd.n5971 gnd.n5967 6.5566
R12327 gnd.n5256 gnd.n5255 6.5566
R12328 gnd.n4466 gnd.t215 6.37362
R12329 gnd.n4519 gnd.n3589 6.37362
R12330 gnd.n4574 gnd.n3580 6.37362
R12331 gnd.n4658 gnd.t31 6.37362
R12332 gnd.n4716 gnd.n3498 6.37362
R12333 gnd.n4728 gnd.n3485 6.37362
R12334 gnd.n4849 gnd.t30 6.37362
R12335 gnd.n4897 gnd.n3409 6.37362
R12336 gnd.n4820 gnd.n3396 6.37362
R12337 gnd.t201 gnd.n3383 6.37362
R12338 gnd.n2668 gnd.n2666 6.20656
R12339 gnd.n5161 gnd.n5004 6.20656
R12340 gnd.t111 gnd.n1685 6.05496
R12341 gnd.n1686 gnd.t156 6.05496
R12342 gnd.t8 gnd.n1100 6.05496
R12343 gnd.t155 gnd.n1852 6.05496
R12344 gnd.n4167 gnd.t187 6.05496
R12345 gnd.t63 gnd.t225 6.05496
R12346 gnd.t19 gnd.t117 6.05496
R12347 gnd.t12 gnd.t314 6.05496
R12348 gnd.n176 gnd.t175 6.05496
R12349 gnd.n2210 gnd.n2180 5.81868
R12350 gnd.n2178 gnd.n2148 5.81868
R12351 gnd.n2146 gnd.n2116 5.81868
R12352 gnd.n2115 gnd.n2085 5.81868
R12353 gnd.n2083 gnd.n2053 5.81868
R12354 gnd.n2051 gnd.n2021 5.81868
R12355 gnd.n2019 gnd.n1989 5.81868
R12356 gnd.n1988 gnd.n1958 5.81868
R12357 gnd.n3546 gnd.n3534 5.73631
R12358 gnd.n4641 gnd.n3527 5.73631
R12359 gnd.t151 gnd.n4697 5.73631
R12360 gnd.n3469 gnd.t32 5.73631
R12361 gnd.n4738 gnd.n4737 5.73631
R12362 gnd.n4808 gnd.n3444 5.73631
R12363 gnd.n5387 gnd.n3263 5.62001
R12364 gnd.n6033 gnd.n2850 5.62001
R12365 gnd.n6033 gnd.n2851 5.62001
R12366 gnd.n5387 gnd.n3264 5.62001
R12367 gnd.n1437 gnd.n1432 5.4308
R12368 gnd.n2255 gnd.n944 5.4308
R12369 gnd.n1753 gnd.t67 5.41765
R12370 gnd.t154 gnd.n1776 5.41765
R12371 gnd.t37 gnd.n1032 5.41765
R12372 gnd.t87 gnd.n4589 5.41765
R12373 gnd.n4828 gnd.t115 5.41765
R12374 gnd.n4496 gnd.t215 5.09899
R12375 gnd.t252 gnd.n3584 5.09899
R12376 gnd.n4582 gnd.n3584 5.09899
R12377 gnd.n4756 gnd.n3489 5.09899
R12378 gnd.n4764 gnd.n3482 5.09899
R12379 gnd.n4923 gnd.n3393 5.09899
R12380 gnd.n2208 gnd.n2207 5.04292
R12381 gnd.n2176 gnd.n2175 5.04292
R12382 gnd.n2144 gnd.n2143 5.04292
R12383 gnd.n2113 gnd.n2112 5.04292
R12384 gnd.n2081 gnd.n2080 5.04292
R12385 gnd.n2049 gnd.n2048 5.04292
R12386 gnd.n2017 gnd.n2016 5.04292
R12387 gnd.n1986 gnd.n1985 5.04292
R12388 gnd.n1716 gnd.t296 4.78034
R12389 gnd.n1055 gnd.t21 4.78034
R12390 gnd.n4423 gnd.t304 4.78034
R12391 gnd.n5193 gnd.t312 4.78034
R12392 gnd.n1158 gnd.n1155 4.74817
R12393 gnd.n1208 gnd.n1106 4.74817
R12394 gnd.n1195 gnd.n1105 4.74817
R12395 gnd.n1104 gnd.n1103 4.74817
R12396 gnd.n1204 gnd.n1155 4.74817
R12397 gnd.n1205 gnd.n1106 4.74817
R12398 gnd.n1207 gnd.n1105 4.74817
R12399 gnd.n1194 gnd.n1104 4.74817
R12400 gnd.n3110 gnd.n82 4.74817
R12401 gnd.n5779 gnd.n81 4.74817
R12402 gnd.n3127 gnd.n80 4.74817
R12403 gnd.n7539 gnd.n75 4.74817
R12404 gnd.n7537 gnd.n76 4.74817
R12405 gnd.n5793 gnd.n82 4.74817
R12406 gnd.n3109 gnd.n81 4.74817
R12407 gnd.n5780 gnd.n80 4.74817
R12408 gnd.n3126 gnd.n75 4.74817
R12409 gnd.n7538 gnd.n7537 4.74817
R12410 gnd.n3795 gnd.n3792 4.74817
R12411 gnd.n3799 gnd.n3791 4.74817
R12412 gnd.n4238 gnd.n3790 4.74817
R12413 gnd.n4236 gnd.n3789 4.74817
R12414 gnd.n4232 gnd.n3788 4.74817
R12415 gnd.n5788 gnd.n3116 4.74817
R12416 gnd.n5786 gnd.n5785 4.74817
R12417 gnd.n3141 gnd.n3140 4.74817
R12418 gnd.n3146 gnd.n3145 4.74817
R12419 gnd.n5766 gnd.n5765 4.74817
R12420 gnd.n5635 gnd.n3116 4.74817
R12421 gnd.n5787 gnd.n5786 4.74817
R12422 gnd.n3140 gnd.n3117 4.74817
R12423 gnd.n3145 gnd.n3144 4.74817
R12424 gnd.n5767 gnd.n5766 4.74817
R12425 gnd.n6245 gnd.n6244 4.74817
R12426 gnd.n2471 gnd.n2455 4.74817
R12427 gnd.n6232 gnd.n6231 4.74817
R12428 gnd.n2488 gnd.n2472 4.74817
R12429 gnd.n6219 gnd.n6218 4.74817
R12430 gnd.n6246 gnd.n6245 4.74817
R12431 gnd.n6243 gnd.n2455 4.74817
R12432 gnd.n6233 gnd.n6232 4.74817
R12433 gnd.n6230 gnd.n2472 4.74817
R12434 gnd.n6220 gnd.n6219 4.74817
R12435 gnd.n4269 gnd.n3792 4.74817
R12436 gnd.n4268 gnd.n3791 4.74817
R12437 gnd.n3798 gnd.n3790 4.74817
R12438 gnd.n4239 gnd.n3789 4.74817
R12439 gnd.n4235 gnd.n3788 4.74817
R12440 gnd.n1153 gnd.n1152 4.74296
R12441 gnd.n62 gnd.n61 4.74296
R12442 gnd.n1129 gnd.n1128 4.7074
R12443 gnd.n1141 gnd.n1140 4.7074
R12444 gnd.n38 gnd.n37 4.7074
R12445 gnd.n50 gnd.n49 4.7074
R12446 gnd.n1153 gnd.n1141 4.65959
R12447 gnd.n62 gnd.n50 4.65959
R12448 gnd.n5478 gnd.n5388 4.6132
R12449 gnd.n6034 gnd.n2849 4.6132
R12450 gnd.n4496 gnd.n4495 4.46168
R12451 gnd.t172 gnd.n2914 4.46168
R12452 gnd.n4502 gnd.t172 4.46168
R12453 gnd.n4627 gnd.t291 4.46168
R12454 gnd.n4638 gnd.n4636 4.46168
R12455 gnd.n4667 gnd.n3529 4.46168
R12456 gnd.n4815 gnd.n3449 4.46168
R12457 gnd.n4859 gnd.n3436 4.46168
R12458 gnd.t92 gnd.n4857 4.46168
R12459 gnd.n5317 gnd.n3304 4.46168
R12460 gnd.n5244 gnd.n5231 4.46111
R12461 gnd.n2193 gnd.n2189 4.38594
R12462 gnd.n2161 gnd.n2157 4.38594
R12463 gnd.n2129 gnd.n2125 4.38594
R12464 gnd.n2098 gnd.n2094 4.38594
R12465 gnd.n2066 gnd.n2062 4.38594
R12466 gnd.n2034 gnd.n2030 4.38594
R12467 gnd.n2002 gnd.n1998 4.38594
R12468 gnd.n1971 gnd.n1967 4.38594
R12469 gnd.n2204 gnd.n2182 4.26717
R12470 gnd.n2172 gnd.n2150 4.26717
R12471 gnd.n2140 gnd.n2118 4.26717
R12472 gnd.n2109 gnd.n2087 4.26717
R12473 gnd.n2077 gnd.n2055 4.26717
R12474 gnd.n2045 gnd.n2023 4.26717
R12475 gnd.n2013 gnd.n1991 4.26717
R12476 gnd.n1982 gnd.n1960 4.26717
R12477 gnd.n1660 gnd.t300 4.14303
R12478 gnd.n1892 gnd.t48 4.14303
R12479 gnd.t211 gnd.n2564 4.14303
R12480 gnd.t194 gnd.n3032 4.14303
R12481 gnd.n2212 gnd.n2211 4.08274
R12482 gnd.n5377 gnd.n5376 4.05904
R12483 gnd.n3616 gnd.n3615 4.05904
R12484 gnd.n5974 gnd.n5967 4.05904
R12485 gnd.n5257 gnd.n5256 4.05904
R12486 gnd.n15 gnd.n7 3.99943
R12487 gnd.n1733 gnd.n1154 3.9165
R12488 gnd.n6030 gnd.t75 3.82437
R12489 gnd.n4538 gnd.n3597 3.82437
R12490 gnd.n4580 gnd.t58 3.82437
R12491 gnd.n4599 gnd.n4598 3.82437
R12492 gnd.n4687 gnd.n3518 3.82437
R12493 gnd.n4689 gnd.t19 3.82437
R12494 gnd.n4730 gnd.t12 3.82437
R12495 gnd.n4773 gnd.n4772 3.82437
R12496 gnd.n4888 gnd.n3407 3.82437
R12497 gnd.n4914 gnd.t11 3.82437
R12498 gnd.n4938 gnd.n4937 3.82437
R12499 gnd.n5384 gnd.t310 3.82437
R12500 gnd.n1141 gnd.n1129 3.72967
R12501 gnd.n50 gnd.n38 3.72967
R12502 gnd.n2212 gnd.n2084 3.70378
R12503 gnd.n15 gnd.n14 3.60163
R12504 gnd.n2203 gnd.n2184 3.49141
R12505 gnd.n2171 gnd.n2152 3.49141
R12506 gnd.n2139 gnd.n2120 3.49141
R12507 gnd.n2108 gnd.n2089 3.49141
R12508 gnd.n2076 gnd.n2057 3.49141
R12509 gnd.n2044 gnd.n2025 3.49141
R12510 gnd.n2012 gnd.n1993 3.49141
R12511 gnd.n1981 gnd.n1962 3.49141
R12512 gnd.n5459 gnd.n5458 3.29747
R12513 gnd.n5458 gnd.n5396 3.29747
R12514 gnd.n7436 gnd.n7433 3.29747
R12515 gnd.n7437 gnd.n7436 3.29747
R12516 gnd.n4016 gnd.n3957 3.29747
R12517 gnd.n3957 gnd.n3952 3.29747
R12518 gnd.n6052 gnd.n6051 3.29747
R12519 gnd.n6051 gnd.n6050 3.29747
R12520 gnd.n4503 gnd.n3604 3.18706
R12521 gnd.n4616 gnd.n4615 3.18706
R12522 gnd.n4678 gnd.n4677 3.18706
R12523 gnd.n4788 gnd.n4787 3.18706
R12524 gnd.n4869 gnd.n4868 3.18706
R12525 gnd.n4820 gnd.t201 3.18706
R12526 gnd.n4955 gnd.n4953 3.18706
R12527 gnd.n1239 gnd.t300 2.8684
R12528 gnd.n3681 gnd.t75 2.8684
R12529 gnd.n1142 gnd.t70 2.82907
R12530 gnd.n1142 gnd.t50 2.82907
R12531 gnd.n1144 gnd.t5 2.82907
R12532 gnd.n1144 gnd.t162 2.82907
R12533 gnd.n1146 gnd.t65 2.82907
R12534 gnd.n1146 gnd.t18 2.82907
R12535 gnd.n1148 gnd.t53 2.82907
R12536 gnd.n1148 gnd.t99 2.82907
R12537 gnd.n1150 gnd.t147 2.82907
R12538 gnd.n1150 gnd.t42 2.82907
R12539 gnd.n1107 gnd.t97 2.82907
R12540 gnd.n1107 gnd.t114 2.82907
R12541 gnd.n1109 gnd.t86 2.82907
R12542 gnd.n1109 gnd.t80 2.82907
R12543 gnd.n1111 gnd.t101 2.82907
R12544 gnd.n1111 gnd.t79 2.82907
R12545 gnd.n1113 gnd.t59 2.82907
R12546 gnd.n1113 gnd.t96 2.82907
R12547 gnd.n1115 gnd.t107 2.82907
R12548 gnd.n1115 gnd.t100 2.82907
R12549 gnd.n1118 gnd.t104 2.82907
R12550 gnd.n1118 gnd.t168 2.82907
R12551 gnd.n1120 gnd.t27 2.82907
R12552 gnd.n1120 gnd.t57 2.82907
R12553 gnd.n1122 gnd.t44 2.82907
R12554 gnd.n1122 gnd.t72 2.82907
R12555 gnd.n1124 gnd.t60 2.82907
R12556 gnd.n1124 gnd.t166 2.82907
R12557 gnd.n1126 gnd.t74 2.82907
R12558 gnd.n1126 gnd.t297 2.82907
R12559 gnd.n1130 gnd.t91 2.82907
R12560 gnd.n1130 gnd.t24 2.82907
R12561 gnd.n1132 gnd.t293 2.82907
R12562 gnd.n1132 gnd.t163 2.82907
R12563 gnd.n1134 gnd.t83 2.82907
R12564 gnd.n1134 gnd.t130 2.82907
R12565 gnd.n1136 gnd.t16 2.82907
R12566 gnd.n1136 gnd.t158 2.82907
R12567 gnd.n1138 gnd.t295 2.82907
R12568 gnd.n1138 gnd.t123 2.82907
R12569 gnd.n59 gnd.t303 2.82907
R12570 gnd.n59 gnd.t294 2.82907
R12571 gnd.n57 gnd.t85 2.82907
R12572 gnd.n57 gnd.t3 2.82907
R12573 gnd.n55 gnd.t84 2.82907
R12574 gnd.n55 gnd.t98 2.82907
R12575 gnd.n53 gnd.t49 2.82907
R12576 gnd.n53 gnd.t140 2.82907
R12577 gnd.n51 gnd.t46 2.82907
R12578 gnd.n51 gnd.t94 2.82907
R12579 gnd.n24 gnd.t160 2.82907
R12580 gnd.n24 gnd.t26 2.82907
R12581 gnd.n22 gnd.t167 2.82907
R12582 gnd.n22 gnd.t108 2.82907
R12583 gnd.n20 gnd.t62 2.82907
R12584 gnd.n20 gnd.t113 2.82907
R12585 gnd.n18 gnd.t170 2.82907
R12586 gnd.n18 gnd.t132 2.82907
R12587 gnd.n16 gnd.t139 2.82907
R12588 gnd.n16 gnd.t14 2.82907
R12589 gnd.n35 gnd.t136 2.82907
R12590 gnd.n35 gnd.t145 2.82907
R12591 gnd.n33 gnd.t36 2.82907
R12592 gnd.n33 gnd.t150 2.82907
R12593 gnd.n31 gnd.t306 2.82907
R12594 gnd.n31 gnd.t71 2.82907
R12595 gnd.n29 gnd.t7 2.82907
R12596 gnd.n29 gnd.t318 2.82907
R12597 gnd.n27 gnd.t169 2.82907
R12598 gnd.n27 gnd.t165 2.82907
R12599 gnd.n47 gnd.t110 2.82907
R12600 gnd.n47 gnd.t164 2.82907
R12601 gnd.n45 gnd.t292 2.82907
R12602 gnd.n45 gnd.t119 2.82907
R12603 gnd.n43 gnd.t128 2.82907
R12604 gnd.n43 gnd.t34 2.82907
R12605 gnd.n41 gnd.t131 2.82907
R12606 gnd.n41 gnd.t52 2.82907
R12607 gnd.n39 gnd.t159 2.82907
R12608 gnd.n39 gnd.t302 2.82907
R12609 gnd.n2200 gnd.n2199 2.71565
R12610 gnd.n2168 gnd.n2167 2.71565
R12611 gnd.n2136 gnd.n2135 2.71565
R12612 gnd.n2105 gnd.n2104 2.71565
R12613 gnd.n2073 gnd.n2072 2.71565
R12614 gnd.n2041 gnd.n2040 2.71565
R12615 gnd.n2009 gnd.n2008 2.71565
R12616 gnd.n1978 gnd.n1977 2.71565
R12617 gnd.n4528 gnd.n4527 2.54975
R12618 gnd.n4617 gnd.n3560 2.54975
R12619 gnd.n4617 gnd.t144 2.54975
R12620 gnd.n4698 gnd.n3511 2.54975
R12621 gnd.n4789 gnd.n3463 2.54975
R12622 gnd.n4878 gnd.t10 2.54975
R12623 gnd.n4878 gnd.n4877 2.54975
R12624 gnd.n3379 gnd.n3372 2.54975
R12625 gnd.n1733 gnd.n1155 2.27742
R12626 gnd.n1733 gnd.n1106 2.27742
R12627 gnd.n1733 gnd.n1105 2.27742
R12628 gnd.n1733 gnd.n1104 2.27742
R12629 gnd.n7536 gnd.n82 2.27742
R12630 gnd.n7536 gnd.n81 2.27742
R12631 gnd.n7536 gnd.n80 2.27742
R12632 gnd.n7536 gnd.n75 2.27742
R12633 gnd.n7537 gnd.n7536 2.27742
R12634 gnd.n3116 gnd.n79 2.27742
R12635 gnd.n5786 gnd.n79 2.27742
R12636 gnd.n3140 gnd.n79 2.27742
R12637 gnd.n3145 gnd.n79 2.27742
R12638 gnd.n5766 gnd.n79 2.27742
R12639 gnd.n6245 gnd.n2454 2.27742
R12640 gnd.n2455 gnd.n2454 2.27742
R12641 gnd.n6232 gnd.n2454 2.27742
R12642 gnd.n2472 gnd.n2454 2.27742
R12643 gnd.n6219 gnd.n2454 2.27742
R12644 gnd.n4275 gnd.n3792 2.27742
R12645 gnd.n4275 gnd.n3791 2.27742
R12646 gnd.n4275 gnd.n3790 2.27742
R12647 gnd.n4275 gnd.n3789 2.27742
R12648 gnd.n4275 gnd.n3788 2.27742
R12649 gnd.n1587 gnd.t245 2.23109
R12650 gnd.n1210 gnd.t296 2.23109
R12651 gnd.t105 gnd.n3529 2.23109
R12652 gnd.t117 gnd.n4687 2.23109
R12653 gnd.n4773 gnd.t314 2.23109
R12654 gnd.t77 gnd.n3449 2.23109
R12655 gnd.n2196 gnd.n2186 1.93989
R12656 gnd.n2164 gnd.n2154 1.93989
R12657 gnd.n2132 gnd.n2122 1.93989
R12658 gnd.n2101 gnd.n2091 1.93989
R12659 gnd.n2069 gnd.n2059 1.93989
R12660 gnd.n2037 gnd.n2027 1.93989
R12661 gnd.n2005 gnd.n1995 1.93989
R12662 gnd.n1974 gnd.n1964 1.93989
R12663 gnd.n4539 gnd.n3596 1.91244
R12664 gnd.t289 gnd.n3597 1.91244
R12665 gnd.n4548 gnd.n4546 1.91244
R12666 gnd.n4707 gnd.n3506 1.91244
R12667 gnd.n3476 gnd.n3475 1.91244
R12668 gnd.n4891 gnd.n4890 1.91244
R12669 gnd.n3386 gnd.n3385 1.91244
R12670 gnd.n5218 gnd.t283 1.91244
R12671 gnd.t28 gnd.n1598 1.59378
R12672 gnd.n1777 gnd.t154 1.59378
R12673 gnd.n1040 gnd.t37 1.59378
R12674 gnd.t89 gnd.n3551 1.59378
R12675 gnd.n4870 gnd.t102 1.59378
R12676 gnd.n5960 gnd.n2911 1.27512
R12677 gnd.n4513 gnd.t207 1.27512
R12678 gnd.n4590 gnd.t58 1.27512
R12679 gnd.n4628 gnd.n4627 1.27512
R12680 gnd.n4651 gnd.n3538 1.27512
R12681 gnd.n4798 gnd.n4797 1.27512
R12682 gnd.n4857 gnd.n3437 1.27512
R12683 gnd.n4827 gnd.t11 1.27512
R12684 gnd.t198 gnd.n3376 1.27512
R12685 gnd.n4945 gnd.t228 1.27512
R12686 gnd.n5225 gnd.n5224 1.27512
R12687 gnd.n1440 gnd.n1432 1.16414
R12688 gnd.n2258 gnd.n944 1.16414
R12689 gnd.n2195 gnd.n2188 1.16414
R12690 gnd.n2163 gnd.n2156 1.16414
R12691 gnd.n2131 gnd.n2124 1.16414
R12692 gnd.n2100 gnd.n2093 1.16414
R12693 gnd.n2068 gnd.n2061 1.16414
R12694 gnd.n2036 gnd.n2029 1.16414
R12695 gnd.n2004 gnd.n1997 1.16414
R12696 gnd.n1973 gnd.n1966 1.16414
R12697 gnd.n5388 gnd.n3262 0.970197
R12698 gnd.n6034 gnd.n2751 0.970197
R12699 gnd.n2179 gnd.n2147 0.962709
R12700 gnd.n2211 gnd.n2179 0.962709
R12701 gnd.n2052 gnd.n2020 0.962709
R12702 gnd.n2084 gnd.n2052 0.962709
R12703 gnd.n1686 gnd.t111 0.956468
R12704 gnd.n1853 gnd.t155 0.956468
R12705 gnd.t126 gnd.n2400 0.956468
R12706 gnd.n4142 gnd.t73 0.956468
R12707 gnd.n4332 gnd.t69 0.956468
R12708 gnd.n4298 gnd.t23 0.956468
R12709 gnd.t134 gnd.n3698 0.956468
R12710 gnd.t283 gnd.t310 0.956468
R12711 gnd.n5206 gnd.t316 0.956468
R12712 gnd.n5589 gnd.t45 0.956468
R12713 gnd.n5644 gnd.t13 0.956468
R12714 gnd.n5749 gnd.t25 0.956468
R12715 gnd.t0 gnd.n138 0.956468
R12716 gnd.n2 gnd.n1 0.672012
R12717 gnd.n3 gnd.n2 0.672012
R12718 gnd.n4 gnd.n3 0.672012
R12719 gnd.n5 gnd.n4 0.672012
R12720 gnd.n6 gnd.n5 0.672012
R12721 gnd.n7 gnd.n6 0.672012
R12722 gnd.n9 gnd.n8 0.672012
R12723 gnd.n10 gnd.n9 0.672012
R12724 gnd.n11 gnd.n10 0.672012
R12725 gnd.n12 gnd.n11 0.672012
R12726 gnd.n13 gnd.n12 0.672012
R12727 gnd.n14 gnd.n13 0.672012
R12728 gnd.t225 gnd.n3606 0.637812
R12729 gnd.n4569 gnd.n4568 0.637812
R12730 gnd.n4589 gnd.n4588 0.637812
R12731 gnd.n4598 gnd.t143 0.637812
R12732 gnd.n4718 gnd.n4717 0.637812
R12733 gnd.n4763 gnd.n4762 0.637812
R12734 gnd.t125 gnd.n4888 0.637812
R12735 gnd.n4829 gnd.n4828 0.637812
R12736 gnd.n4922 gnd.n4920 0.637812
R12737 gnd.n4953 gnd.t267 0.637812
R12738 gnd.n1152 gnd.n1151 0.573776
R12739 gnd.n1151 gnd.n1149 0.573776
R12740 gnd.n1149 gnd.n1147 0.573776
R12741 gnd.n1147 gnd.n1145 0.573776
R12742 gnd.n1145 gnd.n1143 0.573776
R12743 gnd.n1117 gnd.n1116 0.573776
R12744 gnd.n1116 gnd.n1114 0.573776
R12745 gnd.n1114 gnd.n1112 0.573776
R12746 gnd.n1112 gnd.n1110 0.573776
R12747 gnd.n1110 gnd.n1108 0.573776
R12748 gnd.n1128 gnd.n1127 0.573776
R12749 gnd.n1127 gnd.n1125 0.573776
R12750 gnd.n1125 gnd.n1123 0.573776
R12751 gnd.n1123 gnd.n1121 0.573776
R12752 gnd.n1121 gnd.n1119 0.573776
R12753 gnd.n1140 gnd.n1139 0.573776
R12754 gnd.n1139 gnd.n1137 0.573776
R12755 gnd.n1137 gnd.n1135 0.573776
R12756 gnd.n1135 gnd.n1133 0.573776
R12757 gnd.n1133 gnd.n1131 0.573776
R12758 gnd.n54 gnd.n52 0.573776
R12759 gnd.n56 gnd.n54 0.573776
R12760 gnd.n58 gnd.n56 0.573776
R12761 gnd.n60 gnd.n58 0.573776
R12762 gnd.n61 gnd.n60 0.573776
R12763 gnd.n19 gnd.n17 0.573776
R12764 gnd.n21 gnd.n19 0.573776
R12765 gnd.n23 gnd.n21 0.573776
R12766 gnd.n25 gnd.n23 0.573776
R12767 gnd.n26 gnd.n25 0.573776
R12768 gnd.n30 gnd.n28 0.573776
R12769 gnd.n32 gnd.n30 0.573776
R12770 gnd.n34 gnd.n32 0.573776
R12771 gnd.n36 gnd.n34 0.573776
R12772 gnd.n37 gnd.n36 0.573776
R12773 gnd.n42 gnd.n40 0.573776
R12774 gnd.n44 gnd.n42 0.573776
R12775 gnd.n46 gnd.n44 0.573776
R12776 gnd.n48 gnd.n46 0.573776
R12777 gnd.n49 gnd.n48 0.573776
R12778 gnd gnd.n0 0.551497
R12779 gnd.n7474 gnd.n7473 0.532512
R12780 gnd.n3869 gnd.n3868 0.532512
R12781 gnd.n7289 gnd.n166 0.497451
R12782 gnd.n2723 gnd.n2569 0.497451
R12783 gnd.n5414 gnd.n3027 0.497451
R12784 gnd.n3972 gnd.n2370 0.497451
R12785 gnd.n5170 gnd.n5169 0.489829
R12786 gnd.n4386 gnd.n2582 0.489829
R12787 gnd.n4377 gnd.n2605 0.489829
R12788 gnd.n5056 gnd.n2998 0.489829
R12789 gnd.n1915 gnd.n948 0.486781
R12790 gnd.n1489 gnd.n1488 0.48678
R12791 gnd.n2232 gnd.n902 0.480683
R12792 gnd.n1573 gnd.n1572 0.480683
R12793 gnd.n7548 gnd.n7547 0.470187
R12794 gnd.n6497 gnd.n6496 0.468488
R12795 gnd.n7018 gnd.n7017 0.468488
R12796 gnd.n7229 gnd.n7228 0.468488
R12797 gnd.n6326 gnd.n6325 0.468488
R12798 gnd.n7536 gnd.n79 0.4255
R12799 gnd.n4275 gnd.n2454 0.4255
R12800 gnd.n6092 gnd.n2666 0.388379
R12801 gnd.n2192 gnd.n2191 0.388379
R12802 gnd.n2160 gnd.n2159 0.388379
R12803 gnd.n2128 gnd.n2127 0.388379
R12804 gnd.n2097 gnd.n2096 0.388379
R12805 gnd.n2065 gnd.n2064 0.388379
R12806 gnd.n2033 gnd.n2032 0.388379
R12807 gnd.n2001 gnd.n2000 0.388379
R12808 gnd.n1970 gnd.n1969 0.388379
R12809 gnd.n5147 gnd.n5004 0.388379
R12810 gnd.n7548 gnd.n15 0.374463
R12811 gnd.n1003 gnd.t299 0.319156
R12812 gnd.t15 gnd.n2441 0.319156
R12813 gnd.n4220 gnd.t95 0.319156
R12814 gnd.n4241 gnd.t17 0.319156
R12815 gnd.n4251 gnd.t4 0.319156
R12816 gnd.n4393 gnd.t238 0.319156
R12817 gnd.t207 gnd.t63 0.319156
R12818 gnd.t308 gnd.t228 0.319156
R12819 gnd.t218 gnd.n5180 0.319156
R12820 gnd.n5791 gnd.t51 0.319156
R12821 gnd.n5783 gnd.t61 0.319156
R12822 gnd.n5697 gnd.t35 0.319156
R12823 gnd.t2 gnd.n98 0.319156
R12824 gnd.n1407 gnd.n1385 0.311721
R12825 gnd.n6156 gnd.n6155 0.302329
R12826 gnd.n4998 gnd.n4997 0.302329
R12827 gnd gnd.n7548 0.295112
R12828 gnd.n201 gnd.n174 0.293183
R12829 gnd.n4122 gnd.n3909 0.293183
R12830 gnd.n2303 gnd.n2302 0.268793
R12831 gnd.n7350 gnd.n174 0.258122
R12832 gnd.n5564 gnd.n5563 0.258122
R12833 gnd.n2784 gnd.n2577 0.258122
R12834 gnd.n4122 gnd.n4121 0.258122
R12835 gnd.n2302 gnd.n2301 0.241354
R12836 gnd.n5479 gnd.n5478 0.229039
R12837 gnd.n5478 gnd.n3261 0.229039
R12838 gnd.n2849 gnd.n2750 0.229039
R12839 gnd.n2849 gnd.n2848 0.229039
R12840 gnd.n1561 gnd.n1360 0.206293
R12841 gnd.n2209 gnd.n2181 0.155672
R12842 gnd.n2202 gnd.n2181 0.155672
R12843 gnd.n2202 gnd.n2201 0.155672
R12844 gnd.n2201 gnd.n2185 0.155672
R12845 gnd.n2194 gnd.n2185 0.155672
R12846 gnd.n2194 gnd.n2193 0.155672
R12847 gnd.n2177 gnd.n2149 0.155672
R12848 gnd.n2170 gnd.n2149 0.155672
R12849 gnd.n2170 gnd.n2169 0.155672
R12850 gnd.n2169 gnd.n2153 0.155672
R12851 gnd.n2162 gnd.n2153 0.155672
R12852 gnd.n2162 gnd.n2161 0.155672
R12853 gnd.n2145 gnd.n2117 0.155672
R12854 gnd.n2138 gnd.n2117 0.155672
R12855 gnd.n2138 gnd.n2137 0.155672
R12856 gnd.n2137 gnd.n2121 0.155672
R12857 gnd.n2130 gnd.n2121 0.155672
R12858 gnd.n2130 gnd.n2129 0.155672
R12859 gnd.n2114 gnd.n2086 0.155672
R12860 gnd.n2107 gnd.n2086 0.155672
R12861 gnd.n2107 gnd.n2106 0.155672
R12862 gnd.n2106 gnd.n2090 0.155672
R12863 gnd.n2099 gnd.n2090 0.155672
R12864 gnd.n2099 gnd.n2098 0.155672
R12865 gnd.n2082 gnd.n2054 0.155672
R12866 gnd.n2075 gnd.n2054 0.155672
R12867 gnd.n2075 gnd.n2074 0.155672
R12868 gnd.n2074 gnd.n2058 0.155672
R12869 gnd.n2067 gnd.n2058 0.155672
R12870 gnd.n2067 gnd.n2066 0.155672
R12871 gnd.n2050 gnd.n2022 0.155672
R12872 gnd.n2043 gnd.n2022 0.155672
R12873 gnd.n2043 gnd.n2042 0.155672
R12874 gnd.n2042 gnd.n2026 0.155672
R12875 gnd.n2035 gnd.n2026 0.155672
R12876 gnd.n2035 gnd.n2034 0.155672
R12877 gnd.n2018 gnd.n1990 0.155672
R12878 gnd.n2011 gnd.n1990 0.155672
R12879 gnd.n2011 gnd.n2010 0.155672
R12880 gnd.n2010 gnd.n1994 0.155672
R12881 gnd.n2003 gnd.n1994 0.155672
R12882 gnd.n2003 gnd.n2002 0.155672
R12883 gnd.n1987 gnd.n1959 0.155672
R12884 gnd.n1980 gnd.n1959 0.155672
R12885 gnd.n1980 gnd.n1979 0.155672
R12886 gnd.n1979 gnd.n1963 0.155672
R12887 gnd.n1972 gnd.n1963 0.155672
R12888 gnd.n1972 gnd.n1971 0.155672
R12889 gnd.n2334 gnd.n902 0.152939
R12890 gnd.n2334 gnd.n2333 0.152939
R12891 gnd.n2333 gnd.n2332 0.152939
R12892 gnd.n2332 gnd.n904 0.152939
R12893 gnd.n905 gnd.n904 0.152939
R12894 gnd.n906 gnd.n905 0.152939
R12895 gnd.n907 gnd.n906 0.152939
R12896 gnd.n908 gnd.n907 0.152939
R12897 gnd.n909 gnd.n908 0.152939
R12898 gnd.n910 gnd.n909 0.152939
R12899 gnd.n911 gnd.n910 0.152939
R12900 gnd.n912 gnd.n911 0.152939
R12901 gnd.n913 gnd.n912 0.152939
R12902 gnd.n914 gnd.n913 0.152939
R12903 gnd.n2304 gnd.n914 0.152939
R12904 gnd.n2304 gnd.n2303 0.152939
R12905 gnd.n1574 gnd.n1573 0.152939
R12906 gnd.n1574 gnd.n1278 0.152939
R12907 gnd.n1602 gnd.n1278 0.152939
R12908 gnd.n1603 gnd.n1602 0.152939
R12909 gnd.n1604 gnd.n1603 0.152939
R12910 gnd.n1605 gnd.n1604 0.152939
R12911 gnd.n1605 gnd.n1250 0.152939
R12912 gnd.n1632 gnd.n1250 0.152939
R12913 gnd.n1633 gnd.n1632 0.152939
R12914 gnd.n1634 gnd.n1633 0.152939
R12915 gnd.n1634 gnd.n1228 0.152939
R12916 gnd.n1663 gnd.n1228 0.152939
R12917 gnd.n1664 gnd.n1663 0.152939
R12918 gnd.n1665 gnd.n1664 0.152939
R12919 gnd.n1666 gnd.n1665 0.152939
R12920 gnd.n1668 gnd.n1666 0.152939
R12921 gnd.n1668 gnd.n1667 0.152939
R12922 gnd.n1667 gnd.n1177 0.152939
R12923 gnd.n1178 gnd.n1177 0.152939
R12924 gnd.n1179 gnd.n1178 0.152939
R12925 gnd.n1198 gnd.n1179 0.152939
R12926 gnd.n1199 gnd.n1198 0.152939
R12927 gnd.n1199 gnd.n1097 0.152939
R12928 gnd.n1758 gnd.n1097 0.152939
R12929 gnd.n1759 gnd.n1758 0.152939
R12930 gnd.n1760 gnd.n1759 0.152939
R12931 gnd.n1761 gnd.n1760 0.152939
R12932 gnd.n1761 gnd.n1070 0.152939
R12933 gnd.n1798 gnd.n1070 0.152939
R12934 gnd.n1799 gnd.n1798 0.152939
R12935 gnd.n1800 gnd.n1799 0.152939
R12936 gnd.n1801 gnd.n1800 0.152939
R12937 gnd.n1801 gnd.n1044 0.152939
R12938 gnd.n1845 gnd.n1044 0.152939
R12939 gnd.n1846 gnd.n1845 0.152939
R12940 gnd.n1847 gnd.n1846 0.152939
R12941 gnd.n1848 gnd.n1847 0.152939
R12942 gnd.n1848 gnd.n1017 0.152939
R12943 gnd.n1885 gnd.n1017 0.152939
R12944 gnd.n1886 gnd.n1885 0.152939
R12945 gnd.n1887 gnd.n1886 0.152939
R12946 gnd.n1888 gnd.n1887 0.152939
R12947 gnd.n1888 gnd.n990 0.152939
R12948 gnd.n1934 gnd.n990 0.152939
R12949 gnd.n1935 gnd.n1934 0.152939
R12950 gnd.n1936 gnd.n1935 0.152939
R12951 gnd.n1937 gnd.n1936 0.152939
R12952 gnd.n1937 gnd.n963 0.152939
R12953 gnd.n2228 gnd.n963 0.152939
R12954 gnd.n2229 gnd.n2228 0.152939
R12955 gnd.n2230 gnd.n2229 0.152939
R12956 gnd.n2231 gnd.n2230 0.152939
R12957 gnd.n2232 gnd.n2231 0.152939
R12958 gnd.n1572 gnd.n1302 0.152939
R12959 gnd.n1323 gnd.n1302 0.152939
R12960 gnd.n1324 gnd.n1323 0.152939
R12961 gnd.n1330 gnd.n1324 0.152939
R12962 gnd.n1331 gnd.n1330 0.152939
R12963 gnd.n1332 gnd.n1331 0.152939
R12964 gnd.n1332 gnd.n1321 0.152939
R12965 gnd.n1340 gnd.n1321 0.152939
R12966 gnd.n1341 gnd.n1340 0.152939
R12967 gnd.n1342 gnd.n1341 0.152939
R12968 gnd.n1342 gnd.n1319 0.152939
R12969 gnd.n1350 gnd.n1319 0.152939
R12970 gnd.n1351 gnd.n1350 0.152939
R12971 gnd.n1352 gnd.n1351 0.152939
R12972 gnd.n1352 gnd.n1317 0.152939
R12973 gnd.n1360 gnd.n1317 0.152939
R12974 gnd.n2301 gnd.n919 0.152939
R12975 gnd.n921 gnd.n919 0.152939
R12976 gnd.n922 gnd.n921 0.152939
R12977 gnd.n923 gnd.n922 0.152939
R12978 gnd.n924 gnd.n923 0.152939
R12979 gnd.n925 gnd.n924 0.152939
R12980 gnd.n926 gnd.n925 0.152939
R12981 gnd.n927 gnd.n926 0.152939
R12982 gnd.n928 gnd.n927 0.152939
R12983 gnd.n929 gnd.n928 0.152939
R12984 gnd.n930 gnd.n929 0.152939
R12985 gnd.n931 gnd.n930 0.152939
R12986 gnd.n932 gnd.n931 0.152939
R12987 gnd.n933 gnd.n932 0.152939
R12988 gnd.n934 gnd.n933 0.152939
R12989 gnd.n935 gnd.n934 0.152939
R12990 gnd.n936 gnd.n935 0.152939
R12991 gnd.n937 gnd.n936 0.152939
R12992 gnd.n938 gnd.n937 0.152939
R12993 gnd.n939 gnd.n938 0.152939
R12994 gnd.n940 gnd.n939 0.152939
R12995 gnd.n941 gnd.n940 0.152939
R12996 gnd.n945 gnd.n941 0.152939
R12997 gnd.n946 gnd.n945 0.152939
R12998 gnd.n947 gnd.n946 0.152939
R12999 gnd.n948 gnd.n947 0.152939
R13000 gnd.n1735 gnd.n1734 0.152939
R13001 gnd.n1736 gnd.n1735 0.152939
R13002 gnd.n1737 gnd.n1736 0.152939
R13003 gnd.n1738 gnd.n1737 0.152939
R13004 gnd.n1739 gnd.n1738 0.152939
R13005 gnd.n1740 gnd.n1739 0.152939
R13006 gnd.n1740 gnd.n1051 0.152939
R13007 gnd.n1819 gnd.n1051 0.152939
R13008 gnd.n1820 gnd.n1819 0.152939
R13009 gnd.n1821 gnd.n1820 0.152939
R13010 gnd.n1822 gnd.n1821 0.152939
R13011 gnd.n1823 gnd.n1822 0.152939
R13012 gnd.n1824 gnd.n1823 0.152939
R13013 gnd.n1825 gnd.n1824 0.152939
R13014 gnd.n1826 gnd.n1825 0.152939
R13015 gnd.n1827 gnd.n1826 0.152939
R13016 gnd.n1827 gnd.n997 0.152939
R13017 gnd.n1906 gnd.n997 0.152939
R13018 gnd.n1907 gnd.n1906 0.152939
R13019 gnd.n1908 gnd.n1907 0.152939
R13020 gnd.n1909 gnd.n1908 0.152939
R13021 gnd.n1910 gnd.n1909 0.152939
R13022 gnd.n1911 gnd.n1910 0.152939
R13023 gnd.n1912 gnd.n1911 0.152939
R13024 gnd.n1913 gnd.n1912 0.152939
R13025 gnd.n1914 gnd.n1913 0.152939
R13026 gnd.n1916 gnd.n1914 0.152939
R13027 gnd.n1916 gnd.n1915 0.152939
R13028 gnd.n1490 gnd.n1489 0.152939
R13029 gnd.n1490 gnd.n1380 0.152939
R13030 gnd.n1505 gnd.n1380 0.152939
R13031 gnd.n1506 gnd.n1505 0.152939
R13032 gnd.n1507 gnd.n1506 0.152939
R13033 gnd.n1507 gnd.n1368 0.152939
R13034 gnd.n1521 gnd.n1368 0.152939
R13035 gnd.n1522 gnd.n1521 0.152939
R13036 gnd.n1523 gnd.n1522 0.152939
R13037 gnd.n1524 gnd.n1523 0.152939
R13038 gnd.n1525 gnd.n1524 0.152939
R13039 gnd.n1526 gnd.n1525 0.152939
R13040 gnd.n1527 gnd.n1526 0.152939
R13041 gnd.n1528 gnd.n1527 0.152939
R13042 gnd.n1529 gnd.n1528 0.152939
R13043 gnd.n1530 gnd.n1529 0.152939
R13044 gnd.n1531 gnd.n1530 0.152939
R13045 gnd.n1532 gnd.n1531 0.152939
R13046 gnd.n1533 gnd.n1532 0.152939
R13047 gnd.n1534 gnd.n1533 0.152939
R13048 gnd.n1535 gnd.n1534 0.152939
R13049 gnd.n1535 gnd.n1234 0.152939
R13050 gnd.n1652 gnd.n1234 0.152939
R13051 gnd.n1653 gnd.n1652 0.152939
R13052 gnd.n1654 gnd.n1653 0.152939
R13053 gnd.n1655 gnd.n1654 0.152939
R13054 gnd.n1655 gnd.n1156 0.152939
R13055 gnd.n1732 gnd.n1156 0.152939
R13056 gnd.n1408 gnd.n1407 0.152939
R13057 gnd.n1409 gnd.n1408 0.152939
R13058 gnd.n1410 gnd.n1409 0.152939
R13059 gnd.n1411 gnd.n1410 0.152939
R13060 gnd.n1412 gnd.n1411 0.152939
R13061 gnd.n1413 gnd.n1412 0.152939
R13062 gnd.n1414 gnd.n1413 0.152939
R13063 gnd.n1415 gnd.n1414 0.152939
R13064 gnd.n1416 gnd.n1415 0.152939
R13065 gnd.n1417 gnd.n1416 0.152939
R13066 gnd.n1418 gnd.n1417 0.152939
R13067 gnd.n1419 gnd.n1418 0.152939
R13068 gnd.n1420 gnd.n1419 0.152939
R13069 gnd.n1421 gnd.n1420 0.152939
R13070 gnd.n1422 gnd.n1421 0.152939
R13071 gnd.n1423 gnd.n1422 0.152939
R13072 gnd.n1424 gnd.n1423 0.152939
R13073 gnd.n1425 gnd.n1424 0.152939
R13074 gnd.n1426 gnd.n1425 0.152939
R13075 gnd.n1427 gnd.n1426 0.152939
R13076 gnd.n1428 gnd.n1427 0.152939
R13077 gnd.n1429 gnd.n1428 0.152939
R13078 gnd.n1433 gnd.n1429 0.152939
R13079 gnd.n1434 gnd.n1433 0.152939
R13080 gnd.n1434 gnd.n1391 0.152939
R13081 gnd.n1488 gnd.n1391 0.152939
R13082 gnd.n6497 gnd.n702 0.152939
R13083 gnd.n6505 gnd.n702 0.152939
R13084 gnd.n6506 gnd.n6505 0.152939
R13085 gnd.n6507 gnd.n6506 0.152939
R13086 gnd.n6507 gnd.n696 0.152939
R13087 gnd.n6515 gnd.n696 0.152939
R13088 gnd.n6516 gnd.n6515 0.152939
R13089 gnd.n6517 gnd.n6516 0.152939
R13090 gnd.n6517 gnd.n690 0.152939
R13091 gnd.n6525 gnd.n690 0.152939
R13092 gnd.n6526 gnd.n6525 0.152939
R13093 gnd.n6527 gnd.n6526 0.152939
R13094 gnd.n6527 gnd.n684 0.152939
R13095 gnd.n6535 gnd.n684 0.152939
R13096 gnd.n6536 gnd.n6535 0.152939
R13097 gnd.n6537 gnd.n6536 0.152939
R13098 gnd.n6537 gnd.n678 0.152939
R13099 gnd.n6545 gnd.n678 0.152939
R13100 gnd.n6546 gnd.n6545 0.152939
R13101 gnd.n6547 gnd.n6546 0.152939
R13102 gnd.n6547 gnd.n672 0.152939
R13103 gnd.n6555 gnd.n672 0.152939
R13104 gnd.n6556 gnd.n6555 0.152939
R13105 gnd.n6557 gnd.n6556 0.152939
R13106 gnd.n6557 gnd.n666 0.152939
R13107 gnd.n6565 gnd.n666 0.152939
R13108 gnd.n6566 gnd.n6565 0.152939
R13109 gnd.n6567 gnd.n6566 0.152939
R13110 gnd.n6567 gnd.n660 0.152939
R13111 gnd.n6575 gnd.n660 0.152939
R13112 gnd.n6576 gnd.n6575 0.152939
R13113 gnd.n6577 gnd.n6576 0.152939
R13114 gnd.n6577 gnd.n654 0.152939
R13115 gnd.n6585 gnd.n654 0.152939
R13116 gnd.n6586 gnd.n6585 0.152939
R13117 gnd.n6587 gnd.n6586 0.152939
R13118 gnd.n6587 gnd.n648 0.152939
R13119 gnd.n6595 gnd.n648 0.152939
R13120 gnd.n6596 gnd.n6595 0.152939
R13121 gnd.n6597 gnd.n6596 0.152939
R13122 gnd.n6597 gnd.n642 0.152939
R13123 gnd.n6605 gnd.n642 0.152939
R13124 gnd.n6606 gnd.n6605 0.152939
R13125 gnd.n6607 gnd.n6606 0.152939
R13126 gnd.n6607 gnd.n636 0.152939
R13127 gnd.n6615 gnd.n636 0.152939
R13128 gnd.n6616 gnd.n6615 0.152939
R13129 gnd.n6617 gnd.n6616 0.152939
R13130 gnd.n6617 gnd.n630 0.152939
R13131 gnd.n6625 gnd.n630 0.152939
R13132 gnd.n6626 gnd.n6625 0.152939
R13133 gnd.n6627 gnd.n6626 0.152939
R13134 gnd.n6627 gnd.n624 0.152939
R13135 gnd.n6635 gnd.n624 0.152939
R13136 gnd.n6636 gnd.n6635 0.152939
R13137 gnd.n6637 gnd.n6636 0.152939
R13138 gnd.n6637 gnd.n618 0.152939
R13139 gnd.n6645 gnd.n618 0.152939
R13140 gnd.n6646 gnd.n6645 0.152939
R13141 gnd.n6647 gnd.n6646 0.152939
R13142 gnd.n6647 gnd.n612 0.152939
R13143 gnd.n6655 gnd.n612 0.152939
R13144 gnd.n6656 gnd.n6655 0.152939
R13145 gnd.n6657 gnd.n6656 0.152939
R13146 gnd.n6657 gnd.n606 0.152939
R13147 gnd.n6665 gnd.n606 0.152939
R13148 gnd.n6666 gnd.n6665 0.152939
R13149 gnd.n6667 gnd.n6666 0.152939
R13150 gnd.n6667 gnd.n600 0.152939
R13151 gnd.n6675 gnd.n600 0.152939
R13152 gnd.n6676 gnd.n6675 0.152939
R13153 gnd.n6677 gnd.n6676 0.152939
R13154 gnd.n6677 gnd.n594 0.152939
R13155 gnd.n6685 gnd.n594 0.152939
R13156 gnd.n6686 gnd.n6685 0.152939
R13157 gnd.n6687 gnd.n6686 0.152939
R13158 gnd.n6687 gnd.n588 0.152939
R13159 gnd.n6695 gnd.n588 0.152939
R13160 gnd.n6696 gnd.n6695 0.152939
R13161 gnd.n6697 gnd.n6696 0.152939
R13162 gnd.n6697 gnd.n582 0.152939
R13163 gnd.n6705 gnd.n582 0.152939
R13164 gnd.n6706 gnd.n6705 0.152939
R13165 gnd.n6707 gnd.n6706 0.152939
R13166 gnd.n6707 gnd.n576 0.152939
R13167 gnd.n6715 gnd.n576 0.152939
R13168 gnd.n6716 gnd.n6715 0.152939
R13169 gnd.n6717 gnd.n6716 0.152939
R13170 gnd.n6717 gnd.n570 0.152939
R13171 gnd.n6725 gnd.n570 0.152939
R13172 gnd.n6726 gnd.n6725 0.152939
R13173 gnd.n6727 gnd.n6726 0.152939
R13174 gnd.n6727 gnd.n564 0.152939
R13175 gnd.n6735 gnd.n564 0.152939
R13176 gnd.n6736 gnd.n6735 0.152939
R13177 gnd.n6737 gnd.n6736 0.152939
R13178 gnd.n6737 gnd.n558 0.152939
R13179 gnd.n6745 gnd.n558 0.152939
R13180 gnd.n6746 gnd.n6745 0.152939
R13181 gnd.n6747 gnd.n6746 0.152939
R13182 gnd.n6747 gnd.n552 0.152939
R13183 gnd.n6755 gnd.n552 0.152939
R13184 gnd.n6756 gnd.n6755 0.152939
R13185 gnd.n6757 gnd.n6756 0.152939
R13186 gnd.n6757 gnd.n546 0.152939
R13187 gnd.n6765 gnd.n546 0.152939
R13188 gnd.n6766 gnd.n6765 0.152939
R13189 gnd.n6767 gnd.n6766 0.152939
R13190 gnd.n6767 gnd.n540 0.152939
R13191 gnd.n6775 gnd.n540 0.152939
R13192 gnd.n6776 gnd.n6775 0.152939
R13193 gnd.n6777 gnd.n6776 0.152939
R13194 gnd.n6777 gnd.n534 0.152939
R13195 gnd.n6785 gnd.n534 0.152939
R13196 gnd.n6786 gnd.n6785 0.152939
R13197 gnd.n6787 gnd.n6786 0.152939
R13198 gnd.n6787 gnd.n528 0.152939
R13199 gnd.n6795 gnd.n528 0.152939
R13200 gnd.n6796 gnd.n6795 0.152939
R13201 gnd.n6797 gnd.n6796 0.152939
R13202 gnd.n6797 gnd.n522 0.152939
R13203 gnd.n6805 gnd.n522 0.152939
R13204 gnd.n6806 gnd.n6805 0.152939
R13205 gnd.n6807 gnd.n6806 0.152939
R13206 gnd.n6807 gnd.n516 0.152939
R13207 gnd.n6815 gnd.n516 0.152939
R13208 gnd.n6816 gnd.n6815 0.152939
R13209 gnd.n6817 gnd.n6816 0.152939
R13210 gnd.n6817 gnd.n510 0.152939
R13211 gnd.n6825 gnd.n510 0.152939
R13212 gnd.n6826 gnd.n6825 0.152939
R13213 gnd.n6827 gnd.n6826 0.152939
R13214 gnd.n6827 gnd.n504 0.152939
R13215 gnd.n6835 gnd.n504 0.152939
R13216 gnd.n6836 gnd.n6835 0.152939
R13217 gnd.n6837 gnd.n6836 0.152939
R13218 gnd.n6837 gnd.n498 0.152939
R13219 gnd.n6845 gnd.n498 0.152939
R13220 gnd.n6846 gnd.n6845 0.152939
R13221 gnd.n6847 gnd.n6846 0.152939
R13222 gnd.n6847 gnd.n492 0.152939
R13223 gnd.n6855 gnd.n492 0.152939
R13224 gnd.n6856 gnd.n6855 0.152939
R13225 gnd.n6857 gnd.n6856 0.152939
R13226 gnd.n6857 gnd.n486 0.152939
R13227 gnd.n6865 gnd.n486 0.152939
R13228 gnd.n6866 gnd.n6865 0.152939
R13229 gnd.n6867 gnd.n6866 0.152939
R13230 gnd.n6867 gnd.n480 0.152939
R13231 gnd.n6875 gnd.n480 0.152939
R13232 gnd.n6876 gnd.n6875 0.152939
R13233 gnd.n6877 gnd.n6876 0.152939
R13234 gnd.n6877 gnd.n474 0.152939
R13235 gnd.n6885 gnd.n474 0.152939
R13236 gnd.n6886 gnd.n6885 0.152939
R13237 gnd.n6887 gnd.n6886 0.152939
R13238 gnd.n6887 gnd.n468 0.152939
R13239 gnd.n6895 gnd.n468 0.152939
R13240 gnd.n6896 gnd.n6895 0.152939
R13241 gnd.n6897 gnd.n6896 0.152939
R13242 gnd.n6897 gnd.n462 0.152939
R13243 gnd.n6905 gnd.n462 0.152939
R13244 gnd.n6906 gnd.n6905 0.152939
R13245 gnd.n6907 gnd.n6906 0.152939
R13246 gnd.n6907 gnd.n456 0.152939
R13247 gnd.n6915 gnd.n456 0.152939
R13248 gnd.n6916 gnd.n6915 0.152939
R13249 gnd.n6917 gnd.n6916 0.152939
R13250 gnd.n6917 gnd.n450 0.152939
R13251 gnd.n6925 gnd.n450 0.152939
R13252 gnd.n6926 gnd.n6925 0.152939
R13253 gnd.n6927 gnd.n6926 0.152939
R13254 gnd.n6927 gnd.n444 0.152939
R13255 gnd.n6935 gnd.n444 0.152939
R13256 gnd.n6936 gnd.n6935 0.152939
R13257 gnd.n6937 gnd.n6936 0.152939
R13258 gnd.n6937 gnd.n438 0.152939
R13259 gnd.n6945 gnd.n438 0.152939
R13260 gnd.n6946 gnd.n6945 0.152939
R13261 gnd.n6947 gnd.n6946 0.152939
R13262 gnd.n6947 gnd.n432 0.152939
R13263 gnd.n6955 gnd.n432 0.152939
R13264 gnd.n6956 gnd.n6955 0.152939
R13265 gnd.n6957 gnd.n6956 0.152939
R13266 gnd.n6957 gnd.n426 0.152939
R13267 gnd.n6965 gnd.n426 0.152939
R13268 gnd.n6966 gnd.n6965 0.152939
R13269 gnd.n6967 gnd.n6966 0.152939
R13270 gnd.n6967 gnd.n420 0.152939
R13271 gnd.n6975 gnd.n420 0.152939
R13272 gnd.n6976 gnd.n6975 0.152939
R13273 gnd.n6977 gnd.n6976 0.152939
R13274 gnd.n6977 gnd.n414 0.152939
R13275 gnd.n6985 gnd.n414 0.152939
R13276 gnd.n6986 gnd.n6985 0.152939
R13277 gnd.n6987 gnd.n6986 0.152939
R13278 gnd.n6987 gnd.n408 0.152939
R13279 gnd.n6995 gnd.n408 0.152939
R13280 gnd.n6996 gnd.n6995 0.152939
R13281 gnd.n6997 gnd.n6996 0.152939
R13282 gnd.n6997 gnd.n402 0.152939
R13283 gnd.n7005 gnd.n402 0.152939
R13284 gnd.n7006 gnd.n7005 0.152939
R13285 gnd.n7008 gnd.n7006 0.152939
R13286 gnd.n7008 gnd.n7007 0.152939
R13287 gnd.n7007 gnd.n396 0.152939
R13288 gnd.n7017 gnd.n396 0.152939
R13289 gnd.n7018 gnd.n391 0.152939
R13290 gnd.n7026 gnd.n391 0.152939
R13291 gnd.n7027 gnd.n7026 0.152939
R13292 gnd.n7028 gnd.n7027 0.152939
R13293 gnd.n7028 gnd.n385 0.152939
R13294 gnd.n7036 gnd.n385 0.152939
R13295 gnd.n7037 gnd.n7036 0.152939
R13296 gnd.n7038 gnd.n7037 0.152939
R13297 gnd.n7038 gnd.n379 0.152939
R13298 gnd.n7046 gnd.n379 0.152939
R13299 gnd.n7047 gnd.n7046 0.152939
R13300 gnd.n7048 gnd.n7047 0.152939
R13301 gnd.n7048 gnd.n373 0.152939
R13302 gnd.n7056 gnd.n373 0.152939
R13303 gnd.n7057 gnd.n7056 0.152939
R13304 gnd.n7058 gnd.n7057 0.152939
R13305 gnd.n7058 gnd.n367 0.152939
R13306 gnd.n7066 gnd.n367 0.152939
R13307 gnd.n7067 gnd.n7066 0.152939
R13308 gnd.n7068 gnd.n7067 0.152939
R13309 gnd.n7068 gnd.n361 0.152939
R13310 gnd.n7076 gnd.n361 0.152939
R13311 gnd.n7077 gnd.n7076 0.152939
R13312 gnd.n7078 gnd.n7077 0.152939
R13313 gnd.n7078 gnd.n355 0.152939
R13314 gnd.n7086 gnd.n355 0.152939
R13315 gnd.n7087 gnd.n7086 0.152939
R13316 gnd.n7088 gnd.n7087 0.152939
R13317 gnd.n7088 gnd.n349 0.152939
R13318 gnd.n7096 gnd.n349 0.152939
R13319 gnd.n7097 gnd.n7096 0.152939
R13320 gnd.n7098 gnd.n7097 0.152939
R13321 gnd.n7098 gnd.n343 0.152939
R13322 gnd.n7106 gnd.n343 0.152939
R13323 gnd.n7107 gnd.n7106 0.152939
R13324 gnd.n7108 gnd.n7107 0.152939
R13325 gnd.n7108 gnd.n337 0.152939
R13326 gnd.n7116 gnd.n337 0.152939
R13327 gnd.n7117 gnd.n7116 0.152939
R13328 gnd.n7118 gnd.n7117 0.152939
R13329 gnd.n7118 gnd.n331 0.152939
R13330 gnd.n7126 gnd.n331 0.152939
R13331 gnd.n7127 gnd.n7126 0.152939
R13332 gnd.n7128 gnd.n7127 0.152939
R13333 gnd.n7128 gnd.n325 0.152939
R13334 gnd.n7136 gnd.n325 0.152939
R13335 gnd.n7137 gnd.n7136 0.152939
R13336 gnd.n7138 gnd.n7137 0.152939
R13337 gnd.n7138 gnd.n319 0.152939
R13338 gnd.n7146 gnd.n319 0.152939
R13339 gnd.n7147 gnd.n7146 0.152939
R13340 gnd.n7148 gnd.n7147 0.152939
R13341 gnd.n7148 gnd.n313 0.152939
R13342 gnd.n7156 gnd.n313 0.152939
R13343 gnd.n7157 gnd.n7156 0.152939
R13344 gnd.n7158 gnd.n7157 0.152939
R13345 gnd.n7158 gnd.n307 0.152939
R13346 gnd.n7166 gnd.n307 0.152939
R13347 gnd.n7167 gnd.n7166 0.152939
R13348 gnd.n7168 gnd.n7167 0.152939
R13349 gnd.n7168 gnd.n301 0.152939
R13350 gnd.n7176 gnd.n301 0.152939
R13351 gnd.n7177 gnd.n7176 0.152939
R13352 gnd.n7178 gnd.n7177 0.152939
R13353 gnd.n7178 gnd.n295 0.152939
R13354 gnd.n7186 gnd.n295 0.152939
R13355 gnd.n7187 gnd.n7186 0.152939
R13356 gnd.n7188 gnd.n7187 0.152939
R13357 gnd.n7188 gnd.n289 0.152939
R13358 gnd.n7196 gnd.n289 0.152939
R13359 gnd.n7197 gnd.n7196 0.152939
R13360 gnd.n7198 gnd.n7197 0.152939
R13361 gnd.n7198 gnd.n283 0.152939
R13362 gnd.n7206 gnd.n283 0.152939
R13363 gnd.n7207 gnd.n7206 0.152939
R13364 gnd.n7208 gnd.n7207 0.152939
R13365 gnd.n7208 gnd.n277 0.152939
R13366 gnd.n7216 gnd.n277 0.152939
R13367 gnd.n7217 gnd.n7216 0.152939
R13368 gnd.n7218 gnd.n7217 0.152939
R13369 gnd.n7218 gnd.n271 0.152939
R13370 gnd.n7226 gnd.n271 0.152939
R13371 gnd.n7227 gnd.n7226 0.152939
R13372 gnd.n7229 gnd.n7227 0.152939
R13373 gnd.n3150 gnd.n3147 0.152939
R13374 gnd.n3151 gnd.n3150 0.152939
R13375 gnd.n3152 gnd.n3151 0.152939
R13376 gnd.n3153 gnd.n3152 0.152939
R13377 gnd.n3156 gnd.n3153 0.152939
R13378 gnd.n3157 gnd.n3156 0.152939
R13379 gnd.n3158 gnd.n3157 0.152939
R13380 gnd.n3159 gnd.n3158 0.152939
R13381 gnd.n3162 gnd.n3159 0.152939
R13382 gnd.n3163 gnd.n3162 0.152939
R13383 gnd.n3164 gnd.n3163 0.152939
R13384 gnd.n3165 gnd.n3164 0.152939
R13385 gnd.n3168 gnd.n3165 0.152939
R13386 gnd.n3169 gnd.n3168 0.152939
R13387 gnd.n3170 gnd.n3169 0.152939
R13388 gnd.n3172 gnd.n3170 0.152939
R13389 gnd.n3172 gnd.n3171 0.152939
R13390 gnd.n3171 gnd.n247 0.152939
R13391 gnd.n248 gnd.n247 0.152939
R13392 gnd.n249 gnd.n248 0.152939
R13393 gnd.n254 gnd.n249 0.152939
R13394 gnd.n255 gnd.n254 0.152939
R13395 gnd.n256 gnd.n255 0.152939
R13396 gnd.n257 gnd.n256 0.152939
R13397 gnd.n262 gnd.n257 0.152939
R13398 gnd.n263 gnd.n262 0.152939
R13399 gnd.n264 gnd.n263 0.152939
R13400 gnd.n265 gnd.n264 0.152939
R13401 gnd.n7228 gnd.n265 0.152939
R13402 gnd.n7536 gnd.n77 0.152939
R13403 gnd.n103 gnd.n77 0.152939
R13404 gnd.n104 gnd.n103 0.152939
R13405 gnd.n105 gnd.n104 0.152939
R13406 gnd.n122 gnd.n105 0.152939
R13407 gnd.n123 gnd.n122 0.152939
R13408 gnd.n124 gnd.n123 0.152939
R13409 gnd.n125 gnd.n124 0.152939
R13410 gnd.n143 gnd.n125 0.152939
R13411 gnd.n144 gnd.n143 0.152939
R13412 gnd.n145 gnd.n144 0.152939
R13413 gnd.n146 gnd.n145 0.152939
R13414 gnd.n163 gnd.n146 0.152939
R13415 gnd.n164 gnd.n163 0.152939
R13416 gnd.n165 gnd.n164 0.152939
R13417 gnd.n166 gnd.n165 0.152939
R13418 gnd.n7545 gnd.n65 0.152939
R13419 gnd.n5693 gnd.n65 0.152939
R13420 gnd.n5694 gnd.n5693 0.152939
R13421 gnd.n5694 gnd.n3200 0.152939
R13422 gnd.n5706 gnd.n3200 0.152939
R13423 gnd.n5707 gnd.n5706 0.152939
R13424 gnd.n5709 gnd.n5707 0.152939
R13425 gnd.n5709 gnd.n5708 0.152939
R13426 gnd.n5708 gnd.n3193 0.152939
R13427 gnd.n3194 gnd.n3193 0.152939
R13428 gnd.n3195 gnd.n3194 0.152939
R13429 gnd.n5720 gnd.n3195 0.152939
R13430 gnd.n5721 gnd.n5720 0.152939
R13431 gnd.n5722 gnd.n5721 0.152939
R13432 gnd.n5723 gnd.n5722 0.152939
R13433 gnd.n5726 gnd.n5723 0.152939
R13434 gnd.n5728 gnd.n5726 0.152939
R13435 gnd.n5728 gnd.n5727 0.152939
R13436 gnd.n5727 gnd.n178 0.152939
R13437 gnd.n7474 gnd.n178 0.152939
R13438 gnd.n201 gnd.n200 0.152939
R13439 gnd.n208 gnd.n200 0.152939
R13440 gnd.n209 gnd.n208 0.152939
R13441 gnd.n210 gnd.n209 0.152939
R13442 gnd.n210 gnd.n198 0.152939
R13443 gnd.n218 gnd.n198 0.152939
R13444 gnd.n219 gnd.n218 0.152939
R13445 gnd.n220 gnd.n219 0.152939
R13446 gnd.n220 gnd.n196 0.152939
R13447 gnd.n228 gnd.n196 0.152939
R13448 gnd.n229 gnd.n228 0.152939
R13449 gnd.n230 gnd.n229 0.152939
R13450 gnd.n230 gnd.n194 0.152939
R13451 gnd.n237 gnd.n194 0.152939
R13452 gnd.n238 gnd.n237 0.152939
R13453 gnd.n239 gnd.n238 0.152939
R13454 gnd.n239 gnd.n179 0.152939
R13455 gnd.n7473 gnd.n179 0.152939
R13456 gnd.n7290 gnd.n7289 0.152939
R13457 gnd.n7291 gnd.n7290 0.152939
R13458 gnd.n7292 gnd.n7291 0.152939
R13459 gnd.n7293 gnd.n7292 0.152939
R13460 gnd.n7294 gnd.n7293 0.152939
R13461 gnd.n7295 gnd.n7294 0.152939
R13462 gnd.n7296 gnd.n7295 0.152939
R13463 gnd.n7297 gnd.n7296 0.152939
R13464 gnd.n7298 gnd.n7297 0.152939
R13465 gnd.n7299 gnd.n7298 0.152939
R13466 gnd.n7300 gnd.n7299 0.152939
R13467 gnd.n7301 gnd.n7300 0.152939
R13468 gnd.n7302 gnd.n7301 0.152939
R13469 gnd.n7303 gnd.n7302 0.152939
R13470 gnd.n7304 gnd.n7303 0.152939
R13471 gnd.n7305 gnd.n7304 0.152939
R13472 gnd.n7306 gnd.n7305 0.152939
R13473 gnd.n7307 gnd.n7306 0.152939
R13474 gnd.n7308 gnd.n7307 0.152939
R13475 gnd.n7309 gnd.n7308 0.152939
R13476 gnd.n7310 gnd.n7309 0.152939
R13477 gnd.n7311 gnd.n7310 0.152939
R13478 gnd.n7312 gnd.n7311 0.152939
R13479 gnd.n7313 gnd.n7312 0.152939
R13480 gnd.n7314 gnd.n7313 0.152939
R13481 gnd.n7315 gnd.n7314 0.152939
R13482 gnd.n7316 gnd.n7315 0.152939
R13483 gnd.n7317 gnd.n7316 0.152939
R13484 gnd.n7318 gnd.n7317 0.152939
R13485 gnd.n7319 gnd.n7318 0.152939
R13486 gnd.n7320 gnd.n7319 0.152939
R13487 gnd.n7321 gnd.n7320 0.152939
R13488 gnd.n7322 gnd.n7321 0.152939
R13489 gnd.n7323 gnd.n7322 0.152939
R13490 gnd.n7324 gnd.n7323 0.152939
R13491 gnd.n7325 gnd.n7324 0.152939
R13492 gnd.n7393 gnd.n7325 0.152939
R13493 gnd.n7393 gnd.n7392 0.152939
R13494 gnd.n7392 gnd.n7391 0.152939
R13495 gnd.n7391 gnd.n7329 0.152939
R13496 gnd.n7330 gnd.n7329 0.152939
R13497 gnd.n7331 gnd.n7330 0.152939
R13498 gnd.n7332 gnd.n7331 0.152939
R13499 gnd.n7333 gnd.n7332 0.152939
R13500 gnd.n7334 gnd.n7333 0.152939
R13501 gnd.n7335 gnd.n7334 0.152939
R13502 gnd.n7336 gnd.n7335 0.152939
R13503 gnd.n7337 gnd.n7336 0.152939
R13504 gnd.n7338 gnd.n7337 0.152939
R13505 gnd.n7339 gnd.n7338 0.152939
R13506 gnd.n7340 gnd.n7339 0.152939
R13507 gnd.n7341 gnd.n7340 0.152939
R13508 gnd.n7342 gnd.n7341 0.152939
R13509 gnd.n7343 gnd.n7342 0.152939
R13510 gnd.n7344 gnd.n7343 0.152939
R13511 gnd.n7345 gnd.n7344 0.152939
R13512 gnd.n7351 gnd.n7345 0.152939
R13513 gnd.n7351 gnd.n7350 0.152939
R13514 gnd.n5415 gnd.n5414 0.152939
R13515 gnd.n5415 gnd.n5411 0.152939
R13516 gnd.n5423 gnd.n5411 0.152939
R13517 gnd.n5424 gnd.n5423 0.152939
R13518 gnd.n5425 gnd.n5424 0.152939
R13519 gnd.n5425 gnd.n5407 0.152939
R13520 gnd.n5433 gnd.n5407 0.152939
R13521 gnd.n5434 gnd.n5433 0.152939
R13522 gnd.n5435 gnd.n5434 0.152939
R13523 gnd.n5435 gnd.n5403 0.152939
R13524 gnd.n5443 gnd.n5403 0.152939
R13525 gnd.n5444 gnd.n5443 0.152939
R13526 gnd.n5445 gnd.n5444 0.152939
R13527 gnd.n5445 gnd.n5399 0.152939
R13528 gnd.n5453 gnd.n5399 0.152939
R13529 gnd.n5454 gnd.n5453 0.152939
R13530 gnd.n5455 gnd.n5454 0.152939
R13531 gnd.n5455 gnd.n5395 0.152939
R13532 gnd.n5466 gnd.n5395 0.152939
R13533 gnd.n5467 gnd.n5466 0.152939
R13534 gnd.n5468 gnd.n5467 0.152939
R13535 gnd.n5468 gnd.n5391 0.152939
R13536 gnd.n5476 gnd.n5391 0.152939
R13537 gnd.n5477 gnd.n5476 0.152939
R13538 gnd.n5479 gnd.n5477 0.152939
R13539 gnd.n5489 gnd.n3261 0.152939
R13540 gnd.n5490 gnd.n5489 0.152939
R13541 gnd.n5491 gnd.n5490 0.152939
R13542 gnd.n5491 gnd.n3257 0.152939
R13543 gnd.n5499 gnd.n3257 0.152939
R13544 gnd.n5500 gnd.n5499 0.152939
R13545 gnd.n5501 gnd.n5500 0.152939
R13546 gnd.n5501 gnd.n3253 0.152939
R13547 gnd.n5511 gnd.n3253 0.152939
R13548 gnd.n5512 gnd.n5511 0.152939
R13549 gnd.n5513 gnd.n5512 0.152939
R13550 gnd.n5513 gnd.n3249 0.152939
R13551 gnd.n5521 gnd.n3249 0.152939
R13552 gnd.n5522 gnd.n5521 0.152939
R13553 gnd.n5523 gnd.n5522 0.152939
R13554 gnd.n5523 gnd.n3245 0.152939
R13555 gnd.n5531 gnd.n3245 0.152939
R13556 gnd.n5532 gnd.n5531 0.152939
R13557 gnd.n5533 gnd.n5532 0.152939
R13558 gnd.n5533 gnd.n3241 0.152939
R13559 gnd.n5541 gnd.n3241 0.152939
R13560 gnd.n5542 gnd.n5541 0.152939
R13561 gnd.n5543 gnd.n5542 0.152939
R13562 gnd.n5543 gnd.n3237 0.152939
R13563 gnd.n5551 gnd.n3237 0.152939
R13564 gnd.n5552 gnd.n5551 0.152939
R13565 gnd.n5554 gnd.n5552 0.152939
R13566 gnd.n5554 gnd.n5553 0.152939
R13567 gnd.n5553 gnd.n3230 0.152939
R13568 gnd.n5563 gnd.n3230 0.152939
R13569 gnd.n3028 gnd.n3027 0.152939
R13570 gnd.n3029 gnd.n3028 0.152939
R13571 gnd.n3049 gnd.n3029 0.152939
R13572 gnd.n3050 gnd.n3049 0.152939
R13573 gnd.n3051 gnd.n3050 0.152939
R13574 gnd.n3052 gnd.n3051 0.152939
R13575 gnd.n3069 gnd.n3052 0.152939
R13576 gnd.n3070 gnd.n3069 0.152939
R13577 gnd.n3071 gnd.n3070 0.152939
R13578 gnd.n3072 gnd.n3071 0.152939
R13579 gnd.n3089 gnd.n3072 0.152939
R13580 gnd.n3090 gnd.n3089 0.152939
R13581 gnd.n3091 gnd.n3090 0.152939
R13582 gnd.n3092 gnd.n3091 0.152939
R13583 gnd.n3092 gnd.n78 0.152939
R13584 gnd.n7536 gnd.n78 0.152939
R13585 gnd.n4277 gnd.n4276 0.152939
R13586 gnd.n4278 gnd.n4277 0.152939
R13587 gnd.n4278 gnd.n3766 0.152939
R13588 gnd.n4335 gnd.n3766 0.152939
R13589 gnd.n4336 gnd.n4335 0.152939
R13590 gnd.n4337 gnd.n4336 0.152939
R13591 gnd.n4337 gnd.n3762 0.152939
R13592 gnd.n4343 gnd.n3762 0.152939
R13593 gnd.n4344 gnd.n4343 0.152939
R13594 gnd.n4345 gnd.n4344 0.152939
R13595 gnd.n4345 gnd.n3758 0.152939
R13596 gnd.n4351 gnd.n3758 0.152939
R13597 gnd.n4352 gnd.n4351 0.152939
R13598 gnd.n4353 gnd.n4352 0.152939
R13599 gnd.n4353 gnd.n3754 0.152939
R13600 gnd.n4359 gnd.n3754 0.152939
R13601 gnd.n4360 gnd.n4359 0.152939
R13602 gnd.n4361 gnd.n4360 0.152939
R13603 gnd.n4361 gnd.n3750 0.152939
R13604 gnd.n4368 gnd.n3750 0.152939
R13605 gnd.n4369 gnd.n4368 0.152939
R13606 gnd.n4370 gnd.n4369 0.152939
R13607 gnd.n4370 gnd.n3745 0.152939
R13608 gnd.n4396 gnd.n3745 0.152939
R13609 gnd.n4397 gnd.n4396 0.152939
R13610 gnd.n4398 gnd.n4397 0.152939
R13611 gnd.n4399 gnd.n4398 0.152939
R13612 gnd.n4399 gnd.n3720 0.152939
R13613 gnd.n4426 gnd.n3720 0.152939
R13614 gnd.n4427 gnd.n4426 0.152939
R13615 gnd.n4428 gnd.n4427 0.152939
R13616 gnd.n4429 gnd.n4428 0.152939
R13617 gnd.n4429 gnd.n3695 0.152939
R13618 gnd.n4456 gnd.n3695 0.152939
R13619 gnd.n4457 gnd.n4456 0.152939
R13620 gnd.n4458 gnd.n4457 0.152939
R13621 gnd.n4459 gnd.n4458 0.152939
R13622 gnd.n4460 gnd.n4459 0.152939
R13623 gnd.n4462 gnd.n4460 0.152939
R13624 gnd.n4463 gnd.n4462 0.152939
R13625 gnd.n4463 gnd.n3601 0.152939
R13626 gnd.n4531 gnd.n3601 0.152939
R13627 gnd.n4532 gnd.n4531 0.152939
R13628 gnd.n4533 gnd.n4532 0.152939
R13629 gnd.n4534 gnd.n4533 0.152939
R13630 gnd.n4534 gnd.n3575 0.152939
R13631 gnd.n4593 gnd.n3575 0.152939
R13632 gnd.n4594 gnd.n4593 0.152939
R13633 gnd.n4595 gnd.n4594 0.152939
R13634 gnd.n4595 gnd.n3557 0.152939
R13635 gnd.n4620 gnd.n3557 0.152939
R13636 gnd.n4621 gnd.n4620 0.152939
R13637 gnd.n4622 gnd.n4621 0.152939
R13638 gnd.n4623 gnd.n4622 0.152939
R13639 gnd.n4623 gnd.n3524 0.152939
R13640 gnd.n4671 gnd.n3524 0.152939
R13641 gnd.n4672 gnd.n4671 0.152939
R13642 gnd.n4673 gnd.n4672 0.152939
R13643 gnd.n4673 gnd.n3501 0.152939
R13644 gnd.n4711 gnd.n3501 0.152939
R13645 gnd.n4712 gnd.n4711 0.152939
R13646 gnd.n4713 gnd.n4712 0.152939
R13647 gnd.n4713 gnd.n3479 0.152939
R13648 gnd.n4767 gnd.n3479 0.152939
R13649 gnd.n4768 gnd.n4767 0.152939
R13650 gnd.n4769 gnd.n4768 0.152939
R13651 gnd.n4769 gnd.n3460 0.152939
R13652 gnd.n4792 gnd.n3460 0.152939
R13653 gnd.n4793 gnd.n4792 0.152939
R13654 gnd.n4794 gnd.n4793 0.152939
R13655 gnd.n4794 gnd.n3440 0.152939
R13656 gnd.n4852 gnd.n3440 0.152939
R13657 gnd.n4853 gnd.n4852 0.152939
R13658 gnd.n4854 gnd.n4853 0.152939
R13659 gnd.n4854 gnd.n3418 0.152939
R13660 gnd.n4881 gnd.n3418 0.152939
R13661 gnd.n4882 gnd.n4881 0.152939
R13662 gnd.n4883 gnd.n4882 0.152939
R13663 gnd.n4884 gnd.n4883 0.152939
R13664 gnd.n4884 gnd.n3390 0.152939
R13665 gnd.n4926 gnd.n3390 0.152939
R13666 gnd.n4927 gnd.n4926 0.152939
R13667 gnd.n4928 gnd.n4927 0.152939
R13668 gnd.n4929 gnd.n4928 0.152939
R13669 gnd.n4931 gnd.n4929 0.152939
R13670 gnd.n4931 gnd.n4930 0.152939
R13671 gnd.n4930 gnd.n3316 0.152939
R13672 gnd.n3317 gnd.n3316 0.152939
R13673 gnd.n3318 gnd.n3317 0.152939
R13674 gnd.n3325 gnd.n3318 0.152939
R13675 gnd.n3326 gnd.n3325 0.152939
R13676 gnd.n3327 gnd.n3326 0.152939
R13677 gnd.n3328 gnd.n3327 0.152939
R13678 gnd.n3337 gnd.n3328 0.152939
R13679 gnd.n3338 gnd.n3337 0.152939
R13680 gnd.n3339 gnd.n3338 0.152939
R13681 gnd.n3340 gnd.n3339 0.152939
R13682 gnd.n3349 gnd.n3340 0.152939
R13683 gnd.n3350 gnd.n3349 0.152939
R13684 gnd.n3351 gnd.n3350 0.152939
R13685 gnd.n3352 gnd.n3351 0.152939
R13686 gnd.n5175 gnd.n3352 0.152939
R13687 gnd.n5177 gnd.n5175 0.152939
R13688 gnd.n5177 gnd.n5176 0.152939
R13689 gnd.n5176 gnd.n3006 0.152939
R13690 gnd.n3007 gnd.n3006 0.152939
R13691 gnd.n3008 gnd.n3007 0.152939
R13692 gnd.n3014 gnd.n3008 0.152939
R13693 gnd.n3015 gnd.n3014 0.152939
R13694 gnd.n3016 gnd.n3015 0.152939
R13695 gnd.n3017 gnd.n3016 0.152939
R13696 gnd.n5608 gnd.n3017 0.152939
R13697 gnd.n5611 gnd.n5608 0.152939
R13698 gnd.n5612 gnd.n5611 0.152939
R13699 gnd.n5613 gnd.n5612 0.152939
R13700 gnd.n5613 gnd.n5604 0.152939
R13701 gnd.n5619 gnd.n5604 0.152939
R13702 gnd.n5620 gnd.n5619 0.152939
R13703 gnd.n5621 gnd.n5620 0.152939
R13704 gnd.n5621 gnd.n3215 0.152939
R13705 gnd.n5627 gnd.n3215 0.152939
R13706 gnd.n5628 gnd.n5627 0.152939
R13707 gnd.n5629 gnd.n5628 0.152939
R13708 gnd.n5630 gnd.n5629 0.152939
R13709 gnd.n5631 gnd.n5630 0.152939
R13710 gnd.n5633 gnd.n5631 0.152939
R13711 gnd.n5634 gnd.n5633 0.152939
R13712 gnd.n3868 gnd.n3836 0.152939
R13713 gnd.n3837 gnd.n3836 0.152939
R13714 gnd.n3838 gnd.n3837 0.152939
R13715 gnd.n4130 gnd.n3838 0.152939
R13716 gnd.n4131 gnd.n4130 0.152939
R13717 gnd.n4132 gnd.n4131 0.152939
R13718 gnd.n4133 gnd.n4132 0.152939
R13719 gnd.n4138 gnd.n4133 0.152939
R13720 gnd.n4139 gnd.n4138 0.152939
R13721 gnd.n4139 gnd.n3816 0.152939
R13722 gnd.n4200 gnd.n3816 0.152939
R13723 gnd.n4201 gnd.n4200 0.152939
R13724 gnd.n4202 gnd.n4201 0.152939
R13725 gnd.n4202 gnd.n3811 0.152939
R13726 gnd.n4214 gnd.n3811 0.152939
R13727 gnd.n4215 gnd.n4214 0.152939
R13728 gnd.n4217 gnd.n4215 0.152939
R13729 gnd.n4217 gnd.n4216 0.152939
R13730 gnd.n4216 gnd.n3802 0.152939
R13731 gnd.n3803 gnd.n3802 0.152939
R13732 gnd.n3909 gnd.n3841 0.152939
R13733 gnd.n3844 gnd.n3841 0.152939
R13734 gnd.n3845 gnd.n3844 0.152939
R13735 gnd.n3848 gnd.n3845 0.152939
R13736 gnd.n3849 gnd.n3848 0.152939
R13737 gnd.n3850 gnd.n3849 0.152939
R13738 gnd.n3851 gnd.n3850 0.152939
R13739 gnd.n3854 gnd.n3851 0.152939
R13740 gnd.n3855 gnd.n3854 0.152939
R13741 gnd.n3856 gnd.n3855 0.152939
R13742 gnd.n3857 gnd.n3856 0.152939
R13743 gnd.n3860 gnd.n3857 0.152939
R13744 gnd.n3861 gnd.n3860 0.152939
R13745 gnd.n3862 gnd.n3861 0.152939
R13746 gnd.n3863 gnd.n3862 0.152939
R13747 gnd.n3867 gnd.n3863 0.152939
R13748 gnd.n3870 gnd.n3867 0.152939
R13749 gnd.n3870 gnd.n3869 0.152939
R13750 gnd.n2505 gnd.n2454 0.152939
R13751 gnd.n2506 gnd.n2505 0.152939
R13752 gnd.n2507 gnd.n2506 0.152939
R13753 gnd.n2508 gnd.n2507 0.152939
R13754 gnd.n2525 gnd.n2508 0.152939
R13755 gnd.n2526 gnd.n2525 0.152939
R13756 gnd.n2527 gnd.n2526 0.152939
R13757 gnd.n2528 gnd.n2527 0.152939
R13758 gnd.n2545 gnd.n2528 0.152939
R13759 gnd.n2546 gnd.n2545 0.152939
R13760 gnd.n2547 gnd.n2546 0.152939
R13761 gnd.n2548 gnd.n2547 0.152939
R13762 gnd.n2566 gnd.n2548 0.152939
R13763 gnd.n2567 gnd.n2566 0.152939
R13764 gnd.n2568 gnd.n2567 0.152939
R13765 gnd.n2569 gnd.n2568 0.152939
R13766 gnd.n2724 gnd.n2723 0.152939
R13767 gnd.n2725 gnd.n2724 0.152939
R13768 gnd.n2726 gnd.n2725 0.152939
R13769 gnd.n2727 gnd.n2726 0.152939
R13770 gnd.n2728 gnd.n2727 0.152939
R13771 gnd.n2729 gnd.n2728 0.152939
R13772 gnd.n2730 gnd.n2729 0.152939
R13773 gnd.n2731 gnd.n2730 0.152939
R13774 gnd.n2732 gnd.n2731 0.152939
R13775 gnd.n2733 gnd.n2732 0.152939
R13776 gnd.n2734 gnd.n2733 0.152939
R13777 gnd.n2735 gnd.n2734 0.152939
R13778 gnd.n2736 gnd.n2735 0.152939
R13779 gnd.n2737 gnd.n2736 0.152939
R13780 gnd.n2738 gnd.n2737 0.152939
R13781 gnd.n2739 gnd.n2738 0.152939
R13782 gnd.n2740 gnd.n2739 0.152939
R13783 gnd.n2743 gnd.n2740 0.152939
R13784 gnd.n2744 gnd.n2743 0.152939
R13785 gnd.n2745 gnd.n2744 0.152939
R13786 gnd.n2746 gnd.n2745 0.152939
R13787 gnd.n2747 gnd.n2746 0.152939
R13788 gnd.n2748 gnd.n2747 0.152939
R13789 gnd.n2749 gnd.n2748 0.152939
R13790 gnd.n2750 gnd.n2749 0.152939
R13791 gnd.n2848 gnd.n2847 0.152939
R13792 gnd.n2847 gnd.n2753 0.152939
R13793 gnd.n2754 gnd.n2753 0.152939
R13794 gnd.n2755 gnd.n2754 0.152939
R13795 gnd.n2756 gnd.n2755 0.152939
R13796 gnd.n2757 gnd.n2756 0.152939
R13797 gnd.n2758 gnd.n2757 0.152939
R13798 gnd.n2759 gnd.n2758 0.152939
R13799 gnd.n2827 gnd.n2759 0.152939
R13800 gnd.n2827 gnd.n2826 0.152939
R13801 gnd.n2826 gnd.n2825 0.152939
R13802 gnd.n2825 gnd.n2763 0.152939
R13803 gnd.n2764 gnd.n2763 0.152939
R13804 gnd.n2765 gnd.n2764 0.152939
R13805 gnd.n2766 gnd.n2765 0.152939
R13806 gnd.n2767 gnd.n2766 0.152939
R13807 gnd.n2768 gnd.n2767 0.152939
R13808 gnd.n2769 gnd.n2768 0.152939
R13809 gnd.n2770 gnd.n2769 0.152939
R13810 gnd.n2771 gnd.n2770 0.152939
R13811 gnd.n2772 gnd.n2771 0.152939
R13812 gnd.n2773 gnd.n2772 0.152939
R13813 gnd.n2774 gnd.n2773 0.152939
R13814 gnd.n2775 gnd.n2774 0.152939
R13815 gnd.n2776 gnd.n2775 0.152939
R13816 gnd.n2777 gnd.n2776 0.152939
R13817 gnd.n2778 gnd.n2777 0.152939
R13818 gnd.n2779 gnd.n2778 0.152939
R13819 gnd.n2785 gnd.n2779 0.152939
R13820 gnd.n2785 gnd.n2784 0.152939
R13821 gnd.n3977 gnd.n3972 0.152939
R13822 gnd.n3978 gnd.n3977 0.152939
R13823 gnd.n3979 gnd.n3978 0.152939
R13824 gnd.n3979 gnd.n3968 0.152939
R13825 gnd.n3987 gnd.n3968 0.152939
R13826 gnd.n3988 gnd.n3987 0.152939
R13827 gnd.n3989 gnd.n3988 0.152939
R13828 gnd.n3989 gnd.n3964 0.152939
R13829 gnd.n3997 gnd.n3964 0.152939
R13830 gnd.n3998 gnd.n3997 0.152939
R13831 gnd.n3999 gnd.n3998 0.152939
R13832 gnd.n3999 gnd.n3960 0.152939
R13833 gnd.n4007 gnd.n3960 0.152939
R13834 gnd.n4008 gnd.n4007 0.152939
R13835 gnd.n4009 gnd.n4008 0.152939
R13836 gnd.n4009 gnd.n3953 0.152939
R13837 gnd.n4017 gnd.n3953 0.152939
R13838 gnd.n4018 gnd.n4017 0.152939
R13839 gnd.n4019 gnd.n4018 0.152939
R13840 gnd.n4019 gnd.n3949 0.152939
R13841 gnd.n4027 gnd.n3949 0.152939
R13842 gnd.n4028 gnd.n4027 0.152939
R13843 gnd.n4029 gnd.n4028 0.152939
R13844 gnd.n4029 gnd.n3945 0.152939
R13845 gnd.n4037 gnd.n3945 0.152939
R13846 gnd.n4038 gnd.n4037 0.152939
R13847 gnd.n4039 gnd.n4038 0.152939
R13848 gnd.n4039 gnd.n3941 0.152939
R13849 gnd.n4047 gnd.n3941 0.152939
R13850 gnd.n4048 gnd.n4047 0.152939
R13851 gnd.n4049 gnd.n4048 0.152939
R13852 gnd.n4049 gnd.n3937 0.152939
R13853 gnd.n4057 gnd.n3937 0.152939
R13854 gnd.n4058 gnd.n4057 0.152939
R13855 gnd.n4059 gnd.n4058 0.152939
R13856 gnd.n4059 gnd.n3933 0.152939
R13857 gnd.n4069 gnd.n3933 0.152939
R13858 gnd.n4070 gnd.n4069 0.152939
R13859 gnd.n4071 gnd.n4070 0.152939
R13860 gnd.n4071 gnd.n3929 0.152939
R13861 gnd.n4079 gnd.n3929 0.152939
R13862 gnd.n4080 gnd.n4079 0.152939
R13863 gnd.n4081 gnd.n4080 0.152939
R13864 gnd.n4081 gnd.n3925 0.152939
R13865 gnd.n4089 gnd.n3925 0.152939
R13866 gnd.n4090 gnd.n4089 0.152939
R13867 gnd.n4091 gnd.n4090 0.152939
R13868 gnd.n4091 gnd.n3921 0.152939
R13869 gnd.n4099 gnd.n3921 0.152939
R13870 gnd.n4100 gnd.n4099 0.152939
R13871 gnd.n4101 gnd.n4100 0.152939
R13872 gnd.n4101 gnd.n3917 0.152939
R13873 gnd.n4109 gnd.n3917 0.152939
R13874 gnd.n4110 gnd.n4109 0.152939
R13875 gnd.n4112 gnd.n4110 0.152939
R13876 gnd.n4112 gnd.n4111 0.152939
R13877 gnd.n4111 gnd.n3910 0.152939
R13878 gnd.n4121 gnd.n3910 0.152939
R13879 gnd.n2371 gnd.n2370 0.152939
R13880 gnd.n2372 gnd.n2371 0.152939
R13881 gnd.n2391 gnd.n2372 0.152939
R13882 gnd.n2392 gnd.n2391 0.152939
R13883 gnd.n2393 gnd.n2392 0.152939
R13884 gnd.n2394 gnd.n2393 0.152939
R13885 gnd.n2412 gnd.n2394 0.152939
R13886 gnd.n2413 gnd.n2412 0.152939
R13887 gnd.n2414 gnd.n2413 0.152939
R13888 gnd.n2415 gnd.n2414 0.152939
R13889 gnd.n2432 gnd.n2415 0.152939
R13890 gnd.n2433 gnd.n2432 0.152939
R13891 gnd.n2434 gnd.n2433 0.152939
R13892 gnd.n2435 gnd.n2434 0.152939
R13893 gnd.n2453 gnd.n2435 0.152939
R13894 gnd.n2454 gnd.n2453 0.152939
R13895 gnd.n6325 gnd.n874 0.152939
R13896 gnd.n2342 gnd.n874 0.152939
R13897 gnd.n2343 gnd.n2342 0.152939
R13898 gnd.n2344 gnd.n2343 0.152939
R13899 gnd.n2349 gnd.n2344 0.152939
R13900 gnd.n2350 gnd.n2349 0.152939
R13901 gnd.n2351 gnd.n2350 0.152939
R13902 gnd.n2352 gnd.n2351 0.152939
R13903 gnd.n2357 gnd.n2352 0.152939
R13904 gnd.n2358 gnd.n2357 0.152939
R13905 gnd.n2359 gnd.n2358 0.152939
R13906 gnd.n2360 gnd.n2359 0.152939
R13907 gnd.n3830 gnd.n2360 0.152939
R13908 gnd.n3831 gnd.n3830 0.152939
R13909 gnd.n4170 gnd.n3831 0.152939
R13910 gnd.n4171 gnd.n4170 0.152939
R13911 gnd.n4172 gnd.n4171 0.152939
R13912 gnd.n4172 gnd.n3826 0.152939
R13913 gnd.n4178 gnd.n3826 0.152939
R13914 gnd.n4179 gnd.n4178 0.152939
R13915 gnd.n4180 gnd.n4179 0.152939
R13916 gnd.n4180 gnd.n3822 0.152939
R13917 gnd.n4186 gnd.n3822 0.152939
R13918 gnd.n4187 gnd.n4186 0.152939
R13919 gnd.n4188 gnd.n4187 0.152939
R13920 gnd.n4189 gnd.n4188 0.152939
R13921 gnd.n4190 gnd.n4189 0.152939
R13922 gnd.n4190 gnd.n3793 0.152939
R13923 gnd.n4274 gnd.n3793 0.152939
R13924 gnd.n6496 gnd.n707 0.152939
R13925 gnd.n712 gnd.n707 0.152939
R13926 gnd.n713 gnd.n712 0.152939
R13927 gnd.n714 gnd.n713 0.152939
R13928 gnd.n715 gnd.n714 0.152939
R13929 gnd.n720 gnd.n715 0.152939
R13930 gnd.n721 gnd.n720 0.152939
R13931 gnd.n722 gnd.n721 0.152939
R13932 gnd.n723 gnd.n722 0.152939
R13933 gnd.n728 gnd.n723 0.152939
R13934 gnd.n729 gnd.n728 0.152939
R13935 gnd.n730 gnd.n729 0.152939
R13936 gnd.n731 gnd.n730 0.152939
R13937 gnd.n736 gnd.n731 0.152939
R13938 gnd.n737 gnd.n736 0.152939
R13939 gnd.n738 gnd.n737 0.152939
R13940 gnd.n739 gnd.n738 0.152939
R13941 gnd.n744 gnd.n739 0.152939
R13942 gnd.n745 gnd.n744 0.152939
R13943 gnd.n746 gnd.n745 0.152939
R13944 gnd.n747 gnd.n746 0.152939
R13945 gnd.n752 gnd.n747 0.152939
R13946 gnd.n753 gnd.n752 0.152939
R13947 gnd.n754 gnd.n753 0.152939
R13948 gnd.n755 gnd.n754 0.152939
R13949 gnd.n760 gnd.n755 0.152939
R13950 gnd.n761 gnd.n760 0.152939
R13951 gnd.n762 gnd.n761 0.152939
R13952 gnd.n763 gnd.n762 0.152939
R13953 gnd.n768 gnd.n763 0.152939
R13954 gnd.n769 gnd.n768 0.152939
R13955 gnd.n770 gnd.n769 0.152939
R13956 gnd.n771 gnd.n770 0.152939
R13957 gnd.n776 gnd.n771 0.152939
R13958 gnd.n777 gnd.n776 0.152939
R13959 gnd.n778 gnd.n777 0.152939
R13960 gnd.n779 gnd.n778 0.152939
R13961 gnd.n784 gnd.n779 0.152939
R13962 gnd.n785 gnd.n784 0.152939
R13963 gnd.n786 gnd.n785 0.152939
R13964 gnd.n787 gnd.n786 0.152939
R13965 gnd.n792 gnd.n787 0.152939
R13966 gnd.n793 gnd.n792 0.152939
R13967 gnd.n794 gnd.n793 0.152939
R13968 gnd.n795 gnd.n794 0.152939
R13969 gnd.n800 gnd.n795 0.152939
R13970 gnd.n801 gnd.n800 0.152939
R13971 gnd.n802 gnd.n801 0.152939
R13972 gnd.n803 gnd.n802 0.152939
R13973 gnd.n808 gnd.n803 0.152939
R13974 gnd.n809 gnd.n808 0.152939
R13975 gnd.n810 gnd.n809 0.152939
R13976 gnd.n811 gnd.n810 0.152939
R13977 gnd.n816 gnd.n811 0.152939
R13978 gnd.n817 gnd.n816 0.152939
R13979 gnd.n818 gnd.n817 0.152939
R13980 gnd.n819 gnd.n818 0.152939
R13981 gnd.n824 gnd.n819 0.152939
R13982 gnd.n825 gnd.n824 0.152939
R13983 gnd.n826 gnd.n825 0.152939
R13984 gnd.n827 gnd.n826 0.152939
R13985 gnd.n832 gnd.n827 0.152939
R13986 gnd.n833 gnd.n832 0.152939
R13987 gnd.n834 gnd.n833 0.152939
R13988 gnd.n835 gnd.n834 0.152939
R13989 gnd.n840 gnd.n835 0.152939
R13990 gnd.n841 gnd.n840 0.152939
R13991 gnd.n842 gnd.n841 0.152939
R13992 gnd.n843 gnd.n842 0.152939
R13993 gnd.n848 gnd.n843 0.152939
R13994 gnd.n849 gnd.n848 0.152939
R13995 gnd.n850 gnd.n849 0.152939
R13996 gnd.n851 gnd.n850 0.152939
R13997 gnd.n856 gnd.n851 0.152939
R13998 gnd.n857 gnd.n856 0.152939
R13999 gnd.n858 gnd.n857 0.152939
R14000 gnd.n859 gnd.n858 0.152939
R14001 gnd.n864 gnd.n859 0.152939
R14002 gnd.n865 gnd.n864 0.152939
R14003 gnd.n866 gnd.n865 0.152939
R14004 gnd.n867 gnd.n866 0.152939
R14005 gnd.n872 gnd.n867 0.152939
R14006 gnd.n873 gnd.n872 0.152939
R14007 gnd.n6326 gnd.n873 0.152939
R14008 gnd.n4387 gnd.n4386 0.152939
R14009 gnd.n4389 gnd.n4387 0.152939
R14010 gnd.n4389 gnd.n4388 0.152939
R14011 gnd.n4388 gnd.n3726 0.152939
R14012 gnd.n4416 gnd.n3726 0.152939
R14013 gnd.n4417 gnd.n4416 0.152939
R14014 gnd.n4419 gnd.n4417 0.152939
R14015 gnd.n4419 gnd.n4418 0.152939
R14016 gnd.n4418 gnd.n3702 0.152939
R14017 gnd.n4446 gnd.n3702 0.152939
R14018 gnd.n4447 gnd.n4446 0.152939
R14019 gnd.n4449 gnd.n4447 0.152939
R14020 gnd.n4449 gnd.n4448 0.152939
R14021 gnd.n4448 gnd.n3677 0.152939
R14022 gnd.n4486 gnd.n3677 0.152939
R14023 gnd.n4487 gnd.n4486 0.152939
R14024 gnd.n4492 gnd.n4487 0.152939
R14025 gnd.n4492 gnd.n4491 0.152939
R14026 gnd.n4491 gnd.n4490 0.152939
R14027 gnd.n4490 gnd.n3593 0.152939
R14028 gnd.n4542 gnd.n3593 0.152939
R14029 gnd.n4543 gnd.n4542 0.152939
R14030 gnd.n4564 gnd.n4543 0.152939
R14031 gnd.n4564 gnd.n4563 0.152939
R14032 gnd.n4563 gnd.n4562 0.152939
R14033 gnd.n4562 gnd.n4544 0.152939
R14034 gnd.n4558 gnd.n4544 0.152939
R14035 gnd.n4558 gnd.n4557 0.152939
R14036 gnd.n4557 gnd.n4556 0.152939
R14037 gnd.n4556 gnd.n4553 0.152939
R14038 gnd.n4553 gnd.n4552 0.152939
R14039 gnd.n4552 gnd.n3541 0.152939
R14040 gnd.n4644 gnd.n3541 0.152939
R14041 gnd.n4645 gnd.n4644 0.152939
R14042 gnd.n4646 gnd.n4645 0.152939
R14043 gnd.n4646 gnd.n3517 0.152939
R14044 gnd.n4694 gnd.n3517 0.152939
R14045 gnd.n4694 gnd.n4693 0.152939
R14046 gnd.n4693 gnd.n4692 0.152939
R14047 gnd.n4692 gnd.n3494 0.152939
R14048 gnd.n4752 gnd.n3494 0.152939
R14049 gnd.n4752 gnd.n4751 0.152939
R14050 gnd.n4751 gnd.n4750 0.152939
R14051 gnd.n4750 gnd.n3495 0.152939
R14052 gnd.n4746 gnd.n3495 0.152939
R14053 gnd.n4746 gnd.n4745 0.152939
R14054 gnd.n4745 gnd.n4744 0.152939
R14055 gnd.n4744 gnd.n4735 0.152939
R14056 gnd.n4740 gnd.n4735 0.152939
R14057 gnd.n4740 gnd.n3433 0.152939
R14058 gnd.n4862 gnd.n3433 0.152939
R14059 gnd.n4863 gnd.n4862 0.152939
R14060 gnd.n4865 gnd.n4863 0.152939
R14061 gnd.n4865 gnd.n4864 0.152939
R14062 gnd.n4864 gnd.n3404 0.152939
R14063 gnd.n4901 gnd.n3404 0.152939
R14064 gnd.n4902 gnd.n4901 0.152939
R14065 gnd.n4910 gnd.n4902 0.152939
R14066 gnd.n4910 gnd.n4909 0.152939
R14067 gnd.n4909 gnd.n4908 0.152939
R14068 gnd.n4908 gnd.n4903 0.152939
R14069 gnd.n4903 gnd.n3369 0.152939
R14070 gnd.n4958 gnd.n3369 0.152939
R14071 gnd.n4959 gnd.n4958 0.152939
R14072 gnd.n4960 gnd.n4959 0.152939
R14073 gnd.n4960 gnd.n3367 0.152939
R14074 gnd.n4966 gnd.n3367 0.152939
R14075 gnd.n4967 gnd.n4966 0.152939
R14076 gnd.n4968 gnd.n4967 0.152939
R14077 gnd.n4968 gnd.n3365 0.152939
R14078 gnd.n4974 gnd.n3365 0.152939
R14079 gnd.n4975 gnd.n4974 0.152939
R14080 gnd.n4976 gnd.n4975 0.152939
R14081 gnd.n4976 gnd.n3363 0.152939
R14082 gnd.n4982 gnd.n3363 0.152939
R14083 gnd.n4983 gnd.n4982 0.152939
R14084 gnd.n4984 gnd.n4983 0.152939
R14085 gnd.n4984 gnd.n3361 0.152939
R14086 gnd.n4990 gnd.n3361 0.152939
R14087 gnd.n4991 gnd.n4990 0.152939
R14088 gnd.n5171 gnd.n4991 0.152939
R14089 gnd.n5171 gnd.n5170 0.152939
R14090 gnd.n4258 gnd.n4257 0.152939
R14091 gnd.n4257 gnd.n3806 0.152939
R14092 gnd.n4253 gnd.n3806 0.152939
R14093 gnd.n4253 gnd.n3782 0.152939
R14094 gnd.n4286 gnd.n3782 0.152939
R14095 gnd.n4287 gnd.n4286 0.152939
R14096 gnd.n4288 gnd.n4287 0.152939
R14097 gnd.n4288 gnd.n3772 0.152939
R14098 gnd.n4328 gnd.n3772 0.152939
R14099 gnd.n4328 gnd.n4327 0.152939
R14100 gnd.n4327 gnd.n4326 0.152939
R14101 gnd.n4326 gnd.n3773 0.152939
R14102 gnd.n4322 gnd.n3773 0.152939
R14103 gnd.n4322 gnd.n4321 0.152939
R14104 gnd.n4321 gnd.n4320 0.152939
R14105 gnd.n4320 gnd.n3777 0.152939
R14106 gnd.n4316 gnd.n3777 0.152939
R14107 gnd.n4316 gnd.n2581 0.152939
R14108 gnd.n6157 gnd.n2581 0.152939
R14109 gnd.n6157 gnd.n6156 0.152939
R14110 gnd.n6144 gnd.n2605 0.152939
R14111 gnd.n6144 gnd.n6143 0.152939
R14112 gnd.n6143 gnd.n6142 0.152939
R14113 gnd.n6142 gnd.n2607 0.152939
R14114 gnd.n6138 gnd.n2607 0.152939
R14115 gnd.n6138 gnd.n6137 0.152939
R14116 gnd.n4378 gnd.n4377 0.152939
R14117 gnd.n4378 gnd.n3736 0.152939
R14118 gnd.n4407 gnd.n3736 0.152939
R14119 gnd.n4408 gnd.n4407 0.152939
R14120 gnd.n4410 gnd.n4408 0.152939
R14121 gnd.n4410 gnd.n4409 0.152939
R14122 gnd.n4409 gnd.n3711 0.152939
R14123 gnd.n4437 gnd.n3711 0.152939
R14124 gnd.n4438 gnd.n4437 0.152939
R14125 gnd.n4440 gnd.n4438 0.152939
R14126 gnd.n4440 gnd.n4439 0.152939
R14127 gnd.n4439 gnd.n3686 0.152939
R14128 gnd.n4477 gnd.n3686 0.152939
R14129 gnd.n4478 gnd.n4477 0.152939
R14130 gnd.n4480 gnd.n4478 0.152939
R14131 gnd.n4480 gnd.n4479 0.152939
R14132 gnd.n4479 gnd.n2919 0.152939
R14133 gnd.n5956 gnd.n2919 0.152939
R14134 gnd.n5956 gnd.n5955 0.152939
R14135 gnd.n5955 gnd.n5954 0.152939
R14136 gnd.n5954 gnd.n2920 0.152939
R14137 gnd.n5950 gnd.n2920 0.152939
R14138 gnd.n5950 gnd.n5949 0.152939
R14139 gnd.n5949 gnd.n5948 0.152939
R14140 gnd.n5948 gnd.n2925 0.152939
R14141 gnd.n5944 gnd.n2925 0.152939
R14142 gnd.n5944 gnd.n5943 0.152939
R14143 gnd.n5943 gnd.n5942 0.152939
R14144 gnd.n5942 gnd.n2930 0.152939
R14145 gnd.n5938 gnd.n2930 0.152939
R14146 gnd.n5938 gnd.n5937 0.152939
R14147 gnd.n5937 gnd.n5936 0.152939
R14148 gnd.n5936 gnd.n2935 0.152939
R14149 gnd.n5932 gnd.n2935 0.152939
R14150 gnd.n5932 gnd.n5931 0.152939
R14151 gnd.n5931 gnd.n5930 0.152939
R14152 gnd.n5930 gnd.n2940 0.152939
R14153 gnd.n5926 gnd.n2940 0.152939
R14154 gnd.n5926 gnd.n5925 0.152939
R14155 gnd.n5925 gnd.n5924 0.152939
R14156 gnd.n5924 gnd.n2945 0.152939
R14157 gnd.n5920 gnd.n2945 0.152939
R14158 gnd.n5920 gnd.n5919 0.152939
R14159 gnd.n5919 gnd.n5918 0.152939
R14160 gnd.n5918 gnd.n2950 0.152939
R14161 gnd.n5914 gnd.n2950 0.152939
R14162 gnd.n5914 gnd.n5913 0.152939
R14163 gnd.n5913 gnd.n5912 0.152939
R14164 gnd.n5912 gnd.n2955 0.152939
R14165 gnd.n5908 gnd.n2955 0.152939
R14166 gnd.n5908 gnd.n5907 0.152939
R14167 gnd.n5907 gnd.n5906 0.152939
R14168 gnd.n5906 gnd.n2960 0.152939
R14169 gnd.n5902 gnd.n2960 0.152939
R14170 gnd.n5902 gnd.n5901 0.152939
R14171 gnd.n5901 gnd.n5900 0.152939
R14172 gnd.n5900 gnd.n2965 0.152939
R14173 gnd.n5896 gnd.n2965 0.152939
R14174 gnd.n5896 gnd.n5895 0.152939
R14175 gnd.n5895 gnd.n5894 0.152939
R14176 gnd.n5894 gnd.n2970 0.152939
R14177 gnd.n5890 gnd.n2970 0.152939
R14178 gnd.n5890 gnd.n5889 0.152939
R14179 gnd.n5889 gnd.n5888 0.152939
R14180 gnd.n5888 gnd.n2975 0.152939
R14181 gnd.n5884 gnd.n2975 0.152939
R14182 gnd.n5884 gnd.n5883 0.152939
R14183 gnd.n5883 gnd.n5882 0.152939
R14184 gnd.n5882 gnd.n2980 0.152939
R14185 gnd.n5878 gnd.n2980 0.152939
R14186 gnd.n5878 gnd.n5877 0.152939
R14187 gnd.n5877 gnd.n5876 0.152939
R14188 gnd.n5876 gnd.n2985 0.152939
R14189 gnd.n5872 gnd.n2985 0.152939
R14190 gnd.n5872 gnd.n5871 0.152939
R14191 gnd.n5871 gnd.n5870 0.152939
R14192 gnd.n5870 gnd.n2990 0.152939
R14193 gnd.n5866 gnd.n2990 0.152939
R14194 gnd.n5866 gnd.n5865 0.152939
R14195 gnd.n5865 gnd.n5864 0.152939
R14196 gnd.n5864 gnd.n2995 0.152939
R14197 gnd.n2998 gnd.n2995 0.152939
R14198 gnd.n5057 gnd.n5056 0.152939
R14199 gnd.n5057 gnd.n5052 0.152939
R14200 gnd.n5065 gnd.n5052 0.152939
R14201 gnd.n5066 gnd.n5065 0.152939
R14202 gnd.n5068 gnd.n5066 0.152939
R14203 gnd.n5068 gnd.n5067 0.152939
R14204 gnd.n4997 gnd.n4992 0.152939
R14205 gnd.n4992 gnd.n3225 0.152939
R14206 gnd.n5575 gnd.n3225 0.152939
R14207 gnd.n5576 gnd.n5575 0.152939
R14208 gnd.n5577 gnd.n5576 0.152939
R14209 gnd.n5577 gnd.n3220 0.152939
R14210 gnd.n5597 gnd.n3220 0.152939
R14211 gnd.n5597 gnd.n5596 0.152939
R14212 gnd.n5596 gnd.n5595 0.152939
R14213 gnd.n5595 gnd.n3221 0.152939
R14214 gnd.n5591 gnd.n3221 0.152939
R14215 gnd.n5591 gnd.n3208 0.152939
R14216 gnd.n5655 gnd.n3208 0.152939
R14217 gnd.n5656 gnd.n5655 0.152939
R14218 gnd.n5667 gnd.n5656 0.152939
R14219 gnd.n5667 gnd.n5666 0.152939
R14220 gnd.n5666 gnd.n5665 0.152939
R14221 gnd.n5665 gnd.n5657 0.152939
R14222 gnd.n5661 gnd.n5657 0.152939
R14223 gnd.n5661 gnd.n63 0.152939
R14224 gnd.n7546 gnd.n7545 0.145814
R14225 gnd.n4259 gnd.n3803 0.145814
R14226 gnd.n4259 gnd.n4258 0.145814
R14227 gnd.n7546 gnd.n63 0.145814
R14228 gnd.n6137 gnd.n6136 0.128549
R14229 gnd.n5067 gnd.n3229 0.128549
R14230 gnd.n1154 gnd.n0 0.127478
R14231 gnd.n3147 gnd.n79 0.10111
R14232 gnd.n4275 gnd.n4274 0.10111
R14233 gnd.n1734 gnd.n1733 0.0767195
R14234 gnd.n1733 gnd.n1732 0.0767195
R14235 gnd.n6136 gnd.n2577 0.063
R14236 gnd.n5564 gnd.n3229 0.063
R14237 gnd.n5566 gnd.n5564 0.0538288
R14238 gnd.n7482 gnd.n174 0.0538288
R14239 gnd.n4124 gnd.n4122 0.0538288
R14240 gnd.n6164 gnd.n2577 0.0538288
R14241 gnd.n4276 gnd.n4275 0.0523293
R14242 gnd.n5634 gnd.n79 0.0523293
R14243 gnd.n2302 gnd.n918 0.0477147
R14244 gnd.n1497 gnd.n1385 0.0442063
R14245 gnd.n1498 gnd.n1497 0.0442063
R14246 gnd.n1499 gnd.n1498 0.0442063
R14247 gnd.n1499 gnd.n1374 0.0442063
R14248 gnd.n1513 gnd.n1374 0.0442063
R14249 gnd.n1514 gnd.n1513 0.0442063
R14250 gnd.n1515 gnd.n1514 0.0442063
R14251 gnd.n1515 gnd.n1361 0.0442063
R14252 gnd.n1559 gnd.n1361 0.0442063
R14253 gnd.n1560 gnd.n1559 0.0442063
R14254 gnd.n1562 gnd.n1295 0.0344674
R14255 gnd.n5567 gnd.n5566 0.0344674
R14256 gnd.n5567 gnd.n3039 0.0344674
R14257 gnd.n3040 gnd.n3039 0.0344674
R14258 gnd.n3041 gnd.n3040 0.0344674
R14259 gnd.n3223 gnd.n3041 0.0344674
R14260 gnd.n3223 gnd.n3059 0.0344674
R14261 gnd.n3060 gnd.n3059 0.0344674
R14262 gnd.n3061 gnd.n3060 0.0344674
R14263 gnd.n5586 gnd.n3061 0.0344674
R14264 gnd.n5586 gnd.n3080 0.0344674
R14265 gnd.n3081 gnd.n3080 0.0344674
R14266 gnd.n3082 gnd.n3081 0.0344674
R14267 gnd.n5649 gnd.n3082 0.0344674
R14268 gnd.n5649 gnd.n3099 0.0344674
R14269 gnd.n3100 gnd.n3099 0.0344674
R14270 gnd.n3101 gnd.n3100 0.0344674
R14271 gnd.n3203 gnd.n3101 0.0344674
R14272 gnd.n5678 gnd.n3203 0.0344674
R14273 gnd.n5683 gnd.n5678 0.0344674
R14274 gnd.n5684 gnd.n5683 0.0344674
R14275 gnd.n5684 gnd.n3133 0.0344674
R14276 gnd.n3134 gnd.n3133 0.0344674
R14277 gnd.n3135 gnd.n3134 0.0344674
R14278 gnd.n3136 gnd.n3135 0.0344674
R14279 gnd.n5692 gnd.n3136 0.0344674
R14280 gnd.n5692 gnd.n93 0.0344674
R14281 gnd.n94 gnd.n93 0.0344674
R14282 gnd.n95 gnd.n94 0.0344674
R14283 gnd.n3198 gnd.n95 0.0344674
R14284 gnd.n3198 gnd.n112 0.0344674
R14285 gnd.n113 gnd.n112 0.0344674
R14286 gnd.n114 gnd.n113 0.0344674
R14287 gnd.n5718 gnd.n114 0.0344674
R14288 gnd.n5718 gnd.n133 0.0344674
R14289 gnd.n134 gnd.n133 0.0344674
R14290 gnd.n135 gnd.n134 0.0344674
R14291 gnd.n5725 gnd.n135 0.0344674
R14292 gnd.n5725 gnd.n154 0.0344674
R14293 gnd.n155 gnd.n154 0.0344674
R14294 gnd.n156 gnd.n155 0.0344674
R14295 gnd.n173 gnd.n156 0.0344674
R14296 gnd.n7482 gnd.n173 0.0344674
R14297 gnd.n4125 gnd.n4124 0.0344674
R14298 gnd.n4125 gnd.n2381 0.0344674
R14299 gnd.n2382 gnd.n2381 0.0344674
R14300 gnd.n2383 gnd.n2382 0.0344674
R14301 gnd.n4128 gnd.n2383 0.0344674
R14302 gnd.n4128 gnd.n2402 0.0344674
R14303 gnd.n2403 gnd.n2402 0.0344674
R14304 gnd.n2404 gnd.n2403 0.0344674
R14305 gnd.n4135 gnd.n2404 0.0344674
R14306 gnd.n4135 gnd.n2423 0.0344674
R14307 gnd.n2424 gnd.n2423 0.0344674
R14308 gnd.n2425 gnd.n2424 0.0344674
R14309 gnd.n3814 gnd.n2425 0.0344674
R14310 gnd.n3814 gnd.n2443 0.0344674
R14311 gnd.n2444 gnd.n2443 0.0344674
R14312 gnd.n2445 gnd.n2444 0.0344674
R14313 gnd.n3809 gnd.n2445 0.0344674
R14314 gnd.n3809 gnd.n2462 0.0344674
R14315 gnd.n2463 gnd.n2462 0.0344674
R14316 gnd.n2464 gnd.n2463 0.0344674
R14317 gnd.n4226 gnd.n2464 0.0344674
R14318 gnd.n4226 gnd.n2478 0.0344674
R14319 gnd.n2479 gnd.n2478 0.0344674
R14320 gnd.n2480 gnd.n2479 0.0344674
R14321 gnd.n4246 gnd.n2480 0.0344674
R14322 gnd.n4246 gnd.n2496 0.0344674
R14323 gnd.n2497 gnd.n2496 0.0344674
R14324 gnd.n2498 gnd.n2497 0.0344674
R14325 gnd.n3780 gnd.n2498 0.0344674
R14326 gnd.n3780 gnd.n2515 0.0344674
R14327 gnd.n2516 gnd.n2515 0.0344674
R14328 gnd.n2517 gnd.n2516 0.0344674
R14329 gnd.n4297 gnd.n2517 0.0344674
R14330 gnd.n4297 gnd.n2536 0.0344674
R14331 gnd.n2537 gnd.n2536 0.0344674
R14332 gnd.n2538 gnd.n2537 0.0344674
R14333 gnd.n4307 gnd.n2538 0.0344674
R14334 gnd.n4307 gnd.n2556 0.0344674
R14335 gnd.n2557 gnd.n2556 0.0344674
R14336 gnd.n2558 gnd.n2557 0.0344674
R14337 gnd.n2576 gnd.n2558 0.0344674
R14338 gnd.n6164 gnd.n2576 0.0344674
R14339 gnd.n6135 gnd.n2612 0.0344674
R14340 gnd.n5077 gnd.n5076 0.0344674
R14341 gnd.n6155 gnd.n6154 0.029712
R14342 gnd.n5007 gnd.n4998 0.029712
R14343 gnd.n1582 gnd.n1581 0.0269946
R14344 gnd.n1584 gnd.n1583 0.0269946
R14345 gnd.n1290 gnd.n1288 0.0269946
R14346 gnd.n1594 gnd.n1592 0.0269946
R14347 gnd.n1593 gnd.n1269 0.0269946
R14348 gnd.n1613 gnd.n1612 0.0269946
R14349 gnd.n1615 gnd.n1614 0.0269946
R14350 gnd.n1264 gnd.n1263 0.0269946
R14351 gnd.n1625 gnd.n1259 0.0269946
R14352 gnd.n1624 gnd.n1261 0.0269946
R14353 gnd.n1260 gnd.n1242 0.0269946
R14354 gnd.n1645 gnd.n1243 0.0269946
R14355 gnd.n1644 gnd.n1244 0.0269946
R14356 gnd.n1678 gnd.n1219 0.0269946
R14357 gnd.n1680 gnd.n1679 0.0269946
R14358 gnd.n1681 gnd.n1166 0.0269946
R14359 gnd.n1214 gnd.n1167 0.0269946
R14360 gnd.n1216 gnd.n1168 0.0269946
R14361 gnd.n1691 gnd.n1690 0.0269946
R14362 gnd.n1693 gnd.n1692 0.0269946
R14363 gnd.n1694 gnd.n1188 0.0269946
R14364 gnd.n1696 gnd.n1189 0.0269946
R14365 gnd.n1699 gnd.n1190 0.0269946
R14366 gnd.n1702 gnd.n1701 0.0269946
R14367 gnd.n1704 gnd.n1703 0.0269946
R14368 gnd.n1769 gnd.n1089 0.0269946
R14369 gnd.n1771 gnd.n1770 0.0269946
R14370 gnd.n1780 gnd.n1082 0.0269946
R14371 gnd.n1782 gnd.n1781 0.0269946
R14372 gnd.n1783 gnd.n1080 0.0269946
R14373 gnd.n1790 gnd.n1786 0.0269946
R14374 gnd.n1789 gnd.n1788 0.0269946
R14375 gnd.n1787 gnd.n1059 0.0269946
R14376 gnd.n1812 gnd.n1060 0.0269946
R14377 gnd.n1811 gnd.n1061 0.0269946
R14378 gnd.n1856 gnd.n1036 0.0269946
R14379 gnd.n1858 gnd.n1857 0.0269946
R14380 gnd.n1867 gnd.n1029 0.0269946
R14381 gnd.n1869 gnd.n1868 0.0269946
R14382 gnd.n1870 gnd.n1027 0.0269946
R14383 gnd.n1877 gnd.n1873 0.0269946
R14384 gnd.n1876 gnd.n1875 0.0269946
R14385 gnd.n1874 gnd.n1006 0.0269946
R14386 gnd.n1899 gnd.n1007 0.0269946
R14387 gnd.n1898 gnd.n1008 0.0269946
R14388 gnd.n1945 gnd.n982 0.0269946
R14389 gnd.n1947 gnd.n1946 0.0269946
R14390 gnd.n1956 gnd.n975 0.0269946
R14391 gnd.n2215 gnd.n973 0.0269946
R14392 gnd.n2220 gnd.n2218 0.0269946
R14393 gnd.n2219 gnd.n954 0.0269946
R14394 gnd.n2244 gnd.n2243 0.0269946
R14395 gnd.n6131 gnd.n2618 0.0225788
R14396 gnd.n6130 gnd.n2619 0.0225788
R14397 gnd.n6127 gnd.n6126 0.0225788
R14398 gnd.n6123 gnd.n2624 0.0225788
R14399 gnd.n6122 gnd.n2630 0.0225788
R14400 gnd.n6119 gnd.n6118 0.0225788
R14401 gnd.n6115 gnd.n2634 0.0225788
R14402 gnd.n6114 gnd.n2638 0.0225788
R14403 gnd.n6111 gnd.n6110 0.0225788
R14404 gnd.n6107 gnd.n2642 0.0225788
R14405 gnd.n6106 gnd.n2648 0.0225788
R14406 gnd.n6103 gnd.n6102 0.0225788
R14407 gnd.n6099 gnd.n2652 0.0225788
R14408 gnd.n6098 gnd.n2656 0.0225788
R14409 gnd.n6095 gnd.n6094 0.0225788
R14410 gnd.n6091 gnd.n2660 0.0225788
R14411 gnd.n6090 gnd.n2669 0.0225788
R14412 gnd.n2674 gnd.n2673 0.0225788
R14413 gnd.n6154 gnd.n2583 0.0225788
R14414 gnd.n5083 gnd.n5081 0.0225788
R14415 gnd.n5082 gnd.n5044 0.0225788
R14416 gnd.n5092 gnd.n5091 0.0225788
R14417 gnd.n5045 gnd.n5040 0.0225788
R14418 gnd.n5102 gnd.n5100 0.0225788
R14419 gnd.n5101 gnd.n5035 0.0225788
R14420 gnd.n5111 gnd.n5110 0.0225788
R14421 gnd.n5036 gnd.n5031 0.0225788
R14422 gnd.n5121 gnd.n5119 0.0225788
R14423 gnd.n5120 gnd.n5026 0.0225788
R14424 gnd.n5130 gnd.n5129 0.0225788
R14425 gnd.n5027 gnd.n5022 0.0225788
R14426 gnd.n5140 gnd.n5138 0.0225788
R14427 gnd.n5139 gnd.n5017 0.0225788
R14428 gnd.n5150 gnd.n5149 0.0225788
R14429 gnd.n5146 gnd.n5018 0.0225788
R14430 gnd.n5160 gnd.n5005 0.0225788
R14431 gnd.n5159 gnd.n5006 0.0225788
R14432 gnd.n5008 gnd.n5007 0.0225788
R14433 gnd.n5169 gnd.n4998 0.0218415
R14434 gnd.n6155 gnd.n2582 0.0218415
R14435 gnd.n1562 gnd.n1561 0.0202011
R14436 gnd.n1561 gnd.n1560 0.0148637
R14437 gnd.n2213 gnd.n1957 0.0144266
R14438 gnd.n2214 gnd.n2213 0.0130679
R14439 gnd.n2618 gnd.n2612 0.0123886
R14440 gnd.n6131 gnd.n6130 0.0123886
R14441 gnd.n6127 gnd.n2619 0.0123886
R14442 gnd.n6126 gnd.n2624 0.0123886
R14443 gnd.n6123 gnd.n6122 0.0123886
R14444 gnd.n6119 gnd.n2630 0.0123886
R14445 gnd.n6118 gnd.n2634 0.0123886
R14446 gnd.n6115 gnd.n6114 0.0123886
R14447 gnd.n6111 gnd.n2638 0.0123886
R14448 gnd.n6110 gnd.n2642 0.0123886
R14449 gnd.n6107 gnd.n6106 0.0123886
R14450 gnd.n6103 gnd.n2648 0.0123886
R14451 gnd.n6102 gnd.n2652 0.0123886
R14452 gnd.n6099 gnd.n6098 0.0123886
R14453 gnd.n6095 gnd.n2656 0.0123886
R14454 gnd.n6094 gnd.n2660 0.0123886
R14455 gnd.n6091 gnd.n6090 0.0123886
R14456 gnd.n2674 gnd.n2669 0.0123886
R14457 gnd.n2673 gnd.n2583 0.0123886
R14458 gnd.n5081 gnd.n5077 0.0123886
R14459 gnd.n5083 gnd.n5082 0.0123886
R14460 gnd.n5092 gnd.n5044 0.0123886
R14461 gnd.n5091 gnd.n5045 0.0123886
R14462 gnd.n5100 gnd.n5040 0.0123886
R14463 gnd.n5102 gnd.n5101 0.0123886
R14464 gnd.n5111 gnd.n5035 0.0123886
R14465 gnd.n5110 gnd.n5036 0.0123886
R14466 gnd.n5119 gnd.n5031 0.0123886
R14467 gnd.n5121 gnd.n5120 0.0123886
R14468 gnd.n5130 gnd.n5026 0.0123886
R14469 gnd.n5129 gnd.n5027 0.0123886
R14470 gnd.n5138 gnd.n5022 0.0123886
R14471 gnd.n5140 gnd.n5139 0.0123886
R14472 gnd.n5150 gnd.n5017 0.0123886
R14473 gnd.n5149 gnd.n5018 0.0123886
R14474 gnd.n5146 gnd.n5005 0.0123886
R14475 gnd.n5160 gnd.n5159 0.0123886
R14476 gnd.n5008 gnd.n5006 0.0123886
R14477 gnd.n1581 gnd.n1295 0.00797283
R14478 gnd.n1583 gnd.n1582 0.00797283
R14479 gnd.n1584 gnd.n1290 0.00797283
R14480 gnd.n1592 gnd.n1288 0.00797283
R14481 gnd.n1594 gnd.n1593 0.00797283
R14482 gnd.n1612 gnd.n1269 0.00797283
R14483 gnd.n1614 gnd.n1613 0.00797283
R14484 gnd.n1615 gnd.n1264 0.00797283
R14485 gnd.n1263 gnd.n1259 0.00797283
R14486 gnd.n1625 gnd.n1624 0.00797283
R14487 gnd.n1261 gnd.n1260 0.00797283
R14488 gnd.n1243 gnd.n1242 0.00797283
R14489 gnd.n1645 gnd.n1644 0.00797283
R14490 gnd.n1244 gnd.n1219 0.00797283
R14491 gnd.n1679 gnd.n1678 0.00797283
R14492 gnd.n1681 gnd.n1680 0.00797283
R14493 gnd.n1214 gnd.n1166 0.00797283
R14494 gnd.n1216 gnd.n1167 0.00797283
R14495 gnd.n1690 gnd.n1168 0.00797283
R14496 gnd.n1692 gnd.n1691 0.00797283
R14497 gnd.n1694 gnd.n1693 0.00797283
R14498 gnd.n1696 gnd.n1188 0.00797283
R14499 gnd.n1699 gnd.n1189 0.00797283
R14500 gnd.n1701 gnd.n1190 0.00797283
R14501 gnd.n1704 gnd.n1702 0.00797283
R14502 gnd.n1703 gnd.n1089 0.00797283
R14503 gnd.n1771 gnd.n1769 0.00797283
R14504 gnd.n1770 gnd.n1082 0.00797283
R14505 gnd.n1781 gnd.n1780 0.00797283
R14506 gnd.n1783 gnd.n1782 0.00797283
R14507 gnd.n1786 gnd.n1080 0.00797283
R14508 gnd.n1790 gnd.n1789 0.00797283
R14509 gnd.n1788 gnd.n1787 0.00797283
R14510 gnd.n1060 gnd.n1059 0.00797283
R14511 gnd.n1812 gnd.n1811 0.00797283
R14512 gnd.n1061 gnd.n1036 0.00797283
R14513 gnd.n1858 gnd.n1856 0.00797283
R14514 gnd.n1857 gnd.n1029 0.00797283
R14515 gnd.n1868 gnd.n1867 0.00797283
R14516 gnd.n1870 gnd.n1869 0.00797283
R14517 gnd.n1873 gnd.n1027 0.00797283
R14518 gnd.n1877 gnd.n1876 0.00797283
R14519 gnd.n1875 gnd.n1874 0.00797283
R14520 gnd.n1007 gnd.n1006 0.00797283
R14521 gnd.n1899 gnd.n1898 0.00797283
R14522 gnd.n1008 gnd.n982 0.00797283
R14523 gnd.n1947 gnd.n1945 0.00797283
R14524 gnd.n1946 gnd.n975 0.00797283
R14525 gnd.n1957 gnd.n1956 0.00797283
R14526 gnd.n2215 gnd.n2214 0.00797283
R14527 gnd.n2218 gnd.n973 0.00797283
R14528 gnd.n2220 gnd.n2219 0.00797283
R14529 gnd.n2243 gnd.n954 0.00797283
R14530 gnd.n2244 gnd.n918 0.00797283
R14531 gnd.n6136 gnd.n6135 0.00593478
R14532 gnd.n5076 gnd.n3229 0.00593478
R14533 commonsourceibias.n25 commonsourceibias.t22 230.006
R14534 commonsourceibias.n91 commonsourceibias.t73 230.006
R14535 commonsourceibias.n218 commonsourceibias.t98 230.006
R14536 commonsourceibias.n154 commonsourceibias.t70 230.006
R14537 commonsourceibias.n322 commonsourceibias.t40 230.006
R14538 commonsourceibias.n281 commonsourceibias.t111 230.006
R14539 commonsourceibias.n483 commonsourceibias.t113 230.006
R14540 commonsourceibias.n419 commonsourceibias.t52 230.006
R14541 commonsourceibias.n70 commonsourceibias.t8 207.983
R14542 commonsourceibias.n136 commonsourceibias.t89 207.983
R14543 commonsourceibias.n263 commonsourceibias.t109 207.983
R14544 commonsourceibias.n199 commonsourceibias.t54 207.983
R14545 commonsourceibias.n368 commonsourceibias.t26 207.983
R14546 commonsourceibias.n402 commonsourceibias.t69 207.983
R14547 commonsourceibias.n529 commonsourceibias.t63 207.983
R14548 commonsourceibias.n465 commonsourceibias.t112 207.983
R14549 commonsourceibias.n10 commonsourceibias.t38 168.701
R14550 commonsourceibias.n63 commonsourceibias.t0 168.701
R14551 commonsourceibias.n57 commonsourceibias.t6 168.701
R14552 commonsourceibias.n16 commonsourceibias.t44 168.701
R14553 commonsourceibias.n49 commonsourceibias.t12 168.701
R14554 commonsourceibias.n43 commonsourceibias.t20 168.701
R14555 commonsourceibias.n19 commonsourceibias.t2 168.701
R14556 commonsourceibias.n21 commonsourceibias.t10 168.701
R14557 commonsourceibias.n23 commonsourceibias.t34 168.701
R14558 commonsourceibias.n26 commonsourceibias.t16 168.701
R14559 commonsourceibias.n1 commonsourceibias.t51 168.701
R14560 commonsourceibias.n129 commonsourceibias.t95 168.701
R14561 commonsourceibias.n123 commonsourceibias.t90 168.701
R14562 commonsourceibias.n7 commonsourceibias.t101 168.701
R14563 commonsourceibias.n115 commonsourceibias.t86 168.701
R14564 commonsourceibias.n109 commonsourceibias.t77 168.701
R14565 commonsourceibias.n85 commonsourceibias.t94 168.701
R14566 commonsourceibias.n87 commonsourceibias.t87 168.701
R14567 commonsourceibias.n89 commonsourceibias.t58 168.701
R14568 commonsourceibias.n92 commonsourceibias.t80 168.701
R14569 commonsourceibias.n219 commonsourceibias.t102 168.701
R14570 commonsourceibias.n216 commonsourceibias.t48 168.701
R14571 commonsourceibias.n214 commonsourceibias.t103 168.701
R14572 commonsourceibias.n212 commonsourceibias.t108 168.701
R14573 commonsourceibias.n236 commonsourceibias.t88 168.701
R14574 commonsourceibias.n242 commonsourceibias.t68 168.701
R14575 commonsourceibias.n209 commonsourceibias.t115 168.701
R14576 commonsourceibias.n250 commonsourceibias.t93 168.701
R14577 commonsourceibias.n256 commonsourceibias.t96 168.701
R14578 commonsourceibias.n203 commonsourceibias.t57 168.701
R14579 commonsourceibias.n139 commonsourceibias.t119 168.701
R14580 commonsourceibias.n192 commonsourceibias.t110 168.701
R14581 commonsourceibias.n186 commonsourceibias.t60 168.701
R14582 commonsourceibias.n145 commonsourceibias.t117 168.701
R14583 commonsourceibias.n178 commonsourceibias.t65 168.701
R14584 commonsourceibias.n172 commonsourceibias.t59 168.701
R14585 commonsourceibias.n148 commonsourceibias.t118 168.701
R14586 commonsourceibias.n150 commonsourceibias.t71 168.701
R14587 commonsourceibias.n152 commonsourceibias.t83 168.701
R14588 commonsourceibias.n155 commonsourceibias.t116 168.701
R14589 commonsourceibias.n323 commonsourceibias.t32 168.701
R14590 commonsourceibias.n320 commonsourceibias.t42 168.701
R14591 commonsourceibias.n318 commonsourceibias.t28 168.701
R14592 commonsourceibias.n316 commonsourceibias.t18 168.701
R14593 commonsourceibias.n340 commonsourceibias.t36 168.701
R14594 commonsourceibias.n346 commonsourceibias.t30 168.701
R14595 commonsourceibias.n348 commonsourceibias.t4 168.701
R14596 commonsourceibias.n355 commonsourceibias.t24 168.701
R14597 commonsourceibias.n361 commonsourceibias.t14 168.701
R14598 commonsourceibias.n308 commonsourceibias.t46 168.701
R14599 commonsourceibias.n267 commonsourceibias.t99 168.701
R14600 commonsourceibias.n395 commonsourceibias.t84 168.701
R14601 commonsourceibias.n389 commonsourceibias.t72 168.701
R14602 commonsourceibias.n382 commonsourceibias.t92 168.701
R14603 commonsourceibias.n380 commonsourceibias.t66 168.701
R14604 commonsourceibias.n282 commonsourceibias.t64 168.701
R14605 commonsourceibias.n279 commonsourceibias.t104 168.701
R14606 commonsourceibias.n277 commonsourceibias.t67 168.701
R14607 commonsourceibias.n275 commonsourceibias.t79 168.701
R14608 commonsourceibias.n299 commonsourceibias.t56 168.701
R14609 commonsourceibias.n484 commonsourceibias.t97 168.701
R14610 commonsourceibias.n481 commonsourceibias.t78 168.701
R14611 commonsourceibias.n479 commonsourceibias.t53 168.701
R14612 commonsourceibias.n477 commonsourceibias.t62 168.701
R14613 commonsourceibias.n501 commonsourceibias.t82 168.701
R14614 commonsourceibias.n507 commonsourceibias.t85 168.701
R14615 commonsourceibias.n509 commonsourceibias.t76 168.701
R14616 commonsourceibias.n516 commonsourceibias.t100 168.701
R14617 commonsourceibias.n522 commonsourceibias.t91 168.701
R14618 commonsourceibias.n469 commonsourceibias.t81 168.701
R14619 commonsourceibias.n420 commonsourceibias.t61 168.701
R14620 commonsourceibias.n417 commonsourceibias.t75 168.701
R14621 commonsourceibias.n415 commonsourceibias.t55 168.701
R14622 commonsourceibias.n413 commonsourceibias.t105 168.701
R14623 commonsourceibias.n437 commonsourceibias.t74 168.701
R14624 commonsourceibias.n443 commonsourceibias.t49 168.701
R14625 commonsourceibias.n445 commonsourceibias.t106 168.701
R14626 commonsourceibias.n452 commonsourceibias.t114 168.701
R14627 commonsourceibias.n458 commonsourceibias.t50 168.701
R14628 commonsourceibias.n405 commonsourceibias.t107 168.701
R14629 commonsourceibias.n27 commonsourceibias.n24 161.3
R14630 commonsourceibias.n29 commonsourceibias.n28 161.3
R14631 commonsourceibias.n31 commonsourceibias.n30 161.3
R14632 commonsourceibias.n32 commonsourceibias.n22 161.3
R14633 commonsourceibias.n34 commonsourceibias.n33 161.3
R14634 commonsourceibias.n36 commonsourceibias.n35 161.3
R14635 commonsourceibias.n37 commonsourceibias.n20 161.3
R14636 commonsourceibias.n39 commonsourceibias.n38 161.3
R14637 commonsourceibias.n41 commonsourceibias.n40 161.3
R14638 commonsourceibias.n42 commonsourceibias.n18 161.3
R14639 commonsourceibias.n45 commonsourceibias.n44 161.3
R14640 commonsourceibias.n46 commonsourceibias.n17 161.3
R14641 commonsourceibias.n48 commonsourceibias.n47 161.3
R14642 commonsourceibias.n50 commonsourceibias.n15 161.3
R14643 commonsourceibias.n52 commonsourceibias.n51 161.3
R14644 commonsourceibias.n53 commonsourceibias.n14 161.3
R14645 commonsourceibias.n55 commonsourceibias.n54 161.3
R14646 commonsourceibias.n56 commonsourceibias.n13 161.3
R14647 commonsourceibias.n59 commonsourceibias.n58 161.3
R14648 commonsourceibias.n60 commonsourceibias.n12 161.3
R14649 commonsourceibias.n62 commonsourceibias.n61 161.3
R14650 commonsourceibias.n64 commonsourceibias.n11 161.3
R14651 commonsourceibias.n66 commonsourceibias.n65 161.3
R14652 commonsourceibias.n68 commonsourceibias.n67 161.3
R14653 commonsourceibias.n69 commonsourceibias.n9 161.3
R14654 commonsourceibias.n93 commonsourceibias.n90 161.3
R14655 commonsourceibias.n95 commonsourceibias.n94 161.3
R14656 commonsourceibias.n97 commonsourceibias.n96 161.3
R14657 commonsourceibias.n98 commonsourceibias.n88 161.3
R14658 commonsourceibias.n100 commonsourceibias.n99 161.3
R14659 commonsourceibias.n102 commonsourceibias.n101 161.3
R14660 commonsourceibias.n103 commonsourceibias.n86 161.3
R14661 commonsourceibias.n105 commonsourceibias.n104 161.3
R14662 commonsourceibias.n107 commonsourceibias.n106 161.3
R14663 commonsourceibias.n108 commonsourceibias.n84 161.3
R14664 commonsourceibias.n111 commonsourceibias.n110 161.3
R14665 commonsourceibias.n112 commonsourceibias.n8 161.3
R14666 commonsourceibias.n114 commonsourceibias.n113 161.3
R14667 commonsourceibias.n116 commonsourceibias.n6 161.3
R14668 commonsourceibias.n118 commonsourceibias.n117 161.3
R14669 commonsourceibias.n119 commonsourceibias.n5 161.3
R14670 commonsourceibias.n121 commonsourceibias.n120 161.3
R14671 commonsourceibias.n122 commonsourceibias.n4 161.3
R14672 commonsourceibias.n125 commonsourceibias.n124 161.3
R14673 commonsourceibias.n126 commonsourceibias.n3 161.3
R14674 commonsourceibias.n128 commonsourceibias.n127 161.3
R14675 commonsourceibias.n130 commonsourceibias.n2 161.3
R14676 commonsourceibias.n132 commonsourceibias.n131 161.3
R14677 commonsourceibias.n134 commonsourceibias.n133 161.3
R14678 commonsourceibias.n135 commonsourceibias.n0 161.3
R14679 commonsourceibias.n262 commonsourceibias.n202 161.3
R14680 commonsourceibias.n261 commonsourceibias.n260 161.3
R14681 commonsourceibias.n259 commonsourceibias.n258 161.3
R14682 commonsourceibias.n257 commonsourceibias.n204 161.3
R14683 commonsourceibias.n255 commonsourceibias.n254 161.3
R14684 commonsourceibias.n253 commonsourceibias.n205 161.3
R14685 commonsourceibias.n252 commonsourceibias.n251 161.3
R14686 commonsourceibias.n249 commonsourceibias.n206 161.3
R14687 commonsourceibias.n248 commonsourceibias.n247 161.3
R14688 commonsourceibias.n246 commonsourceibias.n207 161.3
R14689 commonsourceibias.n245 commonsourceibias.n244 161.3
R14690 commonsourceibias.n243 commonsourceibias.n208 161.3
R14691 commonsourceibias.n241 commonsourceibias.n240 161.3
R14692 commonsourceibias.n239 commonsourceibias.n210 161.3
R14693 commonsourceibias.n238 commonsourceibias.n237 161.3
R14694 commonsourceibias.n235 commonsourceibias.n211 161.3
R14695 commonsourceibias.n234 commonsourceibias.n233 161.3
R14696 commonsourceibias.n232 commonsourceibias.n231 161.3
R14697 commonsourceibias.n230 commonsourceibias.n213 161.3
R14698 commonsourceibias.n229 commonsourceibias.n228 161.3
R14699 commonsourceibias.n227 commonsourceibias.n226 161.3
R14700 commonsourceibias.n225 commonsourceibias.n215 161.3
R14701 commonsourceibias.n224 commonsourceibias.n223 161.3
R14702 commonsourceibias.n222 commonsourceibias.n221 161.3
R14703 commonsourceibias.n220 commonsourceibias.n217 161.3
R14704 commonsourceibias.n156 commonsourceibias.n153 161.3
R14705 commonsourceibias.n158 commonsourceibias.n157 161.3
R14706 commonsourceibias.n160 commonsourceibias.n159 161.3
R14707 commonsourceibias.n161 commonsourceibias.n151 161.3
R14708 commonsourceibias.n163 commonsourceibias.n162 161.3
R14709 commonsourceibias.n165 commonsourceibias.n164 161.3
R14710 commonsourceibias.n166 commonsourceibias.n149 161.3
R14711 commonsourceibias.n168 commonsourceibias.n167 161.3
R14712 commonsourceibias.n170 commonsourceibias.n169 161.3
R14713 commonsourceibias.n171 commonsourceibias.n147 161.3
R14714 commonsourceibias.n174 commonsourceibias.n173 161.3
R14715 commonsourceibias.n175 commonsourceibias.n146 161.3
R14716 commonsourceibias.n177 commonsourceibias.n176 161.3
R14717 commonsourceibias.n179 commonsourceibias.n144 161.3
R14718 commonsourceibias.n181 commonsourceibias.n180 161.3
R14719 commonsourceibias.n182 commonsourceibias.n143 161.3
R14720 commonsourceibias.n184 commonsourceibias.n183 161.3
R14721 commonsourceibias.n185 commonsourceibias.n142 161.3
R14722 commonsourceibias.n188 commonsourceibias.n187 161.3
R14723 commonsourceibias.n189 commonsourceibias.n141 161.3
R14724 commonsourceibias.n191 commonsourceibias.n190 161.3
R14725 commonsourceibias.n193 commonsourceibias.n140 161.3
R14726 commonsourceibias.n195 commonsourceibias.n194 161.3
R14727 commonsourceibias.n197 commonsourceibias.n196 161.3
R14728 commonsourceibias.n198 commonsourceibias.n138 161.3
R14729 commonsourceibias.n367 commonsourceibias.n307 161.3
R14730 commonsourceibias.n366 commonsourceibias.n365 161.3
R14731 commonsourceibias.n364 commonsourceibias.n363 161.3
R14732 commonsourceibias.n362 commonsourceibias.n309 161.3
R14733 commonsourceibias.n360 commonsourceibias.n359 161.3
R14734 commonsourceibias.n358 commonsourceibias.n310 161.3
R14735 commonsourceibias.n357 commonsourceibias.n356 161.3
R14736 commonsourceibias.n354 commonsourceibias.n311 161.3
R14737 commonsourceibias.n353 commonsourceibias.n352 161.3
R14738 commonsourceibias.n351 commonsourceibias.n312 161.3
R14739 commonsourceibias.n350 commonsourceibias.n349 161.3
R14740 commonsourceibias.n347 commonsourceibias.n313 161.3
R14741 commonsourceibias.n345 commonsourceibias.n344 161.3
R14742 commonsourceibias.n343 commonsourceibias.n314 161.3
R14743 commonsourceibias.n342 commonsourceibias.n341 161.3
R14744 commonsourceibias.n339 commonsourceibias.n315 161.3
R14745 commonsourceibias.n338 commonsourceibias.n337 161.3
R14746 commonsourceibias.n336 commonsourceibias.n335 161.3
R14747 commonsourceibias.n334 commonsourceibias.n317 161.3
R14748 commonsourceibias.n333 commonsourceibias.n332 161.3
R14749 commonsourceibias.n331 commonsourceibias.n330 161.3
R14750 commonsourceibias.n329 commonsourceibias.n319 161.3
R14751 commonsourceibias.n328 commonsourceibias.n327 161.3
R14752 commonsourceibias.n326 commonsourceibias.n325 161.3
R14753 commonsourceibias.n324 commonsourceibias.n321 161.3
R14754 commonsourceibias.n301 commonsourceibias.n300 161.3
R14755 commonsourceibias.n298 commonsourceibias.n274 161.3
R14756 commonsourceibias.n297 commonsourceibias.n296 161.3
R14757 commonsourceibias.n295 commonsourceibias.n294 161.3
R14758 commonsourceibias.n293 commonsourceibias.n276 161.3
R14759 commonsourceibias.n292 commonsourceibias.n291 161.3
R14760 commonsourceibias.n290 commonsourceibias.n289 161.3
R14761 commonsourceibias.n288 commonsourceibias.n278 161.3
R14762 commonsourceibias.n287 commonsourceibias.n286 161.3
R14763 commonsourceibias.n285 commonsourceibias.n284 161.3
R14764 commonsourceibias.n283 commonsourceibias.n280 161.3
R14765 commonsourceibias.n377 commonsourceibias.n273 161.3
R14766 commonsourceibias.n401 commonsourceibias.n266 161.3
R14767 commonsourceibias.n400 commonsourceibias.n399 161.3
R14768 commonsourceibias.n398 commonsourceibias.n397 161.3
R14769 commonsourceibias.n396 commonsourceibias.n268 161.3
R14770 commonsourceibias.n394 commonsourceibias.n393 161.3
R14771 commonsourceibias.n392 commonsourceibias.n269 161.3
R14772 commonsourceibias.n391 commonsourceibias.n390 161.3
R14773 commonsourceibias.n388 commonsourceibias.n270 161.3
R14774 commonsourceibias.n387 commonsourceibias.n386 161.3
R14775 commonsourceibias.n385 commonsourceibias.n271 161.3
R14776 commonsourceibias.n384 commonsourceibias.n383 161.3
R14777 commonsourceibias.n381 commonsourceibias.n272 161.3
R14778 commonsourceibias.n379 commonsourceibias.n378 161.3
R14779 commonsourceibias.n528 commonsourceibias.n468 161.3
R14780 commonsourceibias.n527 commonsourceibias.n526 161.3
R14781 commonsourceibias.n525 commonsourceibias.n524 161.3
R14782 commonsourceibias.n523 commonsourceibias.n470 161.3
R14783 commonsourceibias.n521 commonsourceibias.n520 161.3
R14784 commonsourceibias.n519 commonsourceibias.n471 161.3
R14785 commonsourceibias.n518 commonsourceibias.n517 161.3
R14786 commonsourceibias.n515 commonsourceibias.n472 161.3
R14787 commonsourceibias.n514 commonsourceibias.n513 161.3
R14788 commonsourceibias.n512 commonsourceibias.n473 161.3
R14789 commonsourceibias.n511 commonsourceibias.n510 161.3
R14790 commonsourceibias.n508 commonsourceibias.n474 161.3
R14791 commonsourceibias.n506 commonsourceibias.n505 161.3
R14792 commonsourceibias.n504 commonsourceibias.n475 161.3
R14793 commonsourceibias.n503 commonsourceibias.n502 161.3
R14794 commonsourceibias.n500 commonsourceibias.n476 161.3
R14795 commonsourceibias.n499 commonsourceibias.n498 161.3
R14796 commonsourceibias.n497 commonsourceibias.n496 161.3
R14797 commonsourceibias.n495 commonsourceibias.n478 161.3
R14798 commonsourceibias.n494 commonsourceibias.n493 161.3
R14799 commonsourceibias.n492 commonsourceibias.n491 161.3
R14800 commonsourceibias.n490 commonsourceibias.n480 161.3
R14801 commonsourceibias.n489 commonsourceibias.n488 161.3
R14802 commonsourceibias.n487 commonsourceibias.n486 161.3
R14803 commonsourceibias.n485 commonsourceibias.n482 161.3
R14804 commonsourceibias.n464 commonsourceibias.n404 161.3
R14805 commonsourceibias.n463 commonsourceibias.n462 161.3
R14806 commonsourceibias.n461 commonsourceibias.n460 161.3
R14807 commonsourceibias.n459 commonsourceibias.n406 161.3
R14808 commonsourceibias.n457 commonsourceibias.n456 161.3
R14809 commonsourceibias.n455 commonsourceibias.n407 161.3
R14810 commonsourceibias.n454 commonsourceibias.n453 161.3
R14811 commonsourceibias.n451 commonsourceibias.n408 161.3
R14812 commonsourceibias.n450 commonsourceibias.n449 161.3
R14813 commonsourceibias.n448 commonsourceibias.n409 161.3
R14814 commonsourceibias.n447 commonsourceibias.n446 161.3
R14815 commonsourceibias.n444 commonsourceibias.n410 161.3
R14816 commonsourceibias.n442 commonsourceibias.n441 161.3
R14817 commonsourceibias.n440 commonsourceibias.n411 161.3
R14818 commonsourceibias.n439 commonsourceibias.n438 161.3
R14819 commonsourceibias.n436 commonsourceibias.n412 161.3
R14820 commonsourceibias.n435 commonsourceibias.n434 161.3
R14821 commonsourceibias.n433 commonsourceibias.n432 161.3
R14822 commonsourceibias.n431 commonsourceibias.n414 161.3
R14823 commonsourceibias.n430 commonsourceibias.n429 161.3
R14824 commonsourceibias.n428 commonsourceibias.n427 161.3
R14825 commonsourceibias.n426 commonsourceibias.n416 161.3
R14826 commonsourceibias.n425 commonsourceibias.n424 161.3
R14827 commonsourceibias.n423 commonsourceibias.n422 161.3
R14828 commonsourceibias.n421 commonsourceibias.n418 161.3
R14829 commonsourceibias.n80 commonsourceibias.n78 81.5057
R14830 commonsourceibias.n304 commonsourceibias.n302 81.5057
R14831 commonsourceibias.n80 commonsourceibias.n79 80.9324
R14832 commonsourceibias.n82 commonsourceibias.n81 80.9324
R14833 commonsourceibias.n77 commonsourceibias.n76 80.9324
R14834 commonsourceibias.n75 commonsourceibias.n74 80.9324
R14835 commonsourceibias.n73 commonsourceibias.n72 80.9324
R14836 commonsourceibias.n371 commonsourceibias.n370 80.9324
R14837 commonsourceibias.n373 commonsourceibias.n372 80.9324
R14838 commonsourceibias.n375 commonsourceibias.n374 80.9324
R14839 commonsourceibias.n306 commonsourceibias.n305 80.9324
R14840 commonsourceibias.n304 commonsourceibias.n303 80.9324
R14841 commonsourceibias.n71 commonsourceibias.n70 80.6037
R14842 commonsourceibias.n137 commonsourceibias.n136 80.6037
R14843 commonsourceibias.n264 commonsourceibias.n263 80.6037
R14844 commonsourceibias.n200 commonsourceibias.n199 80.6037
R14845 commonsourceibias.n369 commonsourceibias.n368 80.6037
R14846 commonsourceibias.n403 commonsourceibias.n402 80.6037
R14847 commonsourceibias.n530 commonsourceibias.n529 80.6037
R14848 commonsourceibias.n466 commonsourceibias.n465 80.6037
R14849 commonsourceibias.n65 commonsourceibias.n64 56.5617
R14850 commonsourceibias.n51 commonsourceibias.n50 56.5617
R14851 commonsourceibias.n42 commonsourceibias.n41 56.5617
R14852 commonsourceibias.n28 commonsourceibias.n27 56.5617
R14853 commonsourceibias.n131 commonsourceibias.n130 56.5617
R14854 commonsourceibias.n117 commonsourceibias.n116 56.5617
R14855 commonsourceibias.n108 commonsourceibias.n107 56.5617
R14856 commonsourceibias.n94 commonsourceibias.n93 56.5617
R14857 commonsourceibias.n221 commonsourceibias.n220 56.5617
R14858 commonsourceibias.n235 commonsourceibias.n234 56.5617
R14859 commonsourceibias.n244 commonsourceibias.n243 56.5617
R14860 commonsourceibias.n258 commonsourceibias.n257 56.5617
R14861 commonsourceibias.n194 commonsourceibias.n193 56.5617
R14862 commonsourceibias.n180 commonsourceibias.n179 56.5617
R14863 commonsourceibias.n171 commonsourceibias.n170 56.5617
R14864 commonsourceibias.n157 commonsourceibias.n156 56.5617
R14865 commonsourceibias.n325 commonsourceibias.n324 56.5617
R14866 commonsourceibias.n339 commonsourceibias.n338 56.5617
R14867 commonsourceibias.n349 commonsourceibias.n347 56.5617
R14868 commonsourceibias.n363 commonsourceibias.n362 56.5617
R14869 commonsourceibias.n397 commonsourceibias.n396 56.5617
R14870 commonsourceibias.n383 commonsourceibias.n381 56.5617
R14871 commonsourceibias.n284 commonsourceibias.n283 56.5617
R14872 commonsourceibias.n298 commonsourceibias.n297 56.5617
R14873 commonsourceibias.n486 commonsourceibias.n485 56.5617
R14874 commonsourceibias.n500 commonsourceibias.n499 56.5617
R14875 commonsourceibias.n510 commonsourceibias.n508 56.5617
R14876 commonsourceibias.n524 commonsourceibias.n523 56.5617
R14877 commonsourceibias.n422 commonsourceibias.n421 56.5617
R14878 commonsourceibias.n436 commonsourceibias.n435 56.5617
R14879 commonsourceibias.n446 commonsourceibias.n444 56.5617
R14880 commonsourceibias.n460 commonsourceibias.n459 56.5617
R14881 commonsourceibias.n56 commonsourceibias.n55 56.0773
R14882 commonsourceibias.n37 commonsourceibias.n36 56.0773
R14883 commonsourceibias.n122 commonsourceibias.n121 56.0773
R14884 commonsourceibias.n103 commonsourceibias.n102 56.0773
R14885 commonsourceibias.n230 commonsourceibias.n229 56.0773
R14886 commonsourceibias.n249 commonsourceibias.n248 56.0773
R14887 commonsourceibias.n185 commonsourceibias.n184 56.0773
R14888 commonsourceibias.n166 commonsourceibias.n165 56.0773
R14889 commonsourceibias.n334 commonsourceibias.n333 56.0773
R14890 commonsourceibias.n354 commonsourceibias.n353 56.0773
R14891 commonsourceibias.n388 commonsourceibias.n387 56.0773
R14892 commonsourceibias.n293 commonsourceibias.n292 56.0773
R14893 commonsourceibias.n495 commonsourceibias.n494 56.0773
R14894 commonsourceibias.n515 commonsourceibias.n514 56.0773
R14895 commonsourceibias.n431 commonsourceibias.n430 56.0773
R14896 commonsourceibias.n451 commonsourceibias.n450 56.0773
R14897 commonsourceibias.n70 commonsourceibias.n69 46.0096
R14898 commonsourceibias.n136 commonsourceibias.n135 46.0096
R14899 commonsourceibias.n263 commonsourceibias.n262 46.0096
R14900 commonsourceibias.n199 commonsourceibias.n198 46.0096
R14901 commonsourceibias.n368 commonsourceibias.n367 46.0096
R14902 commonsourceibias.n402 commonsourceibias.n401 46.0096
R14903 commonsourceibias.n529 commonsourceibias.n528 46.0096
R14904 commonsourceibias.n465 commonsourceibias.n464 46.0096
R14905 commonsourceibias.n58 commonsourceibias.n12 41.5458
R14906 commonsourceibias.n33 commonsourceibias.n32 41.5458
R14907 commonsourceibias.n124 commonsourceibias.n3 41.5458
R14908 commonsourceibias.n99 commonsourceibias.n98 41.5458
R14909 commonsourceibias.n226 commonsourceibias.n225 41.5458
R14910 commonsourceibias.n251 commonsourceibias.n205 41.5458
R14911 commonsourceibias.n187 commonsourceibias.n141 41.5458
R14912 commonsourceibias.n162 commonsourceibias.n161 41.5458
R14913 commonsourceibias.n330 commonsourceibias.n329 41.5458
R14914 commonsourceibias.n356 commonsourceibias.n310 41.5458
R14915 commonsourceibias.n390 commonsourceibias.n269 41.5458
R14916 commonsourceibias.n289 commonsourceibias.n288 41.5458
R14917 commonsourceibias.n491 commonsourceibias.n490 41.5458
R14918 commonsourceibias.n517 commonsourceibias.n471 41.5458
R14919 commonsourceibias.n427 commonsourceibias.n426 41.5458
R14920 commonsourceibias.n453 commonsourceibias.n407 41.5458
R14921 commonsourceibias.n48 commonsourceibias.n17 40.577
R14922 commonsourceibias.n44 commonsourceibias.n17 40.577
R14923 commonsourceibias.n114 commonsourceibias.n8 40.577
R14924 commonsourceibias.n110 commonsourceibias.n8 40.577
R14925 commonsourceibias.n237 commonsourceibias.n210 40.577
R14926 commonsourceibias.n241 commonsourceibias.n210 40.577
R14927 commonsourceibias.n177 commonsourceibias.n146 40.577
R14928 commonsourceibias.n173 commonsourceibias.n146 40.577
R14929 commonsourceibias.n341 commonsourceibias.n314 40.577
R14930 commonsourceibias.n345 commonsourceibias.n314 40.577
R14931 commonsourceibias.n379 commonsourceibias.n273 40.577
R14932 commonsourceibias.n300 commonsourceibias.n273 40.577
R14933 commonsourceibias.n502 commonsourceibias.n475 40.577
R14934 commonsourceibias.n506 commonsourceibias.n475 40.577
R14935 commonsourceibias.n438 commonsourceibias.n411 40.577
R14936 commonsourceibias.n442 commonsourceibias.n411 40.577
R14937 commonsourceibias.n62 commonsourceibias.n12 39.6083
R14938 commonsourceibias.n32 commonsourceibias.n31 39.6083
R14939 commonsourceibias.n128 commonsourceibias.n3 39.6083
R14940 commonsourceibias.n98 commonsourceibias.n97 39.6083
R14941 commonsourceibias.n225 commonsourceibias.n224 39.6083
R14942 commonsourceibias.n255 commonsourceibias.n205 39.6083
R14943 commonsourceibias.n191 commonsourceibias.n141 39.6083
R14944 commonsourceibias.n161 commonsourceibias.n160 39.6083
R14945 commonsourceibias.n329 commonsourceibias.n328 39.6083
R14946 commonsourceibias.n360 commonsourceibias.n310 39.6083
R14947 commonsourceibias.n394 commonsourceibias.n269 39.6083
R14948 commonsourceibias.n288 commonsourceibias.n287 39.6083
R14949 commonsourceibias.n490 commonsourceibias.n489 39.6083
R14950 commonsourceibias.n521 commonsourceibias.n471 39.6083
R14951 commonsourceibias.n426 commonsourceibias.n425 39.6083
R14952 commonsourceibias.n457 commonsourceibias.n407 39.6083
R14953 commonsourceibias.n26 commonsourceibias.n25 33.0515
R14954 commonsourceibias.n92 commonsourceibias.n91 33.0515
R14955 commonsourceibias.n155 commonsourceibias.n154 33.0515
R14956 commonsourceibias.n219 commonsourceibias.n218 33.0515
R14957 commonsourceibias.n323 commonsourceibias.n322 33.0515
R14958 commonsourceibias.n282 commonsourceibias.n281 33.0515
R14959 commonsourceibias.n484 commonsourceibias.n483 33.0515
R14960 commonsourceibias.n420 commonsourceibias.n419 33.0515
R14961 commonsourceibias.n25 commonsourceibias.n24 28.5514
R14962 commonsourceibias.n91 commonsourceibias.n90 28.5514
R14963 commonsourceibias.n218 commonsourceibias.n217 28.5514
R14964 commonsourceibias.n154 commonsourceibias.n153 28.5514
R14965 commonsourceibias.n322 commonsourceibias.n321 28.5514
R14966 commonsourceibias.n281 commonsourceibias.n280 28.5514
R14967 commonsourceibias.n483 commonsourceibias.n482 28.5514
R14968 commonsourceibias.n419 commonsourceibias.n418 28.5514
R14969 commonsourceibias.n69 commonsourceibias.n68 26.0455
R14970 commonsourceibias.n135 commonsourceibias.n134 26.0455
R14971 commonsourceibias.n262 commonsourceibias.n261 26.0455
R14972 commonsourceibias.n198 commonsourceibias.n197 26.0455
R14973 commonsourceibias.n367 commonsourceibias.n366 26.0455
R14974 commonsourceibias.n401 commonsourceibias.n400 26.0455
R14975 commonsourceibias.n528 commonsourceibias.n527 26.0455
R14976 commonsourceibias.n464 commonsourceibias.n463 26.0455
R14977 commonsourceibias.n55 commonsourceibias.n14 25.0767
R14978 commonsourceibias.n38 commonsourceibias.n37 25.0767
R14979 commonsourceibias.n121 commonsourceibias.n5 25.0767
R14980 commonsourceibias.n104 commonsourceibias.n103 25.0767
R14981 commonsourceibias.n231 commonsourceibias.n230 25.0767
R14982 commonsourceibias.n248 commonsourceibias.n207 25.0767
R14983 commonsourceibias.n184 commonsourceibias.n143 25.0767
R14984 commonsourceibias.n167 commonsourceibias.n166 25.0767
R14985 commonsourceibias.n335 commonsourceibias.n334 25.0767
R14986 commonsourceibias.n353 commonsourceibias.n312 25.0767
R14987 commonsourceibias.n387 commonsourceibias.n271 25.0767
R14988 commonsourceibias.n294 commonsourceibias.n293 25.0767
R14989 commonsourceibias.n496 commonsourceibias.n495 25.0767
R14990 commonsourceibias.n514 commonsourceibias.n473 25.0767
R14991 commonsourceibias.n432 commonsourceibias.n431 25.0767
R14992 commonsourceibias.n450 commonsourceibias.n409 25.0767
R14993 commonsourceibias.n51 commonsourceibias.n16 24.3464
R14994 commonsourceibias.n41 commonsourceibias.n19 24.3464
R14995 commonsourceibias.n117 commonsourceibias.n7 24.3464
R14996 commonsourceibias.n107 commonsourceibias.n85 24.3464
R14997 commonsourceibias.n234 commonsourceibias.n212 24.3464
R14998 commonsourceibias.n244 commonsourceibias.n209 24.3464
R14999 commonsourceibias.n180 commonsourceibias.n145 24.3464
R15000 commonsourceibias.n170 commonsourceibias.n148 24.3464
R15001 commonsourceibias.n338 commonsourceibias.n316 24.3464
R15002 commonsourceibias.n349 commonsourceibias.n348 24.3464
R15003 commonsourceibias.n383 commonsourceibias.n382 24.3464
R15004 commonsourceibias.n297 commonsourceibias.n275 24.3464
R15005 commonsourceibias.n499 commonsourceibias.n477 24.3464
R15006 commonsourceibias.n510 commonsourceibias.n509 24.3464
R15007 commonsourceibias.n435 commonsourceibias.n413 24.3464
R15008 commonsourceibias.n446 commonsourceibias.n445 24.3464
R15009 commonsourceibias.n65 commonsourceibias.n10 23.8546
R15010 commonsourceibias.n27 commonsourceibias.n26 23.8546
R15011 commonsourceibias.n131 commonsourceibias.n1 23.8546
R15012 commonsourceibias.n93 commonsourceibias.n92 23.8546
R15013 commonsourceibias.n220 commonsourceibias.n219 23.8546
R15014 commonsourceibias.n258 commonsourceibias.n203 23.8546
R15015 commonsourceibias.n194 commonsourceibias.n139 23.8546
R15016 commonsourceibias.n156 commonsourceibias.n155 23.8546
R15017 commonsourceibias.n324 commonsourceibias.n323 23.8546
R15018 commonsourceibias.n363 commonsourceibias.n308 23.8546
R15019 commonsourceibias.n397 commonsourceibias.n267 23.8546
R15020 commonsourceibias.n283 commonsourceibias.n282 23.8546
R15021 commonsourceibias.n485 commonsourceibias.n484 23.8546
R15022 commonsourceibias.n524 commonsourceibias.n469 23.8546
R15023 commonsourceibias.n421 commonsourceibias.n420 23.8546
R15024 commonsourceibias.n460 commonsourceibias.n405 23.8546
R15025 commonsourceibias.n64 commonsourceibias.n63 16.9689
R15026 commonsourceibias.n28 commonsourceibias.n23 16.9689
R15027 commonsourceibias.n130 commonsourceibias.n129 16.9689
R15028 commonsourceibias.n94 commonsourceibias.n89 16.9689
R15029 commonsourceibias.n221 commonsourceibias.n216 16.9689
R15030 commonsourceibias.n257 commonsourceibias.n256 16.9689
R15031 commonsourceibias.n193 commonsourceibias.n192 16.9689
R15032 commonsourceibias.n157 commonsourceibias.n152 16.9689
R15033 commonsourceibias.n325 commonsourceibias.n320 16.9689
R15034 commonsourceibias.n362 commonsourceibias.n361 16.9689
R15035 commonsourceibias.n396 commonsourceibias.n395 16.9689
R15036 commonsourceibias.n284 commonsourceibias.n279 16.9689
R15037 commonsourceibias.n486 commonsourceibias.n481 16.9689
R15038 commonsourceibias.n523 commonsourceibias.n522 16.9689
R15039 commonsourceibias.n422 commonsourceibias.n417 16.9689
R15040 commonsourceibias.n459 commonsourceibias.n458 16.9689
R15041 commonsourceibias.n50 commonsourceibias.n49 16.477
R15042 commonsourceibias.n43 commonsourceibias.n42 16.477
R15043 commonsourceibias.n116 commonsourceibias.n115 16.477
R15044 commonsourceibias.n109 commonsourceibias.n108 16.477
R15045 commonsourceibias.n236 commonsourceibias.n235 16.477
R15046 commonsourceibias.n243 commonsourceibias.n242 16.477
R15047 commonsourceibias.n179 commonsourceibias.n178 16.477
R15048 commonsourceibias.n172 commonsourceibias.n171 16.477
R15049 commonsourceibias.n340 commonsourceibias.n339 16.477
R15050 commonsourceibias.n347 commonsourceibias.n346 16.477
R15051 commonsourceibias.n381 commonsourceibias.n380 16.477
R15052 commonsourceibias.n299 commonsourceibias.n298 16.477
R15053 commonsourceibias.n501 commonsourceibias.n500 16.477
R15054 commonsourceibias.n508 commonsourceibias.n507 16.477
R15055 commonsourceibias.n437 commonsourceibias.n436 16.477
R15056 commonsourceibias.n444 commonsourceibias.n443 16.477
R15057 commonsourceibias.n57 commonsourceibias.n56 15.9852
R15058 commonsourceibias.n36 commonsourceibias.n21 15.9852
R15059 commonsourceibias.n123 commonsourceibias.n122 15.9852
R15060 commonsourceibias.n102 commonsourceibias.n87 15.9852
R15061 commonsourceibias.n229 commonsourceibias.n214 15.9852
R15062 commonsourceibias.n250 commonsourceibias.n249 15.9852
R15063 commonsourceibias.n186 commonsourceibias.n185 15.9852
R15064 commonsourceibias.n165 commonsourceibias.n150 15.9852
R15065 commonsourceibias.n333 commonsourceibias.n318 15.9852
R15066 commonsourceibias.n355 commonsourceibias.n354 15.9852
R15067 commonsourceibias.n389 commonsourceibias.n388 15.9852
R15068 commonsourceibias.n292 commonsourceibias.n277 15.9852
R15069 commonsourceibias.n494 commonsourceibias.n479 15.9852
R15070 commonsourceibias.n516 commonsourceibias.n515 15.9852
R15071 commonsourceibias.n430 commonsourceibias.n415 15.9852
R15072 commonsourceibias.n452 commonsourceibias.n451 15.9852
R15073 commonsourceibias.n73 commonsourceibias.n71 13.2057
R15074 commonsourceibias.n371 commonsourceibias.n369 13.2057
R15075 commonsourceibias.n532 commonsourceibias.n265 10.122
R15076 commonsourceibias.n112 commonsourceibias.n83 9.50363
R15077 commonsourceibias.n377 commonsourceibias.n376 9.50363
R15078 commonsourceibias.n201 commonsourceibias.n137 8.7339
R15079 commonsourceibias.n467 commonsourceibias.n403 8.7339
R15080 commonsourceibias.n58 commonsourceibias.n57 8.60764
R15081 commonsourceibias.n33 commonsourceibias.n21 8.60764
R15082 commonsourceibias.n124 commonsourceibias.n123 8.60764
R15083 commonsourceibias.n99 commonsourceibias.n87 8.60764
R15084 commonsourceibias.n226 commonsourceibias.n214 8.60764
R15085 commonsourceibias.n251 commonsourceibias.n250 8.60764
R15086 commonsourceibias.n187 commonsourceibias.n186 8.60764
R15087 commonsourceibias.n162 commonsourceibias.n150 8.60764
R15088 commonsourceibias.n330 commonsourceibias.n318 8.60764
R15089 commonsourceibias.n356 commonsourceibias.n355 8.60764
R15090 commonsourceibias.n390 commonsourceibias.n389 8.60764
R15091 commonsourceibias.n289 commonsourceibias.n277 8.60764
R15092 commonsourceibias.n491 commonsourceibias.n479 8.60764
R15093 commonsourceibias.n517 commonsourceibias.n516 8.60764
R15094 commonsourceibias.n427 commonsourceibias.n415 8.60764
R15095 commonsourceibias.n453 commonsourceibias.n452 8.60764
R15096 commonsourceibias.n532 commonsourceibias.n531 8.46921
R15097 commonsourceibias.n49 commonsourceibias.n48 8.11581
R15098 commonsourceibias.n44 commonsourceibias.n43 8.11581
R15099 commonsourceibias.n115 commonsourceibias.n114 8.11581
R15100 commonsourceibias.n110 commonsourceibias.n109 8.11581
R15101 commonsourceibias.n237 commonsourceibias.n236 8.11581
R15102 commonsourceibias.n242 commonsourceibias.n241 8.11581
R15103 commonsourceibias.n178 commonsourceibias.n177 8.11581
R15104 commonsourceibias.n173 commonsourceibias.n172 8.11581
R15105 commonsourceibias.n341 commonsourceibias.n340 8.11581
R15106 commonsourceibias.n346 commonsourceibias.n345 8.11581
R15107 commonsourceibias.n380 commonsourceibias.n379 8.11581
R15108 commonsourceibias.n300 commonsourceibias.n299 8.11581
R15109 commonsourceibias.n502 commonsourceibias.n501 8.11581
R15110 commonsourceibias.n507 commonsourceibias.n506 8.11581
R15111 commonsourceibias.n438 commonsourceibias.n437 8.11581
R15112 commonsourceibias.n443 commonsourceibias.n442 8.11581
R15113 commonsourceibias.n63 commonsourceibias.n62 7.62397
R15114 commonsourceibias.n31 commonsourceibias.n23 7.62397
R15115 commonsourceibias.n129 commonsourceibias.n128 7.62397
R15116 commonsourceibias.n97 commonsourceibias.n89 7.62397
R15117 commonsourceibias.n224 commonsourceibias.n216 7.62397
R15118 commonsourceibias.n256 commonsourceibias.n255 7.62397
R15119 commonsourceibias.n192 commonsourceibias.n191 7.62397
R15120 commonsourceibias.n160 commonsourceibias.n152 7.62397
R15121 commonsourceibias.n328 commonsourceibias.n320 7.62397
R15122 commonsourceibias.n361 commonsourceibias.n360 7.62397
R15123 commonsourceibias.n395 commonsourceibias.n394 7.62397
R15124 commonsourceibias.n287 commonsourceibias.n279 7.62397
R15125 commonsourceibias.n489 commonsourceibias.n481 7.62397
R15126 commonsourceibias.n522 commonsourceibias.n521 7.62397
R15127 commonsourceibias.n425 commonsourceibias.n417 7.62397
R15128 commonsourceibias.n458 commonsourceibias.n457 7.62397
R15129 commonsourceibias.n265 commonsourceibias.n264 5.00473
R15130 commonsourceibias.n201 commonsourceibias.n200 5.00473
R15131 commonsourceibias.n531 commonsourceibias.n530 5.00473
R15132 commonsourceibias.n467 commonsourceibias.n466 5.00473
R15133 commonsourceibias commonsourceibias.n532 4.08303
R15134 commonsourceibias.n265 commonsourceibias.n201 3.72967
R15135 commonsourceibias.n531 commonsourceibias.n467 3.72967
R15136 commonsourceibias.n78 commonsourceibias.t17 2.82907
R15137 commonsourceibias.n78 commonsourceibias.t23 2.82907
R15138 commonsourceibias.n79 commonsourceibias.t11 2.82907
R15139 commonsourceibias.n79 commonsourceibias.t35 2.82907
R15140 commonsourceibias.n81 commonsourceibias.t21 2.82907
R15141 commonsourceibias.n81 commonsourceibias.t3 2.82907
R15142 commonsourceibias.n76 commonsourceibias.t45 2.82907
R15143 commonsourceibias.n76 commonsourceibias.t13 2.82907
R15144 commonsourceibias.n74 commonsourceibias.t1 2.82907
R15145 commonsourceibias.n74 commonsourceibias.t7 2.82907
R15146 commonsourceibias.n72 commonsourceibias.t9 2.82907
R15147 commonsourceibias.n72 commonsourceibias.t39 2.82907
R15148 commonsourceibias.n370 commonsourceibias.t47 2.82907
R15149 commonsourceibias.n370 commonsourceibias.t27 2.82907
R15150 commonsourceibias.n372 commonsourceibias.t25 2.82907
R15151 commonsourceibias.n372 commonsourceibias.t15 2.82907
R15152 commonsourceibias.n374 commonsourceibias.t31 2.82907
R15153 commonsourceibias.n374 commonsourceibias.t5 2.82907
R15154 commonsourceibias.n305 commonsourceibias.t19 2.82907
R15155 commonsourceibias.n305 commonsourceibias.t37 2.82907
R15156 commonsourceibias.n303 commonsourceibias.t43 2.82907
R15157 commonsourceibias.n303 commonsourceibias.t29 2.82907
R15158 commonsourceibias.n302 commonsourceibias.t41 2.82907
R15159 commonsourceibias.n302 commonsourceibias.t33 2.82907
R15160 commonsourceibias.n68 commonsourceibias.n10 0.738255
R15161 commonsourceibias.n134 commonsourceibias.n1 0.738255
R15162 commonsourceibias.n261 commonsourceibias.n203 0.738255
R15163 commonsourceibias.n197 commonsourceibias.n139 0.738255
R15164 commonsourceibias.n366 commonsourceibias.n308 0.738255
R15165 commonsourceibias.n400 commonsourceibias.n267 0.738255
R15166 commonsourceibias.n527 commonsourceibias.n469 0.738255
R15167 commonsourceibias.n463 commonsourceibias.n405 0.738255
R15168 commonsourceibias.n75 commonsourceibias.n73 0.573776
R15169 commonsourceibias.n77 commonsourceibias.n75 0.573776
R15170 commonsourceibias.n82 commonsourceibias.n80 0.573776
R15171 commonsourceibias.n306 commonsourceibias.n304 0.573776
R15172 commonsourceibias.n375 commonsourceibias.n373 0.573776
R15173 commonsourceibias.n373 commonsourceibias.n371 0.573776
R15174 commonsourceibias.n83 commonsourceibias.n77 0.287138
R15175 commonsourceibias.n83 commonsourceibias.n82 0.287138
R15176 commonsourceibias.n376 commonsourceibias.n306 0.287138
R15177 commonsourceibias.n376 commonsourceibias.n375 0.287138
R15178 commonsourceibias.n71 commonsourceibias.n9 0.285035
R15179 commonsourceibias.n137 commonsourceibias.n0 0.285035
R15180 commonsourceibias.n264 commonsourceibias.n202 0.285035
R15181 commonsourceibias.n200 commonsourceibias.n138 0.285035
R15182 commonsourceibias.n369 commonsourceibias.n307 0.285035
R15183 commonsourceibias.n403 commonsourceibias.n266 0.285035
R15184 commonsourceibias.n530 commonsourceibias.n468 0.285035
R15185 commonsourceibias.n466 commonsourceibias.n404 0.285035
R15186 commonsourceibias.n16 commonsourceibias.n14 0.246418
R15187 commonsourceibias.n38 commonsourceibias.n19 0.246418
R15188 commonsourceibias.n7 commonsourceibias.n5 0.246418
R15189 commonsourceibias.n104 commonsourceibias.n85 0.246418
R15190 commonsourceibias.n231 commonsourceibias.n212 0.246418
R15191 commonsourceibias.n209 commonsourceibias.n207 0.246418
R15192 commonsourceibias.n145 commonsourceibias.n143 0.246418
R15193 commonsourceibias.n167 commonsourceibias.n148 0.246418
R15194 commonsourceibias.n335 commonsourceibias.n316 0.246418
R15195 commonsourceibias.n348 commonsourceibias.n312 0.246418
R15196 commonsourceibias.n382 commonsourceibias.n271 0.246418
R15197 commonsourceibias.n294 commonsourceibias.n275 0.246418
R15198 commonsourceibias.n496 commonsourceibias.n477 0.246418
R15199 commonsourceibias.n509 commonsourceibias.n473 0.246418
R15200 commonsourceibias.n432 commonsourceibias.n413 0.246418
R15201 commonsourceibias.n445 commonsourceibias.n409 0.246418
R15202 commonsourceibias.n67 commonsourceibias.n9 0.189894
R15203 commonsourceibias.n67 commonsourceibias.n66 0.189894
R15204 commonsourceibias.n66 commonsourceibias.n11 0.189894
R15205 commonsourceibias.n61 commonsourceibias.n11 0.189894
R15206 commonsourceibias.n61 commonsourceibias.n60 0.189894
R15207 commonsourceibias.n60 commonsourceibias.n59 0.189894
R15208 commonsourceibias.n59 commonsourceibias.n13 0.189894
R15209 commonsourceibias.n54 commonsourceibias.n13 0.189894
R15210 commonsourceibias.n54 commonsourceibias.n53 0.189894
R15211 commonsourceibias.n53 commonsourceibias.n52 0.189894
R15212 commonsourceibias.n52 commonsourceibias.n15 0.189894
R15213 commonsourceibias.n47 commonsourceibias.n15 0.189894
R15214 commonsourceibias.n47 commonsourceibias.n46 0.189894
R15215 commonsourceibias.n46 commonsourceibias.n45 0.189894
R15216 commonsourceibias.n45 commonsourceibias.n18 0.189894
R15217 commonsourceibias.n40 commonsourceibias.n18 0.189894
R15218 commonsourceibias.n40 commonsourceibias.n39 0.189894
R15219 commonsourceibias.n39 commonsourceibias.n20 0.189894
R15220 commonsourceibias.n35 commonsourceibias.n20 0.189894
R15221 commonsourceibias.n35 commonsourceibias.n34 0.189894
R15222 commonsourceibias.n34 commonsourceibias.n22 0.189894
R15223 commonsourceibias.n30 commonsourceibias.n22 0.189894
R15224 commonsourceibias.n30 commonsourceibias.n29 0.189894
R15225 commonsourceibias.n29 commonsourceibias.n24 0.189894
R15226 commonsourceibias.n111 commonsourceibias.n84 0.189894
R15227 commonsourceibias.n106 commonsourceibias.n84 0.189894
R15228 commonsourceibias.n106 commonsourceibias.n105 0.189894
R15229 commonsourceibias.n105 commonsourceibias.n86 0.189894
R15230 commonsourceibias.n101 commonsourceibias.n86 0.189894
R15231 commonsourceibias.n101 commonsourceibias.n100 0.189894
R15232 commonsourceibias.n100 commonsourceibias.n88 0.189894
R15233 commonsourceibias.n96 commonsourceibias.n88 0.189894
R15234 commonsourceibias.n96 commonsourceibias.n95 0.189894
R15235 commonsourceibias.n95 commonsourceibias.n90 0.189894
R15236 commonsourceibias.n133 commonsourceibias.n0 0.189894
R15237 commonsourceibias.n133 commonsourceibias.n132 0.189894
R15238 commonsourceibias.n132 commonsourceibias.n2 0.189894
R15239 commonsourceibias.n127 commonsourceibias.n2 0.189894
R15240 commonsourceibias.n127 commonsourceibias.n126 0.189894
R15241 commonsourceibias.n126 commonsourceibias.n125 0.189894
R15242 commonsourceibias.n125 commonsourceibias.n4 0.189894
R15243 commonsourceibias.n120 commonsourceibias.n4 0.189894
R15244 commonsourceibias.n120 commonsourceibias.n119 0.189894
R15245 commonsourceibias.n119 commonsourceibias.n118 0.189894
R15246 commonsourceibias.n118 commonsourceibias.n6 0.189894
R15247 commonsourceibias.n113 commonsourceibias.n6 0.189894
R15248 commonsourceibias.n260 commonsourceibias.n202 0.189894
R15249 commonsourceibias.n260 commonsourceibias.n259 0.189894
R15250 commonsourceibias.n259 commonsourceibias.n204 0.189894
R15251 commonsourceibias.n254 commonsourceibias.n204 0.189894
R15252 commonsourceibias.n254 commonsourceibias.n253 0.189894
R15253 commonsourceibias.n253 commonsourceibias.n252 0.189894
R15254 commonsourceibias.n252 commonsourceibias.n206 0.189894
R15255 commonsourceibias.n247 commonsourceibias.n206 0.189894
R15256 commonsourceibias.n247 commonsourceibias.n246 0.189894
R15257 commonsourceibias.n246 commonsourceibias.n245 0.189894
R15258 commonsourceibias.n245 commonsourceibias.n208 0.189894
R15259 commonsourceibias.n240 commonsourceibias.n208 0.189894
R15260 commonsourceibias.n240 commonsourceibias.n239 0.189894
R15261 commonsourceibias.n239 commonsourceibias.n238 0.189894
R15262 commonsourceibias.n238 commonsourceibias.n211 0.189894
R15263 commonsourceibias.n233 commonsourceibias.n211 0.189894
R15264 commonsourceibias.n233 commonsourceibias.n232 0.189894
R15265 commonsourceibias.n232 commonsourceibias.n213 0.189894
R15266 commonsourceibias.n228 commonsourceibias.n213 0.189894
R15267 commonsourceibias.n228 commonsourceibias.n227 0.189894
R15268 commonsourceibias.n227 commonsourceibias.n215 0.189894
R15269 commonsourceibias.n223 commonsourceibias.n215 0.189894
R15270 commonsourceibias.n223 commonsourceibias.n222 0.189894
R15271 commonsourceibias.n222 commonsourceibias.n217 0.189894
R15272 commonsourceibias.n196 commonsourceibias.n138 0.189894
R15273 commonsourceibias.n196 commonsourceibias.n195 0.189894
R15274 commonsourceibias.n195 commonsourceibias.n140 0.189894
R15275 commonsourceibias.n190 commonsourceibias.n140 0.189894
R15276 commonsourceibias.n190 commonsourceibias.n189 0.189894
R15277 commonsourceibias.n189 commonsourceibias.n188 0.189894
R15278 commonsourceibias.n188 commonsourceibias.n142 0.189894
R15279 commonsourceibias.n183 commonsourceibias.n142 0.189894
R15280 commonsourceibias.n183 commonsourceibias.n182 0.189894
R15281 commonsourceibias.n182 commonsourceibias.n181 0.189894
R15282 commonsourceibias.n181 commonsourceibias.n144 0.189894
R15283 commonsourceibias.n176 commonsourceibias.n144 0.189894
R15284 commonsourceibias.n176 commonsourceibias.n175 0.189894
R15285 commonsourceibias.n175 commonsourceibias.n174 0.189894
R15286 commonsourceibias.n174 commonsourceibias.n147 0.189894
R15287 commonsourceibias.n169 commonsourceibias.n147 0.189894
R15288 commonsourceibias.n169 commonsourceibias.n168 0.189894
R15289 commonsourceibias.n168 commonsourceibias.n149 0.189894
R15290 commonsourceibias.n164 commonsourceibias.n149 0.189894
R15291 commonsourceibias.n164 commonsourceibias.n163 0.189894
R15292 commonsourceibias.n163 commonsourceibias.n151 0.189894
R15293 commonsourceibias.n159 commonsourceibias.n151 0.189894
R15294 commonsourceibias.n159 commonsourceibias.n158 0.189894
R15295 commonsourceibias.n158 commonsourceibias.n153 0.189894
R15296 commonsourceibias.n326 commonsourceibias.n321 0.189894
R15297 commonsourceibias.n327 commonsourceibias.n326 0.189894
R15298 commonsourceibias.n327 commonsourceibias.n319 0.189894
R15299 commonsourceibias.n331 commonsourceibias.n319 0.189894
R15300 commonsourceibias.n332 commonsourceibias.n331 0.189894
R15301 commonsourceibias.n332 commonsourceibias.n317 0.189894
R15302 commonsourceibias.n336 commonsourceibias.n317 0.189894
R15303 commonsourceibias.n337 commonsourceibias.n336 0.189894
R15304 commonsourceibias.n337 commonsourceibias.n315 0.189894
R15305 commonsourceibias.n342 commonsourceibias.n315 0.189894
R15306 commonsourceibias.n343 commonsourceibias.n342 0.189894
R15307 commonsourceibias.n344 commonsourceibias.n343 0.189894
R15308 commonsourceibias.n344 commonsourceibias.n313 0.189894
R15309 commonsourceibias.n350 commonsourceibias.n313 0.189894
R15310 commonsourceibias.n351 commonsourceibias.n350 0.189894
R15311 commonsourceibias.n352 commonsourceibias.n351 0.189894
R15312 commonsourceibias.n352 commonsourceibias.n311 0.189894
R15313 commonsourceibias.n357 commonsourceibias.n311 0.189894
R15314 commonsourceibias.n358 commonsourceibias.n357 0.189894
R15315 commonsourceibias.n359 commonsourceibias.n358 0.189894
R15316 commonsourceibias.n359 commonsourceibias.n309 0.189894
R15317 commonsourceibias.n364 commonsourceibias.n309 0.189894
R15318 commonsourceibias.n365 commonsourceibias.n364 0.189894
R15319 commonsourceibias.n365 commonsourceibias.n307 0.189894
R15320 commonsourceibias.n285 commonsourceibias.n280 0.189894
R15321 commonsourceibias.n286 commonsourceibias.n285 0.189894
R15322 commonsourceibias.n286 commonsourceibias.n278 0.189894
R15323 commonsourceibias.n290 commonsourceibias.n278 0.189894
R15324 commonsourceibias.n291 commonsourceibias.n290 0.189894
R15325 commonsourceibias.n291 commonsourceibias.n276 0.189894
R15326 commonsourceibias.n295 commonsourceibias.n276 0.189894
R15327 commonsourceibias.n296 commonsourceibias.n295 0.189894
R15328 commonsourceibias.n296 commonsourceibias.n274 0.189894
R15329 commonsourceibias.n301 commonsourceibias.n274 0.189894
R15330 commonsourceibias.n378 commonsourceibias.n272 0.189894
R15331 commonsourceibias.n384 commonsourceibias.n272 0.189894
R15332 commonsourceibias.n385 commonsourceibias.n384 0.189894
R15333 commonsourceibias.n386 commonsourceibias.n385 0.189894
R15334 commonsourceibias.n386 commonsourceibias.n270 0.189894
R15335 commonsourceibias.n391 commonsourceibias.n270 0.189894
R15336 commonsourceibias.n392 commonsourceibias.n391 0.189894
R15337 commonsourceibias.n393 commonsourceibias.n392 0.189894
R15338 commonsourceibias.n393 commonsourceibias.n268 0.189894
R15339 commonsourceibias.n398 commonsourceibias.n268 0.189894
R15340 commonsourceibias.n399 commonsourceibias.n398 0.189894
R15341 commonsourceibias.n399 commonsourceibias.n266 0.189894
R15342 commonsourceibias.n487 commonsourceibias.n482 0.189894
R15343 commonsourceibias.n488 commonsourceibias.n487 0.189894
R15344 commonsourceibias.n488 commonsourceibias.n480 0.189894
R15345 commonsourceibias.n492 commonsourceibias.n480 0.189894
R15346 commonsourceibias.n493 commonsourceibias.n492 0.189894
R15347 commonsourceibias.n493 commonsourceibias.n478 0.189894
R15348 commonsourceibias.n497 commonsourceibias.n478 0.189894
R15349 commonsourceibias.n498 commonsourceibias.n497 0.189894
R15350 commonsourceibias.n498 commonsourceibias.n476 0.189894
R15351 commonsourceibias.n503 commonsourceibias.n476 0.189894
R15352 commonsourceibias.n504 commonsourceibias.n503 0.189894
R15353 commonsourceibias.n505 commonsourceibias.n504 0.189894
R15354 commonsourceibias.n505 commonsourceibias.n474 0.189894
R15355 commonsourceibias.n511 commonsourceibias.n474 0.189894
R15356 commonsourceibias.n512 commonsourceibias.n511 0.189894
R15357 commonsourceibias.n513 commonsourceibias.n512 0.189894
R15358 commonsourceibias.n513 commonsourceibias.n472 0.189894
R15359 commonsourceibias.n518 commonsourceibias.n472 0.189894
R15360 commonsourceibias.n519 commonsourceibias.n518 0.189894
R15361 commonsourceibias.n520 commonsourceibias.n519 0.189894
R15362 commonsourceibias.n520 commonsourceibias.n470 0.189894
R15363 commonsourceibias.n525 commonsourceibias.n470 0.189894
R15364 commonsourceibias.n526 commonsourceibias.n525 0.189894
R15365 commonsourceibias.n526 commonsourceibias.n468 0.189894
R15366 commonsourceibias.n423 commonsourceibias.n418 0.189894
R15367 commonsourceibias.n424 commonsourceibias.n423 0.189894
R15368 commonsourceibias.n424 commonsourceibias.n416 0.189894
R15369 commonsourceibias.n428 commonsourceibias.n416 0.189894
R15370 commonsourceibias.n429 commonsourceibias.n428 0.189894
R15371 commonsourceibias.n429 commonsourceibias.n414 0.189894
R15372 commonsourceibias.n433 commonsourceibias.n414 0.189894
R15373 commonsourceibias.n434 commonsourceibias.n433 0.189894
R15374 commonsourceibias.n434 commonsourceibias.n412 0.189894
R15375 commonsourceibias.n439 commonsourceibias.n412 0.189894
R15376 commonsourceibias.n440 commonsourceibias.n439 0.189894
R15377 commonsourceibias.n441 commonsourceibias.n440 0.189894
R15378 commonsourceibias.n441 commonsourceibias.n410 0.189894
R15379 commonsourceibias.n447 commonsourceibias.n410 0.189894
R15380 commonsourceibias.n448 commonsourceibias.n447 0.189894
R15381 commonsourceibias.n449 commonsourceibias.n448 0.189894
R15382 commonsourceibias.n449 commonsourceibias.n408 0.189894
R15383 commonsourceibias.n454 commonsourceibias.n408 0.189894
R15384 commonsourceibias.n455 commonsourceibias.n454 0.189894
R15385 commonsourceibias.n456 commonsourceibias.n455 0.189894
R15386 commonsourceibias.n456 commonsourceibias.n406 0.189894
R15387 commonsourceibias.n461 commonsourceibias.n406 0.189894
R15388 commonsourceibias.n462 commonsourceibias.n461 0.189894
R15389 commonsourceibias.n462 commonsourceibias.n404 0.189894
R15390 commonsourceibias.n112 commonsourceibias.n111 0.170955
R15391 commonsourceibias.n113 commonsourceibias.n112 0.170955
R15392 commonsourceibias.n377 commonsourceibias.n301 0.170955
R15393 commonsourceibias.n378 commonsourceibias.n377 0.170955
R15394 CSoutput.n19 CSoutput.t192 184.661
R15395 CSoutput.n78 CSoutput.n77 165.8
R15396 CSoutput.n76 CSoutput.n0 165.8
R15397 CSoutput.n75 CSoutput.n74 165.8
R15398 CSoutput.n73 CSoutput.n72 165.8
R15399 CSoutput.n71 CSoutput.n2 165.8
R15400 CSoutput.n69 CSoutput.n68 165.8
R15401 CSoutput.n67 CSoutput.n3 165.8
R15402 CSoutput.n66 CSoutput.n65 165.8
R15403 CSoutput.n63 CSoutput.n4 165.8
R15404 CSoutput.n61 CSoutput.n60 165.8
R15405 CSoutput.n59 CSoutput.n5 165.8
R15406 CSoutput.n58 CSoutput.n57 165.8
R15407 CSoutput.n55 CSoutput.n6 165.8
R15408 CSoutput.n54 CSoutput.n53 165.8
R15409 CSoutput.n52 CSoutput.n51 165.8
R15410 CSoutput.n50 CSoutput.n8 165.8
R15411 CSoutput.n48 CSoutput.n47 165.8
R15412 CSoutput.n46 CSoutput.n9 165.8
R15413 CSoutput.n45 CSoutput.n44 165.8
R15414 CSoutput.n42 CSoutput.n10 165.8
R15415 CSoutput.n41 CSoutput.n40 165.8
R15416 CSoutput.n39 CSoutput.n38 165.8
R15417 CSoutput.n37 CSoutput.n12 165.8
R15418 CSoutput.n35 CSoutput.n34 165.8
R15419 CSoutput.n33 CSoutput.n13 165.8
R15420 CSoutput.n32 CSoutput.n31 165.8
R15421 CSoutput.n29 CSoutput.n14 165.8
R15422 CSoutput.n28 CSoutput.n27 165.8
R15423 CSoutput.n26 CSoutput.n25 165.8
R15424 CSoutput.n24 CSoutput.n16 165.8
R15425 CSoutput.n22 CSoutput.n21 165.8
R15426 CSoutput.n20 CSoutput.n17 165.8
R15427 CSoutput.n77 CSoutput.t194 162.194
R15428 CSoutput.n18 CSoutput.t201 120.501
R15429 CSoutput.n23 CSoutput.t203 120.501
R15430 CSoutput.n15 CSoutput.t196 120.501
R15431 CSoutput.n30 CSoutput.t213 120.501
R15432 CSoutput.n36 CSoutput.t204 120.501
R15433 CSoutput.n11 CSoutput.t199 120.501
R15434 CSoutput.n43 CSoutput.t193 120.501
R15435 CSoutput.n49 CSoutput.t210 120.501
R15436 CSoutput.n7 CSoutput.t207 120.501
R15437 CSoutput.n56 CSoutput.t197 120.501
R15438 CSoutput.n62 CSoutput.t212 120.501
R15439 CSoutput.n64 CSoutput.t208 120.501
R15440 CSoutput.n70 CSoutput.t200 120.501
R15441 CSoutput.n1 CSoutput.t202 120.501
R15442 CSoutput.n330 CSoutput.n328 103.469
R15443 CSoutput.n310 CSoutput.n308 103.469
R15444 CSoutput.n291 CSoutput.n289 103.469
R15445 CSoutput.n120 CSoutput.n118 103.469
R15446 CSoutput.n100 CSoutput.n98 103.469
R15447 CSoutput.n81 CSoutput.n79 103.469
R15448 CSoutput.n344 CSoutput.n343 103.111
R15449 CSoutput.n342 CSoutput.n341 103.111
R15450 CSoutput.n340 CSoutput.n339 103.111
R15451 CSoutput.n338 CSoutput.n337 103.111
R15452 CSoutput.n336 CSoutput.n335 103.111
R15453 CSoutput.n334 CSoutput.n333 103.111
R15454 CSoutput.n332 CSoutput.n331 103.111
R15455 CSoutput.n330 CSoutput.n329 103.111
R15456 CSoutput.n326 CSoutput.n325 103.111
R15457 CSoutput.n324 CSoutput.n323 103.111
R15458 CSoutput.n322 CSoutput.n321 103.111
R15459 CSoutput.n320 CSoutput.n319 103.111
R15460 CSoutput.n318 CSoutput.n317 103.111
R15461 CSoutput.n316 CSoutput.n315 103.111
R15462 CSoutput.n314 CSoutput.n313 103.111
R15463 CSoutput.n312 CSoutput.n311 103.111
R15464 CSoutput.n310 CSoutput.n309 103.111
R15465 CSoutput.n307 CSoutput.n306 103.111
R15466 CSoutput.n305 CSoutput.n304 103.111
R15467 CSoutput.n303 CSoutput.n302 103.111
R15468 CSoutput.n301 CSoutput.n300 103.111
R15469 CSoutput.n299 CSoutput.n298 103.111
R15470 CSoutput.n297 CSoutput.n296 103.111
R15471 CSoutput.n295 CSoutput.n294 103.111
R15472 CSoutput.n293 CSoutput.n292 103.111
R15473 CSoutput.n291 CSoutput.n290 103.111
R15474 CSoutput.n120 CSoutput.n119 103.111
R15475 CSoutput.n122 CSoutput.n121 103.111
R15476 CSoutput.n124 CSoutput.n123 103.111
R15477 CSoutput.n126 CSoutput.n125 103.111
R15478 CSoutput.n128 CSoutput.n127 103.111
R15479 CSoutput.n130 CSoutput.n129 103.111
R15480 CSoutput.n132 CSoutput.n131 103.111
R15481 CSoutput.n134 CSoutput.n133 103.111
R15482 CSoutput.n136 CSoutput.n135 103.111
R15483 CSoutput.n100 CSoutput.n99 103.111
R15484 CSoutput.n102 CSoutput.n101 103.111
R15485 CSoutput.n104 CSoutput.n103 103.111
R15486 CSoutput.n106 CSoutput.n105 103.111
R15487 CSoutput.n108 CSoutput.n107 103.111
R15488 CSoutput.n110 CSoutput.n109 103.111
R15489 CSoutput.n112 CSoutput.n111 103.111
R15490 CSoutput.n114 CSoutput.n113 103.111
R15491 CSoutput.n116 CSoutput.n115 103.111
R15492 CSoutput.n81 CSoutput.n80 103.111
R15493 CSoutput.n83 CSoutput.n82 103.111
R15494 CSoutput.n85 CSoutput.n84 103.111
R15495 CSoutput.n87 CSoutput.n86 103.111
R15496 CSoutput.n89 CSoutput.n88 103.111
R15497 CSoutput.n91 CSoutput.n90 103.111
R15498 CSoutput.n93 CSoutput.n92 103.111
R15499 CSoutput.n95 CSoutput.n94 103.111
R15500 CSoutput.n97 CSoutput.n96 103.111
R15501 CSoutput.n346 CSoutput.n345 103.111
R15502 CSoutput.n374 CSoutput.n372 81.5057
R15503 CSoutput.n362 CSoutput.n360 81.5057
R15504 CSoutput.n351 CSoutput.n349 81.5057
R15505 CSoutput.n410 CSoutput.n408 81.5057
R15506 CSoutput.n398 CSoutput.n396 81.5057
R15507 CSoutput.n387 CSoutput.n385 81.5057
R15508 CSoutput.n382 CSoutput.n381 80.9324
R15509 CSoutput.n380 CSoutput.n379 80.9324
R15510 CSoutput.n378 CSoutput.n377 80.9324
R15511 CSoutput.n376 CSoutput.n375 80.9324
R15512 CSoutput.n374 CSoutput.n373 80.9324
R15513 CSoutput.n370 CSoutput.n369 80.9324
R15514 CSoutput.n368 CSoutput.n367 80.9324
R15515 CSoutput.n366 CSoutput.n365 80.9324
R15516 CSoutput.n364 CSoutput.n363 80.9324
R15517 CSoutput.n362 CSoutput.n361 80.9324
R15518 CSoutput.n359 CSoutput.n358 80.9324
R15519 CSoutput.n357 CSoutput.n356 80.9324
R15520 CSoutput.n355 CSoutput.n354 80.9324
R15521 CSoutput.n353 CSoutput.n352 80.9324
R15522 CSoutput.n351 CSoutput.n350 80.9324
R15523 CSoutput.n410 CSoutput.n409 80.9324
R15524 CSoutput.n412 CSoutput.n411 80.9324
R15525 CSoutput.n414 CSoutput.n413 80.9324
R15526 CSoutput.n416 CSoutput.n415 80.9324
R15527 CSoutput.n418 CSoutput.n417 80.9324
R15528 CSoutput.n398 CSoutput.n397 80.9324
R15529 CSoutput.n400 CSoutput.n399 80.9324
R15530 CSoutput.n402 CSoutput.n401 80.9324
R15531 CSoutput.n404 CSoutput.n403 80.9324
R15532 CSoutput.n406 CSoutput.n405 80.9324
R15533 CSoutput.n387 CSoutput.n386 80.9324
R15534 CSoutput.n389 CSoutput.n388 80.9324
R15535 CSoutput.n391 CSoutput.n390 80.9324
R15536 CSoutput.n393 CSoutput.n392 80.9324
R15537 CSoutput.n395 CSoutput.n394 80.9324
R15538 CSoutput.n25 CSoutput.n24 48.1486
R15539 CSoutput.n69 CSoutput.n3 48.1486
R15540 CSoutput.n38 CSoutput.n37 48.1486
R15541 CSoutput.n42 CSoutput.n41 48.1486
R15542 CSoutput.n51 CSoutput.n50 48.1486
R15543 CSoutput.n55 CSoutput.n54 48.1486
R15544 CSoutput.n22 CSoutput.n17 46.462
R15545 CSoutput.n72 CSoutput.n71 46.462
R15546 CSoutput.n20 CSoutput.n19 44.9055
R15547 CSoutput.n29 CSoutput.n28 43.7635
R15548 CSoutput.n65 CSoutput.n63 43.7635
R15549 CSoutput.n35 CSoutput.n13 41.7396
R15550 CSoutput.n57 CSoutput.n5 41.7396
R15551 CSoutput.n44 CSoutput.n9 37.0171
R15552 CSoutput.n48 CSoutput.n9 37.0171
R15553 CSoutput.n76 CSoutput.n75 34.9932
R15554 CSoutput.n31 CSoutput.n13 32.2947
R15555 CSoutput.n61 CSoutput.n5 32.2947
R15556 CSoutput.n30 CSoutput.n29 29.6014
R15557 CSoutput.n63 CSoutput.n62 29.6014
R15558 CSoutput.n19 CSoutput.n18 28.4085
R15559 CSoutput.n18 CSoutput.n17 25.1176
R15560 CSoutput.n72 CSoutput.n1 25.1176
R15561 CSoutput.n43 CSoutput.n42 22.0922
R15562 CSoutput.n50 CSoutput.n49 22.0922
R15563 CSoutput.n77 CSoutput.n76 21.8586
R15564 CSoutput.n37 CSoutput.n36 18.9681
R15565 CSoutput.n56 CSoutput.n55 18.9681
R15566 CSoutput.n25 CSoutput.n15 17.6292
R15567 CSoutput.n64 CSoutput.n3 17.6292
R15568 CSoutput.n24 CSoutput.n23 15.844
R15569 CSoutput.n70 CSoutput.n69 15.844
R15570 CSoutput.n38 CSoutput.n11 14.5051
R15571 CSoutput.n54 CSoutput.n7 14.5051
R15572 CSoutput.n421 CSoutput.n78 11.4967
R15573 CSoutput.n41 CSoutput.n11 11.3811
R15574 CSoutput.n51 CSoutput.n7 11.3811
R15575 CSoutput.n23 CSoutput.n22 10.0422
R15576 CSoutput.n71 CSoutput.n70 10.0422
R15577 CSoutput.n327 CSoutput.n307 9.25285
R15578 CSoutput.n117 CSoutput.n97 9.25285
R15579 CSoutput.n371 CSoutput.n359 8.98182
R15580 CSoutput.n407 CSoutput.n395 8.98182
R15581 CSoutput.n384 CSoutput.n348 8.71742
R15582 CSoutput.n28 CSoutput.n15 8.25698
R15583 CSoutput.n65 CSoutput.n64 8.25698
R15584 CSoutput.n348 CSoutput.n347 7.12641
R15585 CSoutput.n138 CSoutput.n137 7.12641
R15586 CSoutput.n36 CSoutput.n35 6.91809
R15587 CSoutput.n57 CSoutput.n56 6.91809
R15588 CSoutput.n384 CSoutput.n383 6.02792
R15589 CSoutput.n420 CSoutput.n419 6.02792
R15590 CSoutput.n383 CSoutput.n382 5.25266
R15591 CSoutput.n371 CSoutput.n370 5.25266
R15592 CSoutput.n419 CSoutput.n418 5.25266
R15593 CSoutput.n407 CSoutput.n406 5.25266
R15594 CSoutput.n347 CSoutput.n346 5.1449
R15595 CSoutput.n327 CSoutput.n326 5.1449
R15596 CSoutput.n137 CSoutput.n136 5.1449
R15597 CSoutput.n117 CSoutput.n116 5.1449
R15598 CSoutput.n421 CSoutput.n138 4.91834
R15599 CSoutput.n229 CSoutput.n182 4.5005
R15600 CSoutput.n198 CSoutput.n182 4.5005
R15601 CSoutput.n193 CSoutput.n177 4.5005
R15602 CSoutput.n193 CSoutput.n179 4.5005
R15603 CSoutput.n193 CSoutput.n176 4.5005
R15604 CSoutput.n193 CSoutput.n180 4.5005
R15605 CSoutput.n193 CSoutput.n175 4.5005
R15606 CSoutput.n193 CSoutput.t198 4.5005
R15607 CSoutput.n193 CSoutput.n174 4.5005
R15608 CSoutput.n193 CSoutput.n181 4.5005
R15609 CSoutput.n193 CSoutput.n182 4.5005
R15610 CSoutput.n191 CSoutput.n177 4.5005
R15611 CSoutput.n191 CSoutput.n179 4.5005
R15612 CSoutput.n191 CSoutput.n176 4.5005
R15613 CSoutput.n191 CSoutput.n180 4.5005
R15614 CSoutput.n191 CSoutput.n175 4.5005
R15615 CSoutput.n191 CSoutput.t198 4.5005
R15616 CSoutput.n191 CSoutput.n174 4.5005
R15617 CSoutput.n191 CSoutput.n181 4.5005
R15618 CSoutput.n191 CSoutput.n182 4.5005
R15619 CSoutput.n190 CSoutput.n177 4.5005
R15620 CSoutput.n190 CSoutput.n179 4.5005
R15621 CSoutput.n190 CSoutput.n176 4.5005
R15622 CSoutput.n190 CSoutput.n180 4.5005
R15623 CSoutput.n190 CSoutput.n175 4.5005
R15624 CSoutput.n190 CSoutput.t198 4.5005
R15625 CSoutput.n190 CSoutput.n174 4.5005
R15626 CSoutput.n190 CSoutput.n181 4.5005
R15627 CSoutput.n190 CSoutput.n182 4.5005
R15628 CSoutput.n275 CSoutput.n177 4.5005
R15629 CSoutput.n275 CSoutput.n179 4.5005
R15630 CSoutput.n275 CSoutput.n176 4.5005
R15631 CSoutput.n275 CSoutput.n180 4.5005
R15632 CSoutput.n275 CSoutput.n175 4.5005
R15633 CSoutput.n275 CSoutput.t198 4.5005
R15634 CSoutput.n275 CSoutput.n174 4.5005
R15635 CSoutput.n275 CSoutput.n181 4.5005
R15636 CSoutput.n275 CSoutput.n182 4.5005
R15637 CSoutput.n273 CSoutput.n177 4.5005
R15638 CSoutput.n273 CSoutput.n179 4.5005
R15639 CSoutput.n273 CSoutput.n176 4.5005
R15640 CSoutput.n273 CSoutput.n180 4.5005
R15641 CSoutput.n273 CSoutput.n175 4.5005
R15642 CSoutput.n273 CSoutput.t198 4.5005
R15643 CSoutput.n273 CSoutput.n174 4.5005
R15644 CSoutput.n273 CSoutput.n181 4.5005
R15645 CSoutput.n271 CSoutput.n177 4.5005
R15646 CSoutput.n271 CSoutput.n179 4.5005
R15647 CSoutput.n271 CSoutput.n176 4.5005
R15648 CSoutput.n271 CSoutput.n180 4.5005
R15649 CSoutput.n271 CSoutput.n175 4.5005
R15650 CSoutput.n271 CSoutput.t198 4.5005
R15651 CSoutput.n271 CSoutput.n174 4.5005
R15652 CSoutput.n271 CSoutput.n181 4.5005
R15653 CSoutput.n201 CSoutput.n177 4.5005
R15654 CSoutput.n201 CSoutput.n179 4.5005
R15655 CSoutput.n201 CSoutput.n176 4.5005
R15656 CSoutput.n201 CSoutput.n180 4.5005
R15657 CSoutput.n201 CSoutput.n175 4.5005
R15658 CSoutput.n201 CSoutput.t198 4.5005
R15659 CSoutput.n201 CSoutput.n174 4.5005
R15660 CSoutput.n201 CSoutput.n181 4.5005
R15661 CSoutput.n201 CSoutput.n182 4.5005
R15662 CSoutput.n200 CSoutput.n177 4.5005
R15663 CSoutput.n200 CSoutput.n179 4.5005
R15664 CSoutput.n200 CSoutput.n176 4.5005
R15665 CSoutput.n200 CSoutput.n180 4.5005
R15666 CSoutput.n200 CSoutput.n175 4.5005
R15667 CSoutput.n200 CSoutput.t198 4.5005
R15668 CSoutput.n200 CSoutput.n174 4.5005
R15669 CSoutput.n200 CSoutput.n181 4.5005
R15670 CSoutput.n200 CSoutput.n182 4.5005
R15671 CSoutput.n204 CSoutput.n177 4.5005
R15672 CSoutput.n204 CSoutput.n179 4.5005
R15673 CSoutput.n204 CSoutput.n176 4.5005
R15674 CSoutput.n204 CSoutput.n180 4.5005
R15675 CSoutput.n204 CSoutput.n175 4.5005
R15676 CSoutput.n204 CSoutput.t198 4.5005
R15677 CSoutput.n204 CSoutput.n174 4.5005
R15678 CSoutput.n204 CSoutput.n181 4.5005
R15679 CSoutput.n204 CSoutput.n182 4.5005
R15680 CSoutput.n203 CSoutput.n177 4.5005
R15681 CSoutput.n203 CSoutput.n179 4.5005
R15682 CSoutput.n203 CSoutput.n176 4.5005
R15683 CSoutput.n203 CSoutput.n180 4.5005
R15684 CSoutput.n203 CSoutput.n175 4.5005
R15685 CSoutput.n203 CSoutput.t198 4.5005
R15686 CSoutput.n203 CSoutput.n174 4.5005
R15687 CSoutput.n203 CSoutput.n181 4.5005
R15688 CSoutput.n203 CSoutput.n182 4.5005
R15689 CSoutput.n186 CSoutput.n177 4.5005
R15690 CSoutput.n186 CSoutput.n179 4.5005
R15691 CSoutput.n186 CSoutput.n176 4.5005
R15692 CSoutput.n186 CSoutput.n180 4.5005
R15693 CSoutput.n186 CSoutput.n175 4.5005
R15694 CSoutput.n186 CSoutput.t198 4.5005
R15695 CSoutput.n186 CSoutput.n174 4.5005
R15696 CSoutput.n186 CSoutput.n181 4.5005
R15697 CSoutput.n186 CSoutput.n182 4.5005
R15698 CSoutput.n278 CSoutput.n177 4.5005
R15699 CSoutput.n278 CSoutput.n179 4.5005
R15700 CSoutput.n278 CSoutput.n176 4.5005
R15701 CSoutput.n278 CSoutput.n180 4.5005
R15702 CSoutput.n278 CSoutput.n175 4.5005
R15703 CSoutput.n278 CSoutput.t198 4.5005
R15704 CSoutput.n278 CSoutput.n174 4.5005
R15705 CSoutput.n278 CSoutput.n181 4.5005
R15706 CSoutput.n278 CSoutput.n182 4.5005
R15707 CSoutput.n265 CSoutput.n236 4.5005
R15708 CSoutput.n265 CSoutput.n242 4.5005
R15709 CSoutput.n223 CSoutput.n212 4.5005
R15710 CSoutput.n223 CSoutput.n214 4.5005
R15711 CSoutput.n223 CSoutput.n211 4.5005
R15712 CSoutput.n223 CSoutput.n215 4.5005
R15713 CSoutput.n223 CSoutput.n210 4.5005
R15714 CSoutput.n223 CSoutput.t206 4.5005
R15715 CSoutput.n223 CSoutput.n209 4.5005
R15716 CSoutput.n223 CSoutput.n216 4.5005
R15717 CSoutput.n265 CSoutput.n223 4.5005
R15718 CSoutput.n244 CSoutput.n212 4.5005
R15719 CSoutput.n244 CSoutput.n214 4.5005
R15720 CSoutput.n244 CSoutput.n211 4.5005
R15721 CSoutput.n244 CSoutput.n215 4.5005
R15722 CSoutput.n244 CSoutput.n210 4.5005
R15723 CSoutput.n244 CSoutput.t206 4.5005
R15724 CSoutput.n244 CSoutput.n209 4.5005
R15725 CSoutput.n244 CSoutput.n216 4.5005
R15726 CSoutput.n265 CSoutput.n244 4.5005
R15727 CSoutput.n222 CSoutput.n212 4.5005
R15728 CSoutput.n222 CSoutput.n214 4.5005
R15729 CSoutput.n222 CSoutput.n211 4.5005
R15730 CSoutput.n222 CSoutput.n215 4.5005
R15731 CSoutput.n222 CSoutput.n210 4.5005
R15732 CSoutput.n222 CSoutput.t206 4.5005
R15733 CSoutput.n222 CSoutput.n209 4.5005
R15734 CSoutput.n222 CSoutput.n216 4.5005
R15735 CSoutput.n265 CSoutput.n222 4.5005
R15736 CSoutput.n246 CSoutput.n212 4.5005
R15737 CSoutput.n246 CSoutput.n214 4.5005
R15738 CSoutput.n246 CSoutput.n211 4.5005
R15739 CSoutput.n246 CSoutput.n215 4.5005
R15740 CSoutput.n246 CSoutput.n210 4.5005
R15741 CSoutput.n246 CSoutput.t206 4.5005
R15742 CSoutput.n246 CSoutput.n209 4.5005
R15743 CSoutput.n246 CSoutput.n216 4.5005
R15744 CSoutput.n265 CSoutput.n246 4.5005
R15745 CSoutput.n212 CSoutput.n207 4.5005
R15746 CSoutput.n214 CSoutput.n207 4.5005
R15747 CSoutput.n211 CSoutput.n207 4.5005
R15748 CSoutput.n215 CSoutput.n207 4.5005
R15749 CSoutput.n210 CSoutput.n207 4.5005
R15750 CSoutput.t206 CSoutput.n207 4.5005
R15751 CSoutput.n209 CSoutput.n207 4.5005
R15752 CSoutput.n216 CSoutput.n207 4.5005
R15753 CSoutput.n268 CSoutput.n212 4.5005
R15754 CSoutput.n268 CSoutput.n214 4.5005
R15755 CSoutput.n268 CSoutput.n211 4.5005
R15756 CSoutput.n268 CSoutput.n215 4.5005
R15757 CSoutput.n268 CSoutput.n210 4.5005
R15758 CSoutput.n268 CSoutput.t206 4.5005
R15759 CSoutput.n268 CSoutput.n209 4.5005
R15760 CSoutput.n268 CSoutput.n216 4.5005
R15761 CSoutput.n266 CSoutput.n212 4.5005
R15762 CSoutput.n266 CSoutput.n214 4.5005
R15763 CSoutput.n266 CSoutput.n211 4.5005
R15764 CSoutput.n266 CSoutput.n215 4.5005
R15765 CSoutput.n266 CSoutput.n210 4.5005
R15766 CSoutput.n266 CSoutput.t206 4.5005
R15767 CSoutput.n266 CSoutput.n209 4.5005
R15768 CSoutput.n266 CSoutput.n216 4.5005
R15769 CSoutput.n266 CSoutput.n265 4.5005
R15770 CSoutput.n248 CSoutput.n212 4.5005
R15771 CSoutput.n248 CSoutput.n214 4.5005
R15772 CSoutput.n248 CSoutput.n211 4.5005
R15773 CSoutput.n248 CSoutput.n215 4.5005
R15774 CSoutput.n248 CSoutput.n210 4.5005
R15775 CSoutput.n248 CSoutput.t206 4.5005
R15776 CSoutput.n248 CSoutput.n209 4.5005
R15777 CSoutput.n248 CSoutput.n216 4.5005
R15778 CSoutput.n265 CSoutput.n248 4.5005
R15779 CSoutput.n220 CSoutput.n212 4.5005
R15780 CSoutput.n220 CSoutput.n214 4.5005
R15781 CSoutput.n220 CSoutput.n211 4.5005
R15782 CSoutput.n220 CSoutput.n215 4.5005
R15783 CSoutput.n220 CSoutput.n210 4.5005
R15784 CSoutput.n220 CSoutput.t206 4.5005
R15785 CSoutput.n220 CSoutput.n209 4.5005
R15786 CSoutput.n220 CSoutput.n216 4.5005
R15787 CSoutput.n265 CSoutput.n220 4.5005
R15788 CSoutput.n250 CSoutput.n212 4.5005
R15789 CSoutput.n250 CSoutput.n214 4.5005
R15790 CSoutput.n250 CSoutput.n211 4.5005
R15791 CSoutput.n250 CSoutput.n215 4.5005
R15792 CSoutput.n250 CSoutput.n210 4.5005
R15793 CSoutput.n250 CSoutput.t206 4.5005
R15794 CSoutput.n250 CSoutput.n209 4.5005
R15795 CSoutput.n250 CSoutput.n216 4.5005
R15796 CSoutput.n265 CSoutput.n250 4.5005
R15797 CSoutput.n219 CSoutput.n212 4.5005
R15798 CSoutput.n219 CSoutput.n214 4.5005
R15799 CSoutput.n219 CSoutput.n211 4.5005
R15800 CSoutput.n219 CSoutput.n215 4.5005
R15801 CSoutput.n219 CSoutput.n210 4.5005
R15802 CSoutput.n219 CSoutput.t206 4.5005
R15803 CSoutput.n219 CSoutput.n209 4.5005
R15804 CSoutput.n219 CSoutput.n216 4.5005
R15805 CSoutput.n265 CSoutput.n219 4.5005
R15806 CSoutput.n264 CSoutput.n212 4.5005
R15807 CSoutput.n264 CSoutput.n214 4.5005
R15808 CSoutput.n264 CSoutput.n211 4.5005
R15809 CSoutput.n264 CSoutput.n215 4.5005
R15810 CSoutput.n264 CSoutput.n210 4.5005
R15811 CSoutput.n264 CSoutput.t206 4.5005
R15812 CSoutput.n264 CSoutput.n209 4.5005
R15813 CSoutput.n264 CSoutput.n216 4.5005
R15814 CSoutput.n265 CSoutput.n264 4.5005
R15815 CSoutput.n263 CSoutput.n148 4.5005
R15816 CSoutput.n164 CSoutput.n148 4.5005
R15817 CSoutput.n159 CSoutput.n143 4.5005
R15818 CSoutput.n159 CSoutput.n145 4.5005
R15819 CSoutput.n159 CSoutput.n142 4.5005
R15820 CSoutput.n159 CSoutput.n146 4.5005
R15821 CSoutput.n159 CSoutput.n141 4.5005
R15822 CSoutput.n159 CSoutput.t209 4.5005
R15823 CSoutput.n159 CSoutput.n140 4.5005
R15824 CSoutput.n159 CSoutput.n147 4.5005
R15825 CSoutput.n159 CSoutput.n148 4.5005
R15826 CSoutput.n157 CSoutput.n143 4.5005
R15827 CSoutput.n157 CSoutput.n145 4.5005
R15828 CSoutput.n157 CSoutput.n142 4.5005
R15829 CSoutput.n157 CSoutput.n146 4.5005
R15830 CSoutput.n157 CSoutput.n141 4.5005
R15831 CSoutput.n157 CSoutput.t209 4.5005
R15832 CSoutput.n157 CSoutput.n140 4.5005
R15833 CSoutput.n157 CSoutput.n147 4.5005
R15834 CSoutput.n157 CSoutput.n148 4.5005
R15835 CSoutput.n156 CSoutput.n143 4.5005
R15836 CSoutput.n156 CSoutput.n145 4.5005
R15837 CSoutput.n156 CSoutput.n142 4.5005
R15838 CSoutput.n156 CSoutput.n146 4.5005
R15839 CSoutput.n156 CSoutput.n141 4.5005
R15840 CSoutput.n156 CSoutput.t209 4.5005
R15841 CSoutput.n156 CSoutput.n140 4.5005
R15842 CSoutput.n156 CSoutput.n147 4.5005
R15843 CSoutput.n156 CSoutput.n148 4.5005
R15844 CSoutput.n285 CSoutput.n143 4.5005
R15845 CSoutput.n285 CSoutput.n145 4.5005
R15846 CSoutput.n285 CSoutput.n142 4.5005
R15847 CSoutput.n285 CSoutput.n146 4.5005
R15848 CSoutput.n285 CSoutput.n141 4.5005
R15849 CSoutput.n285 CSoutput.t209 4.5005
R15850 CSoutput.n285 CSoutput.n140 4.5005
R15851 CSoutput.n285 CSoutput.n147 4.5005
R15852 CSoutput.n285 CSoutput.n148 4.5005
R15853 CSoutput.n283 CSoutput.n143 4.5005
R15854 CSoutput.n283 CSoutput.n145 4.5005
R15855 CSoutput.n283 CSoutput.n142 4.5005
R15856 CSoutput.n283 CSoutput.n146 4.5005
R15857 CSoutput.n283 CSoutput.n141 4.5005
R15858 CSoutput.n283 CSoutput.t209 4.5005
R15859 CSoutput.n283 CSoutput.n140 4.5005
R15860 CSoutput.n283 CSoutput.n147 4.5005
R15861 CSoutput.n281 CSoutput.n143 4.5005
R15862 CSoutput.n281 CSoutput.n145 4.5005
R15863 CSoutput.n281 CSoutput.n142 4.5005
R15864 CSoutput.n281 CSoutput.n146 4.5005
R15865 CSoutput.n281 CSoutput.n141 4.5005
R15866 CSoutput.n281 CSoutput.t209 4.5005
R15867 CSoutput.n281 CSoutput.n140 4.5005
R15868 CSoutput.n281 CSoutput.n147 4.5005
R15869 CSoutput.n167 CSoutput.n143 4.5005
R15870 CSoutput.n167 CSoutput.n145 4.5005
R15871 CSoutput.n167 CSoutput.n142 4.5005
R15872 CSoutput.n167 CSoutput.n146 4.5005
R15873 CSoutput.n167 CSoutput.n141 4.5005
R15874 CSoutput.n167 CSoutput.t209 4.5005
R15875 CSoutput.n167 CSoutput.n140 4.5005
R15876 CSoutput.n167 CSoutput.n147 4.5005
R15877 CSoutput.n167 CSoutput.n148 4.5005
R15878 CSoutput.n166 CSoutput.n143 4.5005
R15879 CSoutput.n166 CSoutput.n145 4.5005
R15880 CSoutput.n166 CSoutput.n142 4.5005
R15881 CSoutput.n166 CSoutput.n146 4.5005
R15882 CSoutput.n166 CSoutput.n141 4.5005
R15883 CSoutput.n166 CSoutput.t209 4.5005
R15884 CSoutput.n166 CSoutput.n140 4.5005
R15885 CSoutput.n166 CSoutput.n147 4.5005
R15886 CSoutput.n166 CSoutput.n148 4.5005
R15887 CSoutput.n170 CSoutput.n143 4.5005
R15888 CSoutput.n170 CSoutput.n145 4.5005
R15889 CSoutput.n170 CSoutput.n142 4.5005
R15890 CSoutput.n170 CSoutput.n146 4.5005
R15891 CSoutput.n170 CSoutput.n141 4.5005
R15892 CSoutput.n170 CSoutput.t209 4.5005
R15893 CSoutput.n170 CSoutput.n140 4.5005
R15894 CSoutput.n170 CSoutput.n147 4.5005
R15895 CSoutput.n170 CSoutput.n148 4.5005
R15896 CSoutput.n169 CSoutput.n143 4.5005
R15897 CSoutput.n169 CSoutput.n145 4.5005
R15898 CSoutput.n169 CSoutput.n142 4.5005
R15899 CSoutput.n169 CSoutput.n146 4.5005
R15900 CSoutput.n169 CSoutput.n141 4.5005
R15901 CSoutput.n169 CSoutput.t209 4.5005
R15902 CSoutput.n169 CSoutput.n140 4.5005
R15903 CSoutput.n169 CSoutput.n147 4.5005
R15904 CSoutput.n169 CSoutput.n148 4.5005
R15905 CSoutput.n152 CSoutput.n143 4.5005
R15906 CSoutput.n152 CSoutput.n145 4.5005
R15907 CSoutput.n152 CSoutput.n142 4.5005
R15908 CSoutput.n152 CSoutput.n146 4.5005
R15909 CSoutput.n152 CSoutput.n141 4.5005
R15910 CSoutput.n152 CSoutput.t209 4.5005
R15911 CSoutput.n152 CSoutput.n140 4.5005
R15912 CSoutput.n152 CSoutput.n147 4.5005
R15913 CSoutput.n152 CSoutput.n148 4.5005
R15914 CSoutput.n288 CSoutput.n143 4.5005
R15915 CSoutput.n288 CSoutput.n145 4.5005
R15916 CSoutput.n288 CSoutput.n142 4.5005
R15917 CSoutput.n288 CSoutput.n146 4.5005
R15918 CSoutput.n288 CSoutput.n141 4.5005
R15919 CSoutput.n288 CSoutput.t209 4.5005
R15920 CSoutput.n288 CSoutput.n140 4.5005
R15921 CSoutput.n288 CSoutput.n147 4.5005
R15922 CSoutput.n288 CSoutput.n148 4.5005
R15923 CSoutput.n347 CSoutput.n327 4.10845
R15924 CSoutput.n137 CSoutput.n117 4.10845
R15925 CSoutput.n345 CSoutput.t121 4.06363
R15926 CSoutput.n345 CSoutput.t177 4.06363
R15927 CSoutput.n343 CSoutput.t111 4.06363
R15928 CSoutput.n343 CSoutput.t74 4.06363
R15929 CSoutput.n341 CSoutput.t150 4.06363
R15930 CSoutput.n341 CSoutput.t187 4.06363
R15931 CSoutput.n339 CSoutput.t155 4.06363
R15932 CSoutput.n339 CSoutput.t144 4.06363
R15933 CSoutput.n337 CSoutput.t91 4.06363
R15934 CSoutput.n337 CSoutput.t188 4.06363
R15935 CSoutput.n335 CSoutput.t146 4.06363
R15936 CSoutput.n335 CSoutput.t157 4.06363
R15937 CSoutput.n333 CSoutput.t115 4.06363
R15938 CSoutput.n333 CSoutput.t105 4.06363
R15939 CSoutput.n331 CSoutput.t75 4.06363
R15940 CSoutput.n331 CSoutput.t164 4.06363
R15941 CSoutput.n329 CSoutput.t126 4.06363
R15942 CSoutput.n329 CSoutput.t106 4.06363
R15943 CSoutput.n328 CSoutput.t149 4.06363
R15944 CSoutput.n328 CSoutput.t137 4.06363
R15945 CSoutput.n325 CSoutput.t158 4.06363
R15946 CSoutput.n325 CSoutput.t122 4.06363
R15947 CSoutput.n323 CSoutput.t127 4.06363
R15948 CSoutput.n323 CSoutput.t107 4.06363
R15949 CSoutput.n321 CSoutput.t152 4.06363
R15950 CSoutput.n321 CSoutput.t190 4.06363
R15951 CSoutput.n319 CSoutput.t128 4.06363
R15952 CSoutput.n319 CSoutput.t113 4.06363
R15953 CSoutput.n317 CSoutput.t131 4.06363
R15954 CSoutput.n317 CSoutput.t180 4.06363
R15955 CSoutput.n315 CSoutput.t147 4.06363
R15956 CSoutput.n315 CSoutput.t176 4.06363
R15957 CSoutput.n313 CSoutput.t119 4.06363
R15958 CSoutput.n313 CSoutput.t168 4.06363
R15959 CSoutput.n311 CSoutput.t108 4.06363
R15960 CSoutput.n311 CSoutput.t166 4.06363
R15961 CSoutput.n309 CSoutput.t179 4.06363
R15962 CSoutput.n309 CSoutput.t171 4.06363
R15963 CSoutput.n308 CSoutput.t153 4.06363
R15964 CSoutput.n308 CSoutput.t80 4.06363
R15965 CSoutput.n306 CSoutput.t83 4.06363
R15966 CSoutput.n306 CSoutput.t84 4.06363
R15967 CSoutput.n304 CSoutput.t99 4.06363
R15968 CSoutput.n304 CSoutput.t109 4.06363
R15969 CSoutput.n302 CSoutput.t138 4.06363
R15970 CSoutput.n302 CSoutput.t114 4.06363
R15971 CSoutput.n300 CSoutput.t78 4.06363
R15972 CSoutput.n300 CSoutput.t184 4.06363
R15973 CSoutput.n298 CSoutput.t169 4.06363
R15974 CSoutput.n298 CSoutput.t174 4.06363
R15975 CSoutput.n296 CSoutput.t82 4.06363
R15976 CSoutput.n296 CSoutput.t134 4.06363
R15977 CSoutput.n294 CSoutput.t92 4.06363
R15978 CSoutput.n294 CSoutput.t96 4.06363
R15979 CSoutput.n292 CSoutput.t183 4.06363
R15980 CSoutput.n292 CSoutput.t163 4.06363
R15981 CSoutput.n290 CSoutput.t76 4.06363
R15982 CSoutput.n290 CSoutput.t189 4.06363
R15983 CSoutput.n289 CSoutput.t123 4.06363
R15984 CSoutput.n289 CSoutput.t135 4.06363
R15985 CSoutput.n118 CSoutput.t141 4.06363
R15986 CSoutput.n118 CSoutput.t94 4.06363
R15987 CSoutput.n119 CSoutput.t97 4.06363
R15988 CSoutput.n119 CSoutput.t143 4.06363
R15989 CSoutput.n121 CSoutput.t161 4.06363
R15990 CSoutput.n121 CSoutput.t89 4.06363
R15991 CSoutput.n123 CSoutput.t120 4.06363
R15992 CSoutput.n123 CSoutput.t165 4.06363
R15993 CSoutput.n125 CSoutput.t87 4.06363
R15994 CSoutput.n125 CSoutput.t118 4.06363
R15995 CSoutput.n127 CSoutput.t156 4.06363
R15996 CSoutput.n127 CSoutput.t101 4.06363
R15997 CSoutput.n129 CSoutput.t140 4.06363
R15998 CSoutput.n129 CSoutput.t85 4.06363
R15999 CSoutput.n131 CSoutput.t142 4.06363
R16000 CSoutput.n131 CSoutput.t95 4.06363
R16001 CSoutput.n133 CSoutput.t88 4.06363
R16002 CSoutput.n133 CSoutput.t148 4.06363
R16003 CSoutput.n135 CSoutput.t162 4.06363
R16004 CSoutput.n135 CSoutput.t160 4.06363
R16005 CSoutput.n98 CSoutput.t173 4.06363
R16006 CSoutput.n98 CSoutput.t103 4.06363
R16007 CSoutput.n99 CSoutput.t145 4.06363
R16008 CSoutput.n99 CSoutput.t117 4.06363
R16009 CSoutput.n101 CSoutput.t132 4.06363
R16010 CSoutput.n101 CSoutput.t178 4.06363
R16011 CSoutput.n103 CSoutput.t167 4.06363
R16012 CSoutput.n103 CSoutput.t191 4.06363
R16013 CSoutput.n105 CSoutput.t130 4.06363
R16014 CSoutput.n105 CSoutput.t90 4.06363
R16015 CSoutput.n107 CSoutput.t175 4.06363
R16016 CSoutput.n107 CSoutput.t98 4.06363
R16017 CSoutput.n109 CSoutput.t81 4.06363
R16018 CSoutput.n109 CSoutput.t182 4.06363
R16019 CSoutput.n111 CSoutput.t116 4.06363
R16020 CSoutput.n111 CSoutput.t104 4.06363
R16021 CSoutput.n113 CSoutput.t100 4.06363
R16022 CSoutput.n113 CSoutput.t151 4.06363
R16023 CSoutput.n115 CSoutput.t133 4.06363
R16024 CSoutput.n115 CSoutput.t125 4.06363
R16025 CSoutput.n79 CSoutput.t181 4.06363
R16026 CSoutput.n79 CSoutput.t124 4.06363
R16027 CSoutput.n80 CSoutput.t102 4.06363
R16028 CSoutput.n80 CSoutput.t77 4.06363
R16029 CSoutput.n82 CSoutput.t186 4.06363
R16030 CSoutput.n82 CSoutput.t129 4.06363
R16031 CSoutput.n84 CSoutput.t110 4.06363
R16032 CSoutput.n84 CSoutput.t112 4.06363
R16033 CSoutput.n86 CSoutput.t172 4.06363
R16034 CSoutput.n86 CSoutput.t72 4.06363
R16035 CSoutput.n88 CSoutput.t136 4.06363
R16036 CSoutput.n88 CSoutput.t170 4.06363
R16037 CSoutput.n90 CSoutput.t185 4.06363
R16038 CSoutput.n90 CSoutput.t79 4.06363
R16039 CSoutput.n92 CSoutput.t159 4.06363
R16040 CSoutput.n92 CSoutput.t139 4.06363
R16041 CSoutput.n94 CSoutput.t154 4.06363
R16042 CSoutput.n94 CSoutput.t93 4.06363
R16043 CSoutput.n96 CSoutput.t86 4.06363
R16044 CSoutput.n96 CSoutput.t73 4.06363
R16045 CSoutput.n44 CSoutput.n43 3.79402
R16046 CSoutput.n49 CSoutput.n48 3.79402
R16047 CSoutput.n421 CSoutput.n420 3.78008
R16048 CSoutput.n383 CSoutput.n371 3.72967
R16049 CSoutput.n419 CSoutput.n407 3.72967
R16050 CSoutput.n348 CSoutput.n138 3.19963
R16051 CSoutput.n381 CSoutput.t17 2.82907
R16052 CSoutput.n381 CSoutput.t21 2.82907
R16053 CSoutput.n379 CSoutput.t16 2.82907
R16054 CSoutput.n379 CSoutput.t71 2.82907
R16055 CSoutput.n377 CSoutput.t31 2.82907
R16056 CSoutput.n377 CSoutput.t11 2.82907
R16057 CSoutput.n375 CSoutput.t4 2.82907
R16058 CSoutput.n375 CSoutput.t51 2.82907
R16059 CSoutput.n373 CSoutput.t23 2.82907
R16060 CSoutput.n373 CSoutput.t26 2.82907
R16061 CSoutput.n372 CSoutput.t10 2.82907
R16062 CSoutput.n372 CSoutput.t62 2.82907
R16063 CSoutput.n369 CSoutput.t3 2.82907
R16064 CSoutput.n369 CSoutput.t49 2.82907
R16065 CSoutput.n367 CSoutput.t48 2.82907
R16066 CSoutput.n367 CSoutput.t36 2.82907
R16067 CSoutput.n365 CSoutput.t60 2.82907
R16068 CSoutput.n365 CSoutput.t1 2.82907
R16069 CSoutput.n363 CSoutput.t2 2.82907
R16070 CSoutput.n363 CSoutput.t54 2.82907
R16071 CSoutput.n361 CSoutput.t9 2.82907
R16072 CSoutput.n361 CSoutput.t59 2.82907
R16073 CSoutput.n360 CSoutput.t65 2.82907
R16074 CSoutput.n360 CSoutput.t0 2.82907
R16075 CSoutput.n358 CSoutput.t39 2.82907
R16076 CSoutput.n358 CSoutput.t46 2.82907
R16077 CSoutput.n356 CSoutput.t32 2.82907
R16078 CSoutput.n356 CSoutput.t61 2.82907
R16079 CSoutput.n354 CSoutput.t42 2.82907
R16080 CSoutput.n354 CSoutput.t25 2.82907
R16081 CSoutput.n352 CSoutput.t18 2.82907
R16082 CSoutput.n352 CSoutput.t33 2.82907
R16083 CSoutput.n350 CSoutput.t24 2.82907
R16084 CSoutput.n350 CSoutput.t29 2.82907
R16085 CSoutput.n349 CSoutput.t30 2.82907
R16086 CSoutput.n349 CSoutput.t68 2.82907
R16087 CSoutput.n408 CSoutput.t38 2.82907
R16088 CSoutput.n408 CSoutput.t56 2.82907
R16089 CSoutput.n409 CSoutput.t19 2.82907
R16090 CSoutput.n409 CSoutput.t28 2.82907
R16091 CSoutput.n411 CSoutput.t34 2.82907
R16092 CSoutput.n411 CSoutput.t43 2.82907
R16093 CSoutput.n413 CSoutput.t57 2.82907
R16094 CSoutput.n413 CSoutput.t37 2.82907
R16095 CSoutput.n415 CSoutput.t41 2.82907
R16096 CSoutput.n415 CSoutput.t66 2.82907
R16097 CSoutput.n417 CSoutput.t6 2.82907
R16098 CSoutput.n417 CSoutput.t22 2.82907
R16099 CSoutput.n396 CSoutput.t12 2.82907
R16100 CSoutput.n396 CSoutput.t7 2.82907
R16101 CSoutput.n397 CSoutput.t5 2.82907
R16102 CSoutput.n397 CSoutput.t69 2.82907
R16103 CSoutput.n399 CSoutput.t70 2.82907
R16104 CSoutput.n399 CSoutput.t13 2.82907
R16105 CSoutput.n401 CSoutput.t14 2.82907
R16106 CSoutput.n401 CSoutput.t45 2.82907
R16107 CSoutput.n403 CSoutput.t44 2.82907
R16108 CSoutput.n403 CSoutput.t64 2.82907
R16109 CSoutput.n405 CSoutput.t67 2.82907
R16110 CSoutput.n405 CSoutput.t58 2.82907
R16111 CSoutput.n385 CSoutput.t20 2.82907
R16112 CSoutput.n385 CSoutput.t50 2.82907
R16113 CSoutput.n386 CSoutput.t47 2.82907
R16114 CSoutput.n386 CSoutput.t35 2.82907
R16115 CSoutput.n388 CSoutput.t53 2.82907
R16116 CSoutput.n388 CSoutput.t27 2.82907
R16117 CSoutput.n390 CSoutput.t40 2.82907
R16118 CSoutput.n390 CSoutput.t63 2.82907
R16119 CSoutput.n392 CSoutput.t15 2.82907
R16120 CSoutput.n392 CSoutput.t52 2.82907
R16121 CSoutput.n394 CSoutput.t8 2.82907
R16122 CSoutput.n394 CSoutput.t55 2.82907
R16123 CSoutput.n420 CSoutput.n384 2.75627
R16124 CSoutput.n75 CSoutput.n1 2.45513
R16125 CSoutput.n229 CSoutput.n227 2.251
R16126 CSoutput.n229 CSoutput.n226 2.251
R16127 CSoutput.n229 CSoutput.n225 2.251
R16128 CSoutput.n229 CSoutput.n224 2.251
R16129 CSoutput.n198 CSoutput.n197 2.251
R16130 CSoutput.n198 CSoutput.n196 2.251
R16131 CSoutput.n198 CSoutput.n195 2.251
R16132 CSoutput.n198 CSoutput.n194 2.251
R16133 CSoutput.n271 CSoutput.n270 2.251
R16134 CSoutput.n236 CSoutput.n234 2.251
R16135 CSoutput.n236 CSoutput.n233 2.251
R16136 CSoutput.n236 CSoutput.n232 2.251
R16137 CSoutput.n254 CSoutput.n236 2.251
R16138 CSoutput.n242 CSoutput.n241 2.251
R16139 CSoutput.n242 CSoutput.n240 2.251
R16140 CSoutput.n242 CSoutput.n239 2.251
R16141 CSoutput.n242 CSoutput.n238 2.251
R16142 CSoutput.n268 CSoutput.n208 2.251
R16143 CSoutput.n263 CSoutput.n261 2.251
R16144 CSoutput.n263 CSoutput.n260 2.251
R16145 CSoutput.n263 CSoutput.n259 2.251
R16146 CSoutput.n263 CSoutput.n258 2.251
R16147 CSoutput.n164 CSoutput.n163 2.251
R16148 CSoutput.n164 CSoutput.n162 2.251
R16149 CSoutput.n164 CSoutput.n161 2.251
R16150 CSoutput.n164 CSoutput.n160 2.251
R16151 CSoutput.n281 CSoutput.n280 2.251
R16152 CSoutput.n198 CSoutput.n178 2.2505
R16153 CSoutput.n193 CSoutput.n178 2.2505
R16154 CSoutput.n191 CSoutput.n178 2.2505
R16155 CSoutput.n190 CSoutput.n178 2.2505
R16156 CSoutput.n275 CSoutput.n178 2.2505
R16157 CSoutput.n273 CSoutput.n178 2.2505
R16158 CSoutput.n271 CSoutput.n178 2.2505
R16159 CSoutput.n201 CSoutput.n178 2.2505
R16160 CSoutput.n200 CSoutput.n178 2.2505
R16161 CSoutput.n204 CSoutput.n178 2.2505
R16162 CSoutput.n203 CSoutput.n178 2.2505
R16163 CSoutput.n186 CSoutput.n178 2.2505
R16164 CSoutput.n278 CSoutput.n178 2.2505
R16165 CSoutput.n278 CSoutput.n277 2.2505
R16166 CSoutput.n242 CSoutput.n213 2.2505
R16167 CSoutput.n223 CSoutput.n213 2.2505
R16168 CSoutput.n244 CSoutput.n213 2.2505
R16169 CSoutput.n222 CSoutput.n213 2.2505
R16170 CSoutput.n246 CSoutput.n213 2.2505
R16171 CSoutput.n213 CSoutput.n207 2.2505
R16172 CSoutput.n268 CSoutput.n213 2.2505
R16173 CSoutput.n266 CSoutput.n213 2.2505
R16174 CSoutput.n248 CSoutput.n213 2.2505
R16175 CSoutput.n220 CSoutput.n213 2.2505
R16176 CSoutput.n250 CSoutput.n213 2.2505
R16177 CSoutput.n219 CSoutput.n213 2.2505
R16178 CSoutput.n264 CSoutput.n213 2.2505
R16179 CSoutput.n264 CSoutput.n217 2.2505
R16180 CSoutput.n164 CSoutput.n144 2.2505
R16181 CSoutput.n159 CSoutput.n144 2.2505
R16182 CSoutput.n157 CSoutput.n144 2.2505
R16183 CSoutput.n156 CSoutput.n144 2.2505
R16184 CSoutput.n285 CSoutput.n144 2.2505
R16185 CSoutput.n283 CSoutput.n144 2.2505
R16186 CSoutput.n281 CSoutput.n144 2.2505
R16187 CSoutput.n167 CSoutput.n144 2.2505
R16188 CSoutput.n166 CSoutput.n144 2.2505
R16189 CSoutput.n170 CSoutput.n144 2.2505
R16190 CSoutput.n169 CSoutput.n144 2.2505
R16191 CSoutput.n152 CSoutput.n144 2.2505
R16192 CSoutput.n288 CSoutput.n144 2.2505
R16193 CSoutput.n288 CSoutput.n287 2.2505
R16194 CSoutput.n206 CSoutput.n199 2.25024
R16195 CSoutput.n206 CSoutput.n192 2.25024
R16196 CSoutput.n274 CSoutput.n206 2.25024
R16197 CSoutput.n206 CSoutput.n202 2.25024
R16198 CSoutput.n206 CSoutput.n205 2.25024
R16199 CSoutput.n206 CSoutput.n173 2.25024
R16200 CSoutput.n256 CSoutput.n253 2.25024
R16201 CSoutput.n256 CSoutput.n252 2.25024
R16202 CSoutput.n256 CSoutput.n251 2.25024
R16203 CSoutput.n256 CSoutput.n218 2.25024
R16204 CSoutput.n256 CSoutput.n255 2.25024
R16205 CSoutput.n257 CSoutput.n256 2.25024
R16206 CSoutput.n172 CSoutput.n165 2.25024
R16207 CSoutput.n172 CSoutput.n158 2.25024
R16208 CSoutput.n284 CSoutput.n172 2.25024
R16209 CSoutput.n172 CSoutput.n168 2.25024
R16210 CSoutput.n172 CSoutput.n171 2.25024
R16211 CSoutput.n172 CSoutput.n139 2.25024
R16212 CSoutput.n273 CSoutput.n183 1.50111
R16213 CSoutput.n221 CSoutput.n207 1.50111
R16214 CSoutput.n283 CSoutput.n149 1.50111
R16215 CSoutput.n229 CSoutput.n228 1.501
R16216 CSoutput.n236 CSoutput.n235 1.501
R16217 CSoutput.n263 CSoutput.n262 1.501
R16218 CSoutput.n277 CSoutput.n188 1.12536
R16219 CSoutput.n277 CSoutput.n189 1.12536
R16220 CSoutput.n277 CSoutput.n276 1.12536
R16221 CSoutput.n237 CSoutput.n217 1.12536
R16222 CSoutput.n243 CSoutput.n217 1.12536
R16223 CSoutput.n245 CSoutput.n217 1.12536
R16224 CSoutput.n287 CSoutput.n154 1.12536
R16225 CSoutput.n287 CSoutput.n155 1.12536
R16226 CSoutput.n287 CSoutput.n286 1.12536
R16227 CSoutput.n277 CSoutput.n184 1.12536
R16228 CSoutput.n277 CSoutput.n185 1.12536
R16229 CSoutput.n277 CSoutput.n187 1.12536
R16230 CSoutput.n267 CSoutput.n217 1.12536
R16231 CSoutput.n247 CSoutput.n217 1.12536
R16232 CSoutput.n249 CSoutput.n217 1.12536
R16233 CSoutput.n287 CSoutput.n150 1.12536
R16234 CSoutput.n287 CSoutput.n151 1.12536
R16235 CSoutput.n287 CSoutput.n153 1.12536
R16236 CSoutput.n31 CSoutput.n30 0.669944
R16237 CSoutput.n62 CSoutput.n61 0.669944
R16238 CSoutput.n376 CSoutput.n374 0.573776
R16239 CSoutput.n378 CSoutput.n376 0.573776
R16240 CSoutput.n380 CSoutput.n378 0.573776
R16241 CSoutput.n382 CSoutput.n380 0.573776
R16242 CSoutput.n364 CSoutput.n362 0.573776
R16243 CSoutput.n366 CSoutput.n364 0.573776
R16244 CSoutput.n368 CSoutput.n366 0.573776
R16245 CSoutput.n370 CSoutput.n368 0.573776
R16246 CSoutput.n353 CSoutput.n351 0.573776
R16247 CSoutput.n355 CSoutput.n353 0.573776
R16248 CSoutput.n357 CSoutput.n355 0.573776
R16249 CSoutput.n359 CSoutput.n357 0.573776
R16250 CSoutput.n418 CSoutput.n416 0.573776
R16251 CSoutput.n416 CSoutput.n414 0.573776
R16252 CSoutput.n414 CSoutput.n412 0.573776
R16253 CSoutput.n412 CSoutput.n410 0.573776
R16254 CSoutput.n406 CSoutput.n404 0.573776
R16255 CSoutput.n404 CSoutput.n402 0.573776
R16256 CSoutput.n402 CSoutput.n400 0.573776
R16257 CSoutput.n400 CSoutput.n398 0.573776
R16258 CSoutput.n395 CSoutput.n393 0.573776
R16259 CSoutput.n393 CSoutput.n391 0.573776
R16260 CSoutput.n391 CSoutput.n389 0.573776
R16261 CSoutput.n389 CSoutput.n387 0.573776
R16262 CSoutput.n421 CSoutput.n288 0.534303
R16263 CSoutput.n332 CSoutput.n330 0.358259
R16264 CSoutput.n334 CSoutput.n332 0.358259
R16265 CSoutput.n336 CSoutput.n334 0.358259
R16266 CSoutput.n338 CSoutput.n336 0.358259
R16267 CSoutput.n340 CSoutput.n338 0.358259
R16268 CSoutput.n342 CSoutput.n340 0.358259
R16269 CSoutput.n344 CSoutput.n342 0.358259
R16270 CSoutput.n346 CSoutput.n344 0.358259
R16271 CSoutput.n312 CSoutput.n310 0.358259
R16272 CSoutput.n314 CSoutput.n312 0.358259
R16273 CSoutput.n316 CSoutput.n314 0.358259
R16274 CSoutput.n318 CSoutput.n316 0.358259
R16275 CSoutput.n320 CSoutput.n318 0.358259
R16276 CSoutput.n322 CSoutput.n320 0.358259
R16277 CSoutput.n324 CSoutput.n322 0.358259
R16278 CSoutput.n326 CSoutput.n324 0.358259
R16279 CSoutput.n293 CSoutput.n291 0.358259
R16280 CSoutput.n295 CSoutput.n293 0.358259
R16281 CSoutput.n297 CSoutput.n295 0.358259
R16282 CSoutput.n299 CSoutput.n297 0.358259
R16283 CSoutput.n301 CSoutput.n299 0.358259
R16284 CSoutput.n303 CSoutput.n301 0.358259
R16285 CSoutput.n305 CSoutput.n303 0.358259
R16286 CSoutput.n307 CSoutput.n305 0.358259
R16287 CSoutput.n136 CSoutput.n134 0.358259
R16288 CSoutput.n134 CSoutput.n132 0.358259
R16289 CSoutput.n132 CSoutput.n130 0.358259
R16290 CSoutput.n130 CSoutput.n128 0.358259
R16291 CSoutput.n128 CSoutput.n126 0.358259
R16292 CSoutput.n126 CSoutput.n124 0.358259
R16293 CSoutput.n124 CSoutput.n122 0.358259
R16294 CSoutput.n122 CSoutput.n120 0.358259
R16295 CSoutput.n116 CSoutput.n114 0.358259
R16296 CSoutput.n114 CSoutput.n112 0.358259
R16297 CSoutput.n112 CSoutput.n110 0.358259
R16298 CSoutput.n110 CSoutput.n108 0.358259
R16299 CSoutput.n108 CSoutput.n106 0.358259
R16300 CSoutput.n106 CSoutput.n104 0.358259
R16301 CSoutput.n104 CSoutput.n102 0.358259
R16302 CSoutput.n102 CSoutput.n100 0.358259
R16303 CSoutput.n97 CSoutput.n95 0.358259
R16304 CSoutput.n95 CSoutput.n93 0.358259
R16305 CSoutput.n93 CSoutput.n91 0.358259
R16306 CSoutput.n91 CSoutput.n89 0.358259
R16307 CSoutput.n89 CSoutput.n87 0.358259
R16308 CSoutput.n87 CSoutput.n85 0.358259
R16309 CSoutput.n85 CSoutput.n83 0.358259
R16310 CSoutput.n83 CSoutput.n81 0.358259
R16311 CSoutput.n21 CSoutput.n20 0.169105
R16312 CSoutput.n21 CSoutput.n16 0.169105
R16313 CSoutput.n26 CSoutput.n16 0.169105
R16314 CSoutput.n27 CSoutput.n26 0.169105
R16315 CSoutput.n27 CSoutput.n14 0.169105
R16316 CSoutput.n32 CSoutput.n14 0.169105
R16317 CSoutput.n33 CSoutput.n32 0.169105
R16318 CSoutput.n34 CSoutput.n33 0.169105
R16319 CSoutput.n34 CSoutput.n12 0.169105
R16320 CSoutput.n39 CSoutput.n12 0.169105
R16321 CSoutput.n40 CSoutput.n39 0.169105
R16322 CSoutput.n40 CSoutput.n10 0.169105
R16323 CSoutput.n45 CSoutput.n10 0.169105
R16324 CSoutput.n46 CSoutput.n45 0.169105
R16325 CSoutput.n47 CSoutput.n46 0.169105
R16326 CSoutput.n47 CSoutput.n8 0.169105
R16327 CSoutput.n52 CSoutput.n8 0.169105
R16328 CSoutput.n53 CSoutput.n52 0.169105
R16329 CSoutput.n53 CSoutput.n6 0.169105
R16330 CSoutput.n58 CSoutput.n6 0.169105
R16331 CSoutput.n59 CSoutput.n58 0.169105
R16332 CSoutput.n60 CSoutput.n59 0.169105
R16333 CSoutput.n60 CSoutput.n4 0.169105
R16334 CSoutput.n66 CSoutput.n4 0.169105
R16335 CSoutput.n67 CSoutput.n66 0.169105
R16336 CSoutput.n68 CSoutput.n67 0.169105
R16337 CSoutput.n68 CSoutput.n2 0.169105
R16338 CSoutput.n73 CSoutput.n2 0.169105
R16339 CSoutput.n74 CSoutput.n73 0.169105
R16340 CSoutput.n74 CSoutput.n0 0.169105
R16341 CSoutput.n78 CSoutput.n0 0.169105
R16342 CSoutput.n231 CSoutput.n230 0.0910737
R16343 CSoutput.n282 CSoutput.n279 0.0723685
R16344 CSoutput.n236 CSoutput.n231 0.0522944
R16345 CSoutput.n279 CSoutput.n278 0.0499135
R16346 CSoutput.n230 CSoutput.n229 0.0499135
R16347 CSoutput.n264 CSoutput.n263 0.0464294
R16348 CSoutput.n272 CSoutput.n269 0.0391444
R16349 CSoutput.n231 CSoutput.t211 0.023435
R16350 CSoutput.n279 CSoutput.t195 0.02262
R16351 CSoutput.n230 CSoutput.t205 0.02262
R16352 CSoutput CSoutput.n421 0.0052
R16353 CSoutput.n201 CSoutput.n184 0.00365111
R16354 CSoutput.n204 CSoutput.n185 0.00365111
R16355 CSoutput.n187 CSoutput.n186 0.00365111
R16356 CSoutput.n229 CSoutput.n188 0.00365111
R16357 CSoutput.n193 CSoutput.n189 0.00365111
R16358 CSoutput.n276 CSoutput.n190 0.00365111
R16359 CSoutput.n267 CSoutput.n266 0.00365111
R16360 CSoutput.n247 CSoutput.n220 0.00365111
R16361 CSoutput.n249 CSoutput.n219 0.00365111
R16362 CSoutput.n237 CSoutput.n236 0.00365111
R16363 CSoutput.n243 CSoutput.n223 0.00365111
R16364 CSoutput.n245 CSoutput.n222 0.00365111
R16365 CSoutput.n167 CSoutput.n150 0.00365111
R16366 CSoutput.n170 CSoutput.n151 0.00365111
R16367 CSoutput.n153 CSoutput.n152 0.00365111
R16368 CSoutput.n263 CSoutput.n154 0.00365111
R16369 CSoutput.n159 CSoutput.n155 0.00365111
R16370 CSoutput.n286 CSoutput.n156 0.00365111
R16371 CSoutput.n198 CSoutput.n188 0.00340054
R16372 CSoutput.n191 CSoutput.n189 0.00340054
R16373 CSoutput.n276 CSoutput.n275 0.00340054
R16374 CSoutput.n271 CSoutput.n184 0.00340054
R16375 CSoutput.n200 CSoutput.n185 0.00340054
R16376 CSoutput.n203 CSoutput.n187 0.00340054
R16377 CSoutput.n242 CSoutput.n237 0.00340054
R16378 CSoutput.n244 CSoutput.n243 0.00340054
R16379 CSoutput.n246 CSoutput.n245 0.00340054
R16380 CSoutput.n268 CSoutput.n267 0.00340054
R16381 CSoutput.n248 CSoutput.n247 0.00340054
R16382 CSoutput.n250 CSoutput.n249 0.00340054
R16383 CSoutput.n164 CSoutput.n154 0.00340054
R16384 CSoutput.n157 CSoutput.n155 0.00340054
R16385 CSoutput.n286 CSoutput.n285 0.00340054
R16386 CSoutput.n281 CSoutput.n150 0.00340054
R16387 CSoutput.n166 CSoutput.n151 0.00340054
R16388 CSoutput.n169 CSoutput.n153 0.00340054
R16389 CSoutput.n199 CSoutput.n193 0.00252698
R16390 CSoutput.n192 CSoutput.n190 0.00252698
R16391 CSoutput.n274 CSoutput.n273 0.00252698
R16392 CSoutput.n202 CSoutput.n200 0.00252698
R16393 CSoutput.n205 CSoutput.n203 0.00252698
R16394 CSoutput.n278 CSoutput.n173 0.00252698
R16395 CSoutput.n199 CSoutput.n198 0.00252698
R16396 CSoutput.n192 CSoutput.n191 0.00252698
R16397 CSoutput.n275 CSoutput.n274 0.00252698
R16398 CSoutput.n202 CSoutput.n201 0.00252698
R16399 CSoutput.n205 CSoutput.n204 0.00252698
R16400 CSoutput.n186 CSoutput.n173 0.00252698
R16401 CSoutput.n253 CSoutput.n223 0.00252698
R16402 CSoutput.n252 CSoutput.n222 0.00252698
R16403 CSoutput.n251 CSoutput.n207 0.00252698
R16404 CSoutput.n248 CSoutput.n218 0.00252698
R16405 CSoutput.n255 CSoutput.n250 0.00252698
R16406 CSoutput.n264 CSoutput.n257 0.00252698
R16407 CSoutput.n253 CSoutput.n242 0.00252698
R16408 CSoutput.n252 CSoutput.n244 0.00252698
R16409 CSoutput.n251 CSoutput.n246 0.00252698
R16410 CSoutput.n266 CSoutput.n218 0.00252698
R16411 CSoutput.n255 CSoutput.n220 0.00252698
R16412 CSoutput.n257 CSoutput.n219 0.00252698
R16413 CSoutput.n165 CSoutput.n159 0.00252698
R16414 CSoutput.n158 CSoutput.n156 0.00252698
R16415 CSoutput.n284 CSoutput.n283 0.00252698
R16416 CSoutput.n168 CSoutput.n166 0.00252698
R16417 CSoutput.n171 CSoutput.n169 0.00252698
R16418 CSoutput.n288 CSoutput.n139 0.00252698
R16419 CSoutput.n165 CSoutput.n164 0.00252698
R16420 CSoutput.n158 CSoutput.n157 0.00252698
R16421 CSoutput.n285 CSoutput.n284 0.00252698
R16422 CSoutput.n168 CSoutput.n167 0.00252698
R16423 CSoutput.n171 CSoutput.n170 0.00252698
R16424 CSoutput.n152 CSoutput.n139 0.00252698
R16425 CSoutput.n273 CSoutput.n272 0.0020275
R16426 CSoutput.n272 CSoutput.n271 0.0020275
R16427 CSoutput.n269 CSoutput.n207 0.0020275
R16428 CSoutput.n269 CSoutput.n268 0.0020275
R16429 CSoutput.n283 CSoutput.n282 0.0020275
R16430 CSoutput.n282 CSoutput.n281 0.0020275
R16431 CSoutput.n183 CSoutput.n182 0.00166668
R16432 CSoutput.n265 CSoutput.n221 0.00166668
R16433 CSoutput.n149 CSoutput.n148 0.00166668
R16434 CSoutput.n287 CSoutput.n149 0.00133328
R16435 CSoutput.n221 CSoutput.n217 0.00133328
R16436 CSoutput.n277 CSoutput.n183 0.00133328
R16437 CSoutput.n280 CSoutput.n172 0.001
R16438 CSoutput.n258 CSoutput.n172 0.001
R16439 CSoutput.n160 CSoutput.n140 0.001
R16440 CSoutput.n259 CSoutput.n140 0.001
R16441 CSoutput.n161 CSoutput.n141 0.001
R16442 CSoutput.n260 CSoutput.n141 0.001
R16443 CSoutput.n162 CSoutput.n142 0.001
R16444 CSoutput.n261 CSoutput.n142 0.001
R16445 CSoutput.n163 CSoutput.n143 0.001
R16446 CSoutput.n262 CSoutput.n143 0.001
R16447 CSoutput.n256 CSoutput.n208 0.001
R16448 CSoutput.n256 CSoutput.n254 0.001
R16449 CSoutput.n238 CSoutput.n209 0.001
R16450 CSoutput.n232 CSoutput.n209 0.001
R16451 CSoutput.n239 CSoutput.n210 0.001
R16452 CSoutput.n233 CSoutput.n210 0.001
R16453 CSoutput.n240 CSoutput.n211 0.001
R16454 CSoutput.n234 CSoutput.n211 0.001
R16455 CSoutput.n241 CSoutput.n212 0.001
R16456 CSoutput.n235 CSoutput.n212 0.001
R16457 CSoutput.n270 CSoutput.n206 0.001
R16458 CSoutput.n224 CSoutput.n206 0.001
R16459 CSoutput.n194 CSoutput.n174 0.001
R16460 CSoutput.n225 CSoutput.n174 0.001
R16461 CSoutput.n195 CSoutput.n175 0.001
R16462 CSoutput.n226 CSoutput.n175 0.001
R16463 CSoutput.n196 CSoutput.n176 0.001
R16464 CSoutput.n227 CSoutput.n176 0.001
R16465 CSoutput.n197 CSoutput.n177 0.001
R16466 CSoutput.n228 CSoutput.n177 0.001
R16467 CSoutput.n228 CSoutput.n178 0.001
R16468 CSoutput.n227 CSoutput.n179 0.001
R16469 CSoutput.n226 CSoutput.n180 0.001
R16470 CSoutput.n225 CSoutput.t198 0.001
R16471 CSoutput.n224 CSoutput.n181 0.001
R16472 CSoutput.n197 CSoutput.n179 0.001
R16473 CSoutput.n196 CSoutput.n180 0.001
R16474 CSoutput.n195 CSoutput.t198 0.001
R16475 CSoutput.n194 CSoutput.n181 0.001
R16476 CSoutput.n270 CSoutput.n182 0.001
R16477 CSoutput.n235 CSoutput.n213 0.001
R16478 CSoutput.n234 CSoutput.n214 0.001
R16479 CSoutput.n233 CSoutput.n215 0.001
R16480 CSoutput.n232 CSoutput.t206 0.001
R16481 CSoutput.n254 CSoutput.n216 0.001
R16482 CSoutput.n241 CSoutput.n214 0.001
R16483 CSoutput.n240 CSoutput.n215 0.001
R16484 CSoutput.n239 CSoutput.t206 0.001
R16485 CSoutput.n238 CSoutput.n216 0.001
R16486 CSoutput.n265 CSoutput.n208 0.001
R16487 CSoutput.n262 CSoutput.n144 0.001
R16488 CSoutput.n261 CSoutput.n145 0.001
R16489 CSoutput.n260 CSoutput.n146 0.001
R16490 CSoutput.n259 CSoutput.t209 0.001
R16491 CSoutput.n258 CSoutput.n147 0.001
R16492 CSoutput.n163 CSoutput.n145 0.001
R16493 CSoutput.n162 CSoutput.n146 0.001
R16494 CSoutput.n161 CSoutput.t209 0.001
R16495 CSoutput.n160 CSoutput.n147 0.001
R16496 CSoutput.n280 CSoutput.n148 0.001
R16497 a_n2982_13878.n8 a_n2982_13878.t102 538.698
R16498 a_n2982_13878.n104 a_n2982_13878.t79 512.366
R16499 a_n2982_13878.n103 a_n2982_13878.t84 512.366
R16500 a_n2982_13878.n95 a_n2982_13878.t72 512.366
R16501 a_n2982_13878.n102 a_n2982_13878.t89 512.366
R16502 a_n2982_13878.n101 a_n2982_13878.t98 512.366
R16503 a_n2982_13878.n96 a_n2982_13878.t99 512.366
R16504 a_n2982_13878.n100 a_n2982_13878.t66 512.366
R16505 a_n2982_13878.n99 a_n2982_13878.t81 512.366
R16506 a_n2982_13878.n97 a_n2982_13878.t69 512.366
R16507 a_n2982_13878.n98 a_n2982_13878.t76 512.366
R16508 a_n2982_13878.n66 a_n2982_13878.t29 532.5
R16509 a_n2982_13878.n119 a_n2982_13878.t47 512.366
R16510 a_n2982_13878.n118 a_n2982_13878.t49 512.366
R16511 a_n2982_13878.n92 a_n2982_13878.t25 512.366
R16512 a_n2982_13878.n117 a_n2982_13878.t53 512.366
R16513 a_n2982_13878.n116 a_n2982_13878.t13 512.366
R16514 a_n2982_13878.n93 a_n2982_13878.t19 512.366
R16515 a_n2982_13878.n115 a_n2982_13878.t27 512.366
R16516 a_n2982_13878.n114 a_n2982_13878.t55 512.366
R16517 a_n2982_13878.n94 a_n2982_13878.t21 512.366
R16518 a_n2982_13878.n113 a_n2982_13878.t31 512.366
R16519 a_n2982_13878.n26 a_n2982_13878.t41 538.698
R16520 a_n2982_13878.n145 a_n2982_13878.t17 512.366
R16521 a_n2982_13878.n87 a_n2982_13878.t39 512.366
R16522 a_n2982_13878.n146 a_n2982_13878.t11 512.366
R16523 a_n2982_13878.n86 a_n2982_13878.t35 512.366
R16524 a_n2982_13878.n147 a_n2982_13878.t45 512.366
R16525 a_n2982_13878.n148 a_n2982_13878.t15 512.366
R16526 a_n2982_13878.n85 a_n2982_13878.t51 512.366
R16527 a_n2982_13878.n149 a_n2982_13878.t43 512.366
R16528 a_n2982_13878.n84 a_n2982_13878.t23 512.366
R16529 a_n2982_13878.n150 a_n2982_13878.t37 512.366
R16530 a_n2982_13878.n32 a_n2982_13878.t101 538.698
R16531 a_n2982_13878.n139 a_n2982_13878.t70 512.366
R16532 a_n2982_13878.n91 a_n2982_13878.t71 512.366
R16533 a_n2982_13878.n140 a_n2982_13878.t96 512.366
R16534 a_n2982_13878.n90 a_n2982_13878.t97 512.366
R16535 a_n2982_13878.n141 a_n2982_13878.t68 512.366
R16536 a_n2982_13878.n142 a_n2982_13878.t92 512.366
R16537 a_n2982_13878.n89 a_n2982_13878.t93 512.366
R16538 a_n2982_13878.n143 a_n2982_13878.t65 512.366
R16539 a_n2982_13878.n88 a_n2982_13878.t78 512.366
R16540 a_n2982_13878.n144 a_n2982_13878.t88 512.366
R16541 a_n2982_13878.n131 a_n2982_13878.t86 512.366
R16542 a_n2982_13878.n130 a_n2982_13878.t75 512.366
R16543 a_n2982_13878.n129 a_n2982_13878.t64 512.366
R16544 a_n2982_13878.n133 a_n2982_13878.t94 512.366
R16545 a_n2982_13878.n132 a_n2982_13878.t83 512.366
R16546 a_n2982_13878.n128 a_n2982_13878.t82 512.366
R16547 a_n2982_13878.n135 a_n2982_13878.t90 512.366
R16548 a_n2982_13878.n134 a_n2982_13878.t73 512.366
R16549 a_n2982_13878.n127 a_n2982_13878.t74 512.366
R16550 a_n2982_13878.n137 a_n2982_13878.t77 512.366
R16551 a_n2982_13878.n136 a_n2982_13878.t87 512.366
R16552 a_n2982_13878.n126 a_n2982_13878.t103 512.366
R16553 a_n2982_13878.n82 a_n2982_13878.n3 70.5844
R16554 a_n2982_13878.n34 a_n2982_13878.n33 44.7878
R16555 a_n2982_13878.n22 a_n2982_13878.n56 70.5844
R16556 a_n2982_13878.n28 a_n2982_13878.n48 70.5844
R16557 a_n2982_13878.n47 a_n2982_13878.n28 70.1674
R16558 a_n2982_13878.n47 a_n2982_13878.n88 20.9683
R16559 a_n2982_13878.n27 a_n2982_13878.n46 74.73
R16560 a_n2982_13878.n143 a_n2982_13878.n46 11.843
R16561 a_n2982_13878.n45 a_n2982_13878.n27 80.4688
R16562 a_n2982_13878.n45 a_n2982_13878.n89 0.365327
R16563 a_n2982_13878.n29 a_n2982_13878.n44 75.0448
R16564 a_n2982_13878.n43 a_n2982_13878.n29 70.1674
R16565 a_n2982_13878.n43 a_n2982_13878.n90 20.9683
R16566 a_n2982_13878.n30 a_n2982_13878.n42 70.3058
R16567 a_n2982_13878.n140 a_n2982_13878.n42 20.6913
R16568 a_n2982_13878.n41 a_n2982_13878.n30 75.3623
R16569 a_n2982_13878.n41 a_n2982_13878.n91 10.5784
R16570 a_n2982_13878.n32 a_n2982_13878.n31 44.7878
R16571 a_n2982_13878.n55 a_n2982_13878.n22 70.1674
R16572 a_n2982_13878.n55 a_n2982_13878.n84 20.9683
R16573 a_n2982_13878.n21 a_n2982_13878.n54 74.73
R16574 a_n2982_13878.n149 a_n2982_13878.n54 11.843
R16575 a_n2982_13878.n53 a_n2982_13878.n21 80.4688
R16576 a_n2982_13878.n53 a_n2982_13878.n85 0.365327
R16577 a_n2982_13878.n23 a_n2982_13878.n52 75.0448
R16578 a_n2982_13878.n51 a_n2982_13878.n23 70.1674
R16579 a_n2982_13878.n51 a_n2982_13878.n86 20.9683
R16580 a_n2982_13878.n24 a_n2982_13878.n50 70.3058
R16581 a_n2982_13878.n146 a_n2982_13878.n50 20.6913
R16582 a_n2982_13878.n49 a_n2982_13878.n24 75.3623
R16583 a_n2982_13878.n49 a_n2982_13878.n87 10.5784
R16584 a_n2982_13878.n26 a_n2982_13878.n25 44.7878
R16585 a_n2982_13878.n13 a_n2982_13878.n65 70.1674
R16586 a_n2982_13878.n15 a_n2982_13878.n62 70.1674
R16587 a_n2982_13878.n17 a_n2982_13878.n60 70.1674
R16588 a_n2982_13878.n19 a_n2982_13878.n58 70.1674
R16589 a_n2982_13878.n58 a_n2982_13878.n126 20.9683
R16590 a_n2982_13878.n57 a_n2982_13878.n20 75.0448
R16591 a_n2982_13878.n136 a_n2982_13878.n57 11.2134
R16592 a_n2982_13878.n20 a_n2982_13878.n137 161.3
R16593 a_n2982_13878.n60 a_n2982_13878.n127 20.9683
R16594 a_n2982_13878.n59 a_n2982_13878.n18 75.0448
R16595 a_n2982_13878.n134 a_n2982_13878.n59 11.2134
R16596 a_n2982_13878.n18 a_n2982_13878.n135 161.3
R16597 a_n2982_13878.n62 a_n2982_13878.n128 20.9683
R16598 a_n2982_13878.n61 a_n2982_13878.n16 75.0448
R16599 a_n2982_13878.n132 a_n2982_13878.n61 11.2134
R16600 a_n2982_13878.n16 a_n2982_13878.n133 161.3
R16601 a_n2982_13878.n65 a_n2982_13878.n129 20.9683
R16602 a_n2982_13878.n63 a_n2982_13878.n14 75.0448
R16603 a_n2982_13878.n130 a_n2982_13878.n63 11.2134
R16604 a_n2982_13878.n14 a_n2982_13878.n131 161.3
R16605 a_n2982_13878.n34 a_n2982_13878.n113 14.1668
R16606 a_n2982_13878.n74 a_n2982_13878.n73 75.3623
R16607 a_n2982_13878.n72 a_n2982_13878.n9 70.3058
R16608 a_n2982_13878.n9 a_n2982_13878.n71 70.1674
R16609 a_n2982_13878.n71 a_n2982_13878.n93 20.9683
R16610 a_n2982_13878.n70 a_n2982_13878.n10 75.0448
R16611 a_n2982_13878.n116 a_n2982_13878.n70 11.2134
R16612 a_n2982_13878.n69 a_n2982_13878.n10 80.4688
R16613 a_n2982_13878.n12 a_n2982_13878.n68 74.73
R16614 a_n2982_13878.n67 a_n2982_13878.n12 70.1674
R16615 a_n2982_13878.n119 a_n2982_13878.n67 20.9683
R16616 a_n2982_13878.n11 a_n2982_13878.n66 70.5844
R16617 a_n2982_13878.n3 a_n2982_13878.n81 70.1674
R16618 a_n2982_13878.n81 a_n2982_13878.n97 20.9683
R16619 a_n2982_13878.n80 a_n2982_13878.n4 74.73
R16620 a_n2982_13878.n99 a_n2982_13878.n80 11.843
R16621 a_n2982_13878.n79 a_n2982_13878.n4 80.4688
R16622 a_n2982_13878.n79 a_n2982_13878.n100 0.365327
R16623 a_n2982_13878.n5 a_n2982_13878.n78 75.0448
R16624 a_n2982_13878.n77 a_n2982_13878.n5 70.1674
R16625 a_n2982_13878.n102 a_n2982_13878.n77 20.9683
R16626 a_n2982_13878.n7 a_n2982_13878.n76 70.3058
R16627 a_n2982_13878.n76 a_n2982_13878.n95 20.6913
R16628 a_n2982_13878.n75 a_n2982_13878.n7 75.3623
R16629 a_n2982_13878.n103 a_n2982_13878.n75 10.5784
R16630 a_n2982_13878.n6 a_n2982_13878.n8 44.7878
R16631 a_n2982_13878.n1 a_n2982_13878.n111 81.3764
R16632 a_n2982_13878.n2 a_n2982_13878.n107 81.3764
R16633 a_n2982_13878.n2 a_n2982_13878.n105 81.3764
R16634 a_n2982_13878.n1 a_n2982_13878.n112 80.9324
R16635 a_n2982_13878.n1 a_n2982_13878.n110 80.9324
R16636 a_n2982_13878.n0 a_n2982_13878.n109 80.9324
R16637 a_n2982_13878.n2 a_n2982_13878.n108 80.9324
R16638 a_n2982_13878.n2 a_n2982_13878.n106 80.9324
R16639 a_n2982_13878.n39 a_n2982_13878.t42 74.6477
R16640 a_n2982_13878.n37 a_n2982_13878.t34 74.6477
R16641 a_n2982_13878.n36 a_n2982_13878.t30 74.2899
R16642 a_n2982_13878.n40 a_n2982_13878.t58 74.2897
R16643 a_n2982_13878.n40 a_n2982_13878.n152 70.6783
R16644 a_n2982_13878.n38 a_n2982_13878.n153 70.6783
R16645 a_n2982_13878.n38 a_n2982_13878.n154 70.6783
R16646 a_n2982_13878.n39 a_n2982_13878.n83 70.6783
R16647 a_n2982_13878.n37 a_n2982_13878.n120 70.6783
R16648 a_n2982_13878.n37 a_n2982_13878.n121 70.6783
R16649 a_n2982_13878.n35 a_n2982_13878.n122 70.6783
R16650 a_n2982_13878.n35 a_n2982_13878.n123 70.6783
R16651 a_n2982_13878.n36 a_n2982_13878.n124 70.6783
R16652 a_n2982_13878.n155 a_n2982_13878.n39 70.6782
R16653 a_n2982_13878.n104 a_n2982_13878.n103 48.2005
R16654 a_n2982_13878.n77 a_n2982_13878.n101 20.9683
R16655 a_n2982_13878.n100 a_n2982_13878.n96 48.2005
R16656 a_n2982_13878.n98 a_n2982_13878.n81 20.9683
R16657 a_n2982_13878.n67 a_n2982_13878.n118 20.9683
R16658 a_n2982_13878.n117 a_n2982_13878.n116 48.2005
R16659 a_n2982_13878.n115 a_n2982_13878.n71 20.9683
R16660 a_n2982_13878.n113 a_n2982_13878.n94 48.2005
R16661 a_n2982_13878.n145 a_n2982_13878.n87 48.2005
R16662 a_n2982_13878.n147 a_n2982_13878.n51 20.9683
R16663 a_n2982_13878.n148 a_n2982_13878.n85 48.2005
R16664 a_n2982_13878.n150 a_n2982_13878.n55 20.9683
R16665 a_n2982_13878.n139 a_n2982_13878.n91 48.2005
R16666 a_n2982_13878.n141 a_n2982_13878.n43 20.9683
R16667 a_n2982_13878.n142 a_n2982_13878.n89 48.2005
R16668 a_n2982_13878.n144 a_n2982_13878.n47 20.9683
R16669 a_n2982_13878.n131 a_n2982_13878.n130 48.2005
R16670 a_n2982_13878.t91 a_n2982_13878.n65 533.335
R16671 a_n2982_13878.n133 a_n2982_13878.n132 48.2005
R16672 a_n2982_13878.t100 a_n2982_13878.n62 533.335
R16673 a_n2982_13878.n135 a_n2982_13878.n134 48.2005
R16674 a_n2982_13878.t85 a_n2982_13878.n60 533.335
R16675 a_n2982_13878.n137 a_n2982_13878.n136 48.2005
R16676 a_n2982_13878.t80 a_n2982_13878.n58 533.335
R16677 a_n2982_13878.n102 a_n2982_13878.n76 21.4216
R16678 a_n2982_13878.n69 a_n2982_13878.n92 47.835
R16679 a_n2982_13878.n72 a_n2982_13878.n114 20.6913
R16680 a_n2982_13878.n86 a_n2982_13878.n50 21.4216
R16681 a_n2982_13878.n90 a_n2982_13878.n42 21.4216
R16682 a_n2982_13878.n82 a_n2982_13878.t95 532.5
R16683 a_n2982_13878.t57 a_n2982_13878.n56 532.5
R16684 a_n2982_13878.t67 a_n2982_13878.n48 532.5
R16685 a_n2982_13878.n80 a_n2982_13878.n97 34.4824
R16686 a_n2982_13878.n68 a_n2982_13878.n92 11.843
R16687 a_n2982_13878.n114 a_n2982_13878.n73 36.139
R16688 a_n2982_13878.n84 a_n2982_13878.n54 34.4824
R16689 a_n2982_13878.n88 a_n2982_13878.n46 34.4824
R16690 a_n2982_13878.n101 a_n2982_13878.n78 35.3134
R16691 a_n2982_13878.n78 a_n2982_13878.n96 11.2134
R16692 a_n2982_13878.n70 a_n2982_13878.n93 35.3134
R16693 a_n2982_13878.n52 a_n2982_13878.n147 35.3134
R16694 a_n2982_13878.n148 a_n2982_13878.n52 11.2134
R16695 a_n2982_13878.n44 a_n2982_13878.n141 35.3134
R16696 a_n2982_13878.n142 a_n2982_13878.n44 11.2134
R16697 a_n2982_13878.n63 a_n2982_13878.n129 35.3134
R16698 a_n2982_13878.n61 a_n2982_13878.n128 35.3134
R16699 a_n2982_13878.n59 a_n2982_13878.n127 35.3134
R16700 a_n2982_13878.n57 a_n2982_13878.n126 35.3134
R16701 a_n2982_13878.n33 a_n2982_13878.n1 23.891
R16702 a_n2982_13878.n75 a_n2982_13878.n95 36.139
R16703 a_n2982_13878.n118 a_n2982_13878.n68 34.4824
R16704 a_n2982_13878.n73 a_n2982_13878.n94 10.5784
R16705 a_n2982_13878.n146 a_n2982_13878.n49 36.139
R16706 a_n2982_13878.n140 a_n2982_13878.n41 36.139
R16707 a_n2982_13878.n31 a_n2982_13878.n138 13.9285
R16708 a_n2982_13878.n3 a_n2982_13878.n64 13.724
R16709 a_n2982_13878.n125 a_n2982_13878.n11 12.4191
R16710 a_n2982_13878.n13 a_n2982_13878.n64 11.2486
R16711 a_n2982_13878.n138 a_n2982_13878.n20 11.2486
R16712 a_n2982_13878.n40 a_n2982_13878.n151 10.5745
R16713 a_n2982_13878.n151 a_n2982_13878.n22 8.58383
R16714 a_n2982_13878.n125 a_n2982_13878.n36 6.7311
R16715 a_n2982_13878.n151 a_n2982_13878.n64 5.3452
R16716 a_n2982_13878.n25 a_n2982_13878.n28 3.94368
R16717 a_n2982_13878.n33 a_n2982_13878.n6 3.7202
R16718 a_n2982_13878.n152 a_n2982_13878.t24 3.61217
R16719 a_n2982_13878.n152 a_n2982_13878.t38 3.61217
R16720 a_n2982_13878.n153 a_n2982_13878.t52 3.61217
R16721 a_n2982_13878.n153 a_n2982_13878.t44 3.61217
R16722 a_n2982_13878.n154 a_n2982_13878.t46 3.61217
R16723 a_n2982_13878.n154 a_n2982_13878.t16 3.61217
R16724 a_n2982_13878.n83 a_n2982_13878.t18 3.61217
R16725 a_n2982_13878.n83 a_n2982_13878.t40 3.61217
R16726 a_n2982_13878.n120 a_n2982_13878.t22 3.61217
R16727 a_n2982_13878.n120 a_n2982_13878.t32 3.61217
R16728 a_n2982_13878.n121 a_n2982_13878.t28 3.61217
R16729 a_n2982_13878.n121 a_n2982_13878.t56 3.61217
R16730 a_n2982_13878.n122 a_n2982_13878.t14 3.61217
R16731 a_n2982_13878.n122 a_n2982_13878.t20 3.61217
R16732 a_n2982_13878.n123 a_n2982_13878.t26 3.61217
R16733 a_n2982_13878.n123 a_n2982_13878.t54 3.61217
R16734 a_n2982_13878.n124 a_n2982_13878.t48 3.61217
R16735 a_n2982_13878.n124 a_n2982_13878.t50 3.61217
R16736 a_n2982_13878.t12 a_n2982_13878.n155 3.61217
R16737 a_n2982_13878.n155 a_n2982_13878.t36 3.61217
R16738 a_n2982_13878.n111 a_n2982_13878.t62 2.82907
R16739 a_n2982_13878.n111 a_n2982_13878.t3 2.82907
R16740 a_n2982_13878.n112 a_n2982_13878.t5 2.82907
R16741 a_n2982_13878.n112 a_n2982_13878.t61 2.82907
R16742 a_n2982_13878.n110 a_n2982_13878.t60 2.82907
R16743 a_n2982_13878.n110 a_n2982_13878.t63 2.82907
R16744 a_n2982_13878.n109 a_n2982_13878.t7 2.82907
R16745 a_n2982_13878.n109 a_n2982_13878.t59 2.82907
R16746 a_n2982_13878.n107 a_n2982_13878.t10 2.82907
R16747 a_n2982_13878.n107 a_n2982_13878.t1 2.82907
R16748 a_n2982_13878.n108 a_n2982_13878.t8 2.82907
R16749 a_n2982_13878.n108 a_n2982_13878.t0 2.82907
R16750 a_n2982_13878.n106 a_n2982_13878.t9 2.82907
R16751 a_n2982_13878.n106 a_n2982_13878.t4 2.82907
R16752 a_n2982_13878.n105 a_n2982_13878.t2 2.82907
R16753 a_n2982_13878.n105 a_n2982_13878.t6 2.82907
R16754 a_n2982_13878.n8 a_n2982_13878.n104 14.1668
R16755 a_n2982_13878.n98 a_n2982_13878.n82 22.3251
R16756 a_n2982_13878.n66 a_n2982_13878.n119 22.3251
R16757 a_n2982_13878.n34 a_n2982_13878.t33 538.698
R16758 a_n2982_13878.n145 a_n2982_13878.n26 14.1668
R16759 a_n2982_13878.n56 a_n2982_13878.n150 22.3251
R16760 a_n2982_13878.n139 a_n2982_13878.n32 14.1668
R16761 a_n2982_13878.n48 a_n2982_13878.n144 22.3251
R16762 a_n2982_13878.n138 a_n2982_13878.n125 1.30542
R16763 a_n2982_13878.n17 a_n2982_13878.n16 1.04595
R16764 a_n2982_13878.n79 a_n2982_13878.n99 47.835
R16765 a_n2982_13878.n69 a_n2982_13878.n117 0.365327
R16766 a_n2982_13878.n115 a_n2982_13878.n72 21.4216
R16767 a_n2982_13878.n149 a_n2982_13878.n53 47.835
R16768 a_n2982_13878.n143 a_n2982_13878.n45 47.835
R16769 a_n2982_13878.n0 a_n2982_13878.n2 31.7919
R16770 a_n2982_13878.n28 a_n2982_13878.n27 1.13686
R16771 a_n2982_13878.n22 a_n2982_13878.n21 1.13686
R16772 a_n2982_13878.n4 a_n2982_13878.n3 1.13686
R16773 a_n2982_13878.n39 a_n2982_13878.n38 1.07378
R16774 a_n2982_13878.n36 a_n2982_13878.n35 1.07378
R16775 a_n2982_13878.n1 a_n2982_13878.n0 0.888431
R16776 a_n2982_13878.n30 a_n2982_13878.n31 0.758076
R16777 a_n2982_13878.n29 a_n2982_13878.n30 0.758076
R16778 a_n2982_13878.n27 a_n2982_13878.n29 0.758076
R16779 a_n2982_13878.n24 a_n2982_13878.n25 0.758076
R16780 a_n2982_13878.n23 a_n2982_13878.n24 0.758076
R16781 a_n2982_13878.n21 a_n2982_13878.n23 0.758076
R16782 a_n2982_13878.n20 a_n2982_13878.n19 0.758076
R16783 a_n2982_13878.n18 a_n2982_13878.n17 0.758076
R16784 a_n2982_13878.n16 a_n2982_13878.n15 0.758076
R16785 a_n2982_13878.n14 a_n2982_13878.n13 0.758076
R16786 a_n2982_13878.n12 a_n2982_13878.n10 0.758076
R16787 a_n2982_13878.n10 a_n2982_13878.n9 0.758076
R16788 a_n2982_13878.n74 a_n2982_13878.n9 0.758076
R16789 a_n2982_13878.n7 a_n2982_13878.n6 0.758076
R16790 a_n2982_13878.n7 a_n2982_13878.n5 0.758076
R16791 a_n2982_13878.n5 a_n2982_13878.n4 0.758076
R16792 a_n2982_13878.n74 a_n2982_13878.n33 0.754288
R16793 a_n2982_13878.n38 a_n2982_13878.n40 0.716017
R16794 a_n2982_13878.n35 a_n2982_13878.n37 0.716017
R16795 a_n2982_13878.n19 a_n2982_13878.n18 0.67853
R16796 a_n2982_13878.n15 a_n2982_13878.n14 0.67853
R16797 a_n2982_13878.n12 a_n2982_13878.n11 0.568682
R16798 vdd.n327 vdd.n291 756.745
R16799 vdd.n268 vdd.n232 756.745
R16800 vdd.n225 vdd.n189 756.745
R16801 vdd.n166 vdd.n130 756.745
R16802 vdd.n124 vdd.n88 756.745
R16803 vdd.n65 vdd.n29 756.745
R16804 vdd.n2201 vdd.n2165 756.745
R16805 vdd.n2260 vdd.n2224 756.745
R16806 vdd.n2099 vdd.n2063 756.745
R16807 vdd.n2158 vdd.n2122 756.745
R16808 vdd.n1998 vdd.n1962 756.745
R16809 vdd.n2057 vdd.n2021 756.745
R16810 vdd.n1315 vdd.t164 640.208
R16811 vdd.n1010 vdd.t205 640.208
R16812 vdd.n1319 vdd.t202 640.208
R16813 vdd.n1001 vdd.t227 640.208
R16814 vdd.n896 vdd.t189 640.208
R16815 vdd.n2823 vdd.t220 640.208
R16816 vdd.n832 vdd.t182 640.208
R16817 vdd.n2820 vdd.t212 640.208
R16818 vdd.n799 vdd.t160 640.208
R16819 vdd.n1071 vdd.t216 640.208
R16820 vdd.n1772 vdd.t230 592.009
R16821 vdd.n1810 vdd.t223 592.009
R16822 vdd.n1706 vdd.t233 592.009
R16823 vdd.n2362 vdd.t193 592.009
R16824 vdd.n1248 vdd.t168 592.009
R16825 vdd.n1208 vdd.t176 592.009
R16826 vdd.n426 vdd.t199 592.009
R16827 vdd.n440 vdd.t172 592.009
R16828 vdd.n452 vdd.t179 592.009
R16829 vdd.n768 vdd.t196 592.009
R16830 vdd.n3456 vdd.t209 592.009
R16831 vdd.n688 vdd.t185 592.009
R16832 vdd.n328 vdd.n327 585
R16833 vdd.n326 vdd.n293 585
R16834 vdd.n325 vdd.n324 585
R16835 vdd.n296 vdd.n294 585
R16836 vdd.n319 vdd.n318 585
R16837 vdd.n317 vdd.n316 585
R16838 vdd.n300 vdd.n299 585
R16839 vdd.n311 vdd.n310 585
R16840 vdd.n309 vdd.n308 585
R16841 vdd.n304 vdd.n303 585
R16842 vdd.n269 vdd.n268 585
R16843 vdd.n267 vdd.n234 585
R16844 vdd.n266 vdd.n265 585
R16845 vdd.n237 vdd.n235 585
R16846 vdd.n260 vdd.n259 585
R16847 vdd.n258 vdd.n257 585
R16848 vdd.n241 vdd.n240 585
R16849 vdd.n252 vdd.n251 585
R16850 vdd.n250 vdd.n249 585
R16851 vdd.n245 vdd.n244 585
R16852 vdd.n226 vdd.n225 585
R16853 vdd.n224 vdd.n191 585
R16854 vdd.n223 vdd.n222 585
R16855 vdd.n194 vdd.n192 585
R16856 vdd.n217 vdd.n216 585
R16857 vdd.n215 vdd.n214 585
R16858 vdd.n198 vdd.n197 585
R16859 vdd.n209 vdd.n208 585
R16860 vdd.n207 vdd.n206 585
R16861 vdd.n202 vdd.n201 585
R16862 vdd.n167 vdd.n166 585
R16863 vdd.n165 vdd.n132 585
R16864 vdd.n164 vdd.n163 585
R16865 vdd.n135 vdd.n133 585
R16866 vdd.n158 vdd.n157 585
R16867 vdd.n156 vdd.n155 585
R16868 vdd.n139 vdd.n138 585
R16869 vdd.n150 vdd.n149 585
R16870 vdd.n148 vdd.n147 585
R16871 vdd.n143 vdd.n142 585
R16872 vdd.n125 vdd.n124 585
R16873 vdd.n123 vdd.n90 585
R16874 vdd.n122 vdd.n121 585
R16875 vdd.n93 vdd.n91 585
R16876 vdd.n116 vdd.n115 585
R16877 vdd.n114 vdd.n113 585
R16878 vdd.n97 vdd.n96 585
R16879 vdd.n108 vdd.n107 585
R16880 vdd.n106 vdd.n105 585
R16881 vdd.n101 vdd.n100 585
R16882 vdd.n66 vdd.n65 585
R16883 vdd.n64 vdd.n31 585
R16884 vdd.n63 vdd.n62 585
R16885 vdd.n34 vdd.n32 585
R16886 vdd.n57 vdd.n56 585
R16887 vdd.n55 vdd.n54 585
R16888 vdd.n38 vdd.n37 585
R16889 vdd.n49 vdd.n48 585
R16890 vdd.n47 vdd.n46 585
R16891 vdd.n42 vdd.n41 585
R16892 vdd.n2202 vdd.n2201 585
R16893 vdd.n2200 vdd.n2167 585
R16894 vdd.n2199 vdd.n2198 585
R16895 vdd.n2170 vdd.n2168 585
R16896 vdd.n2193 vdd.n2192 585
R16897 vdd.n2191 vdd.n2190 585
R16898 vdd.n2174 vdd.n2173 585
R16899 vdd.n2185 vdd.n2184 585
R16900 vdd.n2183 vdd.n2182 585
R16901 vdd.n2178 vdd.n2177 585
R16902 vdd.n2261 vdd.n2260 585
R16903 vdd.n2259 vdd.n2226 585
R16904 vdd.n2258 vdd.n2257 585
R16905 vdd.n2229 vdd.n2227 585
R16906 vdd.n2252 vdd.n2251 585
R16907 vdd.n2250 vdd.n2249 585
R16908 vdd.n2233 vdd.n2232 585
R16909 vdd.n2244 vdd.n2243 585
R16910 vdd.n2242 vdd.n2241 585
R16911 vdd.n2237 vdd.n2236 585
R16912 vdd.n2100 vdd.n2099 585
R16913 vdd.n2098 vdd.n2065 585
R16914 vdd.n2097 vdd.n2096 585
R16915 vdd.n2068 vdd.n2066 585
R16916 vdd.n2091 vdd.n2090 585
R16917 vdd.n2089 vdd.n2088 585
R16918 vdd.n2072 vdd.n2071 585
R16919 vdd.n2083 vdd.n2082 585
R16920 vdd.n2081 vdd.n2080 585
R16921 vdd.n2076 vdd.n2075 585
R16922 vdd.n2159 vdd.n2158 585
R16923 vdd.n2157 vdd.n2124 585
R16924 vdd.n2156 vdd.n2155 585
R16925 vdd.n2127 vdd.n2125 585
R16926 vdd.n2150 vdd.n2149 585
R16927 vdd.n2148 vdd.n2147 585
R16928 vdd.n2131 vdd.n2130 585
R16929 vdd.n2142 vdd.n2141 585
R16930 vdd.n2140 vdd.n2139 585
R16931 vdd.n2135 vdd.n2134 585
R16932 vdd.n1999 vdd.n1998 585
R16933 vdd.n1997 vdd.n1964 585
R16934 vdd.n1996 vdd.n1995 585
R16935 vdd.n1967 vdd.n1965 585
R16936 vdd.n1990 vdd.n1989 585
R16937 vdd.n1988 vdd.n1987 585
R16938 vdd.n1971 vdd.n1970 585
R16939 vdd.n1982 vdd.n1981 585
R16940 vdd.n1980 vdd.n1979 585
R16941 vdd.n1975 vdd.n1974 585
R16942 vdd.n2058 vdd.n2057 585
R16943 vdd.n2056 vdd.n2023 585
R16944 vdd.n2055 vdd.n2054 585
R16945 vdd.n2026 vdd.n2024 585
R16946 vdd.n2049 vdd.n2048 585
R16947 vdd.n2047 vdd.n2046 585
R16948 vdd.n2030 vdd.n2029 585
R16949 vdd.n2041 vdd.n2040 585
R16950 vdd.n2039 vdd.n2038 585
R16951 vdd.n2034 vdd.n2033 585
R16952 vdd.n3628 vdd.n392 509.269
R16953 vdd.n3624 vdd.n393 509.269
R16954 vdd.n3496 vdd.n685 509.269
R16955 vdd.n3493 vdd.n684 509.269
R16956 vdd.n2357 vdd.n1530 509.269
R16957 vdd.n2360 vdd.n2359 509.269
R16958 vdd.n1679 vdd.n1643 509.269
R16959 vdd.n1875 vdd.n1644 509.269
R16960 vdd.n305 vdd.t36 329.043
R16961 vdd.n246 vdd.t152 329.043
R16962 vdd.n203 vdd.t15 329.043
R16963 vdd.n144 vdd.t141 329.043
R16964 vdd.n102 vdd.t122 329.043
R16965 vdd.n43 vdd.t82 329.043
R16966 vdd.n2179 vdd.t62 329.043
R16967 vdd.n2238 vdd.t105 329.043
R16968 vdd.n2077 vdd.t43 329.043
R16969 vdd.n2136 vdd.t88 329.043
R16970 vdd.n1976 vdd.t83 329.043
R16971 vdd.n2035 vdd.t124 329.043
R16972 vdd.n1772 vdd.t232 319.788
R16973 vdd.n1810 vdd.t226 319.788
R16974 vdd.n1706 vdd.t235 319.788
R16975 vdd.n2362 vdd.t194 319.788
R16976 vdd.n1248 vdd.t170 319.788
R16977 vdd.n1208 vdd.t177 319.788
R16978 vdd.n426 vdd.t200 319.788
R16979 vdd.n440 vdd.t174 319.788
R16980 vdd.n452 vdd.t180 319.788
R16981 vdd.n768 vdd.t198 319.788
R16982 vdd.n3456 vdd.t211 319.788
R16983 vdd.n688 vdd.t188 319.788
R16984 vdd.n1773 vdd.t231 303.69
R16985 vdd.n1811 vdd.t225 303.69
R16986 vdd.n1707 vdd.t234 303.69
R16987 vdd.n2363 vdd.t195 303.69
R16988 vdd.n1249 vdd.t171 303.69
R16989 vdd.n1209 vdd.t178 303.69
R16990 vdd.n427 vdd.t201 303.69
R16991 vdd.n441 vdd.t175 303.69
R16992 vdd.n453 vdd.t181 303.69
R16993 vdd.n769 vdd.t197 303.69
R16994 vdd.n3457 vdd.t210 303.69
R16995 vdd.n689 vdd.t187 303.69
R16996 vdd.n3090 vdd.n960 279.512
R16997 vdd.n3330 vdd.n809 279.512
R16998 vdd.n3267 vdd.n806 279.512
R16999 vdd.n3022 vdd.n3021 279.512
R17000 vdd.n2783 vdd.n998 279.512
R17001 vdd.n2714 vdd.n2713 279.512
R17002 vdd.n1355 vdd.n1354 279.512
R17003 vdd.n2508 vdd.n1138 279.512
R17004 vdd.n3246 vdd.n807 279.512
R17005 vdd.n3333 vdd.n3332 279.512
R17006 vdd.n2895 vdd.n2818 279.512
R17007 vdd.n2826 vdd.n956 279.512
R17008 vdd.n2711 vdd.n1008 279.512
R17009 vdd.n1006 vdd.n980 279.512
R17010 vdd.n1480 vdd.n1175 279.512
R17011 vdd.n1280 vdd.n1133 279.512
R17012 vdd.n2506 vdd.n1141 254.619
R17013 vdd.n3495 vdd.n692 254.619
R17014 vdd.n3248 vdd.n807 185
R17015 vdd.n3331 vdd.n807 185
R17016 vdd.n3250 vdd.n3249 185
R17017 vdd.n3249 vdd.n805 185
R17018 vdd.n3251 vdd.n839 185
R17019 vdd.n3261 vdd.n839 185
R17020 vdd.n3252 vdd.n848 185
R17021 vdd.n848 vdd.n846 185
R17022 vdd.n3254 vdd.n3253 185
R17023 vdd.n3255 vdd.n3254 185
R17024 vdd.n3207 vdd.n847 185
R17025 vdd.n847 vdd.n843 185
R17026 vdd.n3206 vdd.n3205 185
R17027 vdd.n3205 vdd.n3204 185
R17028 vdd.n850 vdd.n849 185
R17029 vdd.n851 vdd.n850 185
R17030 vdd.n3197 vdd.n3196 185
R17031 vdd.n3198 vdd.n3197 185
R17032 vdd.n3195 vdd.n859 185
R17033 vdd.n864 vdd.n859 185
R17034 vdd.n3194 vdd.n3193 185
R17035 vdd.n3193 vdd.n3192 185
R17036 vdd.n861 vdd.n860 185
R17037 vdd.n870 vdd.n861 185
R17038 vdd.n3185 vdd.n3184 185
R17039 vdd.n3186 vdd.n3185 185
R17040 vdd.n3183 vdd.n871 185
R17041 vdd.n877 vdd.n871 185
R17042 vdd.n3182 vdd.n3181 185
R17043 vdd.n3181 vdd.n3180 185
R17044 vdd.n873 vdd.n872 185
R17045 vdd.n874 vdd.n873 185
R17046 vdd.n3173 vdd.n3172 185
R17047 vdd.n3174 vdd.n3173 185
R17048 vdd.n3171 vdd.n884 185
R17049 vdd.n884 vdd.n881 185
R17050 vdd.n3170 vdd.n3169 185
R17051 vdd.n3169 vdd.n3168 185
R17052 vdd.n886 vdd.n885 185
R17053 vdd.n887 vdd.n886 185
R17054 vdd.n3161 vdd.n3160 185
R17055 vdd.n3162 vdd.n3161 185
R17056 vdd.n3159 vdd.n895 185
R17057 vdd.n901 vdd.n895 185
R17058 vdd.n3158 vdd.n3157 185
R17059 vdd.n3157 vdd.n3156 185
R17060 vdd.n3147 vdd.n898 185
R17061 vdd.n908 vdd.n898 185
R17062 vdd.n3149 vdd.n3148 185
R17063 vdd.n3150 vdd.n3149 185
R17064 vdd.n3146 vdd.n909 185
R17065 vdd.n909 vdd.n905 185
R17066 vdd.n3145 vdd.n3144 185
R17067 vdd.n3144 vdd.n3143 185
R17068 vdd.n911 vdd.n910 185
R17069 vdd.n912 vdd.n911 185
R17070 vdd.n3136 vdd.n3135 185
R17071 vdd.n3137 vdd.n3136 185
R17072 vdd.n3134 vdd.n920 185
R17073 vdd.n925 vdd.n920 185
R17074 vdd.n3133 vdd.n3132 185
R17075 vdd.n3132 vdd.n3131 185
R17076 vdd.n922 vdd.n921 185
R17077 vdd.n931 vdd.n922 185
R17078 vdd.n3124 vdd.n3123 185
R17079 vdd.n3125 vdd.n3124 185
R17080 vdd.n3122 vdd.n932 185
R17081 vdd.n2998 vdd.n932 185
R17082 vdd.n3121 vdd.n3120 185
R17083 vdd.n3120 vdd.n3119 185
R17084 vdd.n934 vdd.n933 185
R17085 vdd.n3004 vdd.n934 185
R17086 vdd.n3112 vdd.n3111 185
R17087 vdd.n3113 vdd.n3112 185
R17088 vdd.n3110 vdd.n943 185
R17089 vdd.n943 vdd.n940 185
R17090 vdd.n3109 vdd.n3108 185
R17091 vdd.n3108 vdd.n3107 185
R17092 vdd.n945 vdd.n944 185
R17093 vdd.n946 vdd.n945 185
R17094 vdd.n3100 vdd.n3099 185
R17095 vdd.n3101 vdd.n3100 185
R17096 vdd.n3098 vdd.n954 185
R17097 vdd.n3016 vdd.n954 185
R17098 vdd.n3097 vdd.n3096 185
R17099 vdd.n3096 vdd.n3095 185
R17100 vdd.n956 vdd.n955 185
R17101 vdd.n957 vdd.n956 185
R17102 vdd.n2827 vdd.n2826 185
R17103 vdd.n2829 vdd.n2828 185
R17104 vdd.n2831 vdd.n2830 185
R17105 vdd.n2833 vdd.n2832 185
R17106 vdd.n2835 vdd.n2834 185
R17107 vdd.n2837 vdd.n2836 185
R17108 vdd.n2839 vdd.n2838 185
R17109 vdd.n2841 vdd.n2840 185
R17110 vdd.n2843 vdd.n2842 185
R17111 vdd.n2845 vdd.n2844 185
R17112 vdd.n2847 vdd.n2846 185
R17113 vdd.n2849 vdd.n2848 185
R17114 vdd.n2851 vdd.n2850 185
R17115 vdd.n2853 vdd.n2852 185
R17116 vdd.n2855 vdd.n2854 185
R17117 vdd.n2857 vdd.n2856 185
R17118 vdd.n2859 vdd.n2858 185
R17119 vdd.n2861 vdd.n2860 185
R17120 vdd.n2863 vdd.n2862 185
R17121 vdd.n2865 vdd.n2864 185
R17122 vdd.n2867 vdd.n2866 185
R17123 vdd.n2869 vdd.n2868 185
R17124 vdd.n2871 vdd.n2870 185
R17125 vdd.n2873 vdd.n2872 185
R17126 vdd.n2875 vdd.n2874 185
R17127 vdd.n2877 vdd.n2876 185
R17128 vdd.n2879 vdd.n2878 185
R17129 vdd.n2881 vdd.n2880 185
R17130 vdd.n2883 vdd.n2882 185
R17131 vdd.n2885 vdd.n2884 185
R17132 vdd.n2887 vdd.n2886 185
R17133 vdd.n2889 vdd.n2888 185
R17134 vdd.n2891 vdd.n2890 185
R17135 vdd.n2893 vdd.n2892 185
R17136 vdd.n2894 vdd.n2818 185
R17137 vdd.n3088 vdd.n2818 185
R17138 vdd.n3334 vdd.n3333 185
R17139 vdd.n3335 vdd.n798 185
R17140 vdd.n3337 vdd.n3336 185
R17141 vdd.n3339 vdd.n796 185
R17142 vdd.n3341 vdd.n3340 185
R17143 vdd.n3342 vdd.n795 185
R17144 vdd.n3344 vdd.n3343 185
R17145 vdd.n3346 vdd.n793 185
R17146 vdd.n3348 vdd.n3347 185
R17147 vdd.n3349 vdd.n792 185
R17148 vdd.n3351 vdd.n3350 185
R17149 vdd.n3353 vdd.n790 185
R17150 vdd.n3355 vdd.n3354 185
R17151 vdd.n3356 vdd.n789 185
R17152 vdd.n3358 vdd.n3357 185
R17153 vdd.n3360 vdd.n788 185
R17154 vdd.n3361 vdd.n786 185
R17155 vdd.n3364 vdd.n3363 185
R17156 vdd.n787 vdd.n785 185
R17157 vdd.n3220 vdd.n3219 185
R17158 vdd.n3222 vdd.n3221 185
R17159 vdd.n3224 vdd.n3216 185
R17160 vdd.n3226 vdd.n3225 185
R17161 vdd.n3227 vdd.n3215 185
R17162 vdd.n3229 vdd.n3228 185
R17163 vdd.n3231 vdd.n3213 185
R17164 vdd.n3233 vdd.n3232 185
R17165 vdd.n3234 vdd.n3212 185
R17166 vdd.n3236 vdd.n3235 185
R17167 vdd.n3238 vdd.n3210 185
R17168 vdd.n3240 vdd.n3239 185
R17169 vdd.n3241 vdd.n3209 185
R17170 vdd.n3243 vdd.n3242 185
R17171 vdd.n3245 vdd.n3208 185
R17172 vdd.n3247 vdd.n3246 185
R17173 vdd.n3246 vdd.n692 185
R17174 vdd.n3332 vdd.n802 185
R17175 vdd.n3332 vdd.n3331 185
R17176 vdd.n2949 vdd.n804 185
R17177 vdd.n805 vdd.n804 185
R17178 vdd.n2950 vdd.n838 185
R17179 vdd.n3261 vdd.n838 185
R17180 vdd.n2952 vdd.n2951 185
R17181 vdd.n2951 vdd.n846 185
R17182 vdd.n2953 vdd.n845 185
R17183 vdd.n3255 vdd.n845 185
R17184 vdd.n2955 vdd.n2954 185
R17185 vdd.n2954 vdd.n843 185
R17186 vdd.n2956 vdd.n853 185
R17187 vdd.n3204 vdd.n853 185
R17188 vdd.n2958 vdd.n2957 185
R17189 vdd.n2957 vdd.n851 185
R17190 vdd.n2959 vdd.n858 185
R17191 vdd.n3198 vdd.n858 185
R17192 vdd.n2961 vdd.n2960 185
R17193 vdd.n2960 vdd.n864 185
R17194 vdd.n2962 vdd.n863 185
R17195 vdd.n3192 vdd.n863 185
R17196 vdd.n2964 vdd.n2963 185
R17197 vdd.n2963 vdd.n870 185
R17198 vdd.n2965 vdd.n869 185
R17199 vdd.n3186 vdd.n869 185
R17200 vdd.n2967 vdd.n2966 185
R17201 vdd.n2966 vdd.n877 185
R17202 vdd.n2968 vdd.n876 185
R17203 vdd.n3180 vdd.n876 185
R17204 vdd.n2970 vdd.n2969 185
R17205 vdd.n2969 vdd.n874 185
R17206 vdd.n2971 vdd.n883 185
R17207 vdd.n3174 vdd.n883 185
R17208 vdd.n2973 vdd.n2972 185
R17209 vdd.n2972 vdd.n881 185
R17210 vdd.n2974 vdd.n889 185
R17211 vdd.n3168 vdd.n889 185
R17212 vdd.n2976 vdd.n2975 185
R17213 vdd.n2975 vdd.n887 185
R17214 vdd.n2977 vdd.n894 185
R17215 vdd.n3162 vdd.n894 185
R17216 vdd.n2979 vdd.n2978 185
R17217 vdd.n2978 vdd.n901 185
R17218 vdd.n2980 vdd.n900 185
R17219 vdd.n3156 vdd.n900 185
R17220 vdd.n2982 vdd.n2981 185
R17221 vdd.n2981 vdd.n908 185
R17222 vdd.n2983 vdd.n907 185
R17223 vdd.n3150 vdd.n907 185
R17224 vdd.n2985 vdd.n2984 185
R17225 vdd.n2984 vdd.n905 185
R17226 vdd.n2986 vdd.n914 185
R17227 vdd.n3143 vdd.n914 185
R17228 vdd.n2988 vdd.n2987 185
R17229 vdd.n2987 vdd.n912 185
R17230 vdd.n2989 vdd.n919 185
R17231 vdd.n3137 vdd.n919 185
R17232 vdd.n2991 vdd.n2990 185
R17233 vdd.n2990 vdd.n925 185
R17234 vdd.n2992 vdd.n924 185
R17235 vdd.n3131 vdd.n924 185
R17236 vdd.n2994 vdd.n2993 185
R17237 vdd.n2993 vdd.n931 185
R17238 vdd.n2995 vdd.n930 185
R17239 vdd.n3125 vdd.n930 185
R17240 vdd.n2997 vdd.n2996 185
R17241 vdd.n2998 vdd.n2997 185
R17242 vdd.n2898 vdd.n936 185
R17243 vdd.n3119 vdd.n936 185
R17244 vdd.n3006 vdd.n3005 185
R17245 vdd.n3005 vdd.n3004 185
R17246 vdd.n3007 vdd.n942 185
R17247 vdd.n3113 vdd.n942 185
R17248 vdd.n3009 vdd.n3008 185
R17249 vdd.n3008 vdd.n940 185
R17250 vdd.n3010 vdd.n948 185
R17251 vdd.n3107 vdd.n948 185
R17252 vdd.n3012 vdd.n3011 185
R17253 vdd.n3011 vdd.n946 185
R17254 vdd.n3013 vdd.n953 185
R17255 vdd.n3101 vdd.n953 185
R17256 vdd.n3015 vdd.n3014 185
R17257 vdd.n3016 vdd.n3015 185
R17258 vdd.n2897 vdd.n959 185
R17259 vdd.n3095 vdd.n959 185
R17260 vdd.n2896 vdd.n2895 185
R17261 vdd.n2895 vdd.n957 185
R17262 vdd.n2357 vdd.n2356 185
R17263 vdd.n2358 vdd.n2357 185
R17264 vdd.n1531 vdd.n1529 185
R17265 vdd.n2349 vdd.n1529 185
R17266 vdd.n2352 vdd.n2351 185
R17267 vdd.n2351 vdd.n2350 185
R17268 vdd.n1534 vdd.n1533 185
R17269 vdd.n1535 vdd.n1534 185
R17270 vdd.n2338 vdd.n2337 185
R17271 vdd.n2339 vdd.n2338 185
R17272 vdd.n1543 vdd.n1542 185
R17273 vdd.n2330 vdd.n1542 185
R17274 vdd.n2333 vdd.n2332 185
R17275 vdd.n2332 vdd.n2331 185
R17276 vdd.n1546 vdd.n1545 185
R17277 vdd.n1553 vdd.n1546 185
R17278 vdd.n2321 vdd.n2320 185
R17279 vdd.n2322 vdd.n2321 185
R17280 vdd.n1555 vdd.n1554 185
R17281 vdd.n1554 vdd.n1552 185
R17282 vdd.n2316 vdd.n2315 185
R17283 vdd.n2315 vdd.n2314 185
R17284 vdd.n1558 vdd.n1557 185
R17285 vdd.n1559 vdd.n1558 185
R17286 vdd.n2305 vdd.n2304 185
R17287 vdd.n2306 vdd.n2305 185
R17288 vdd.n1566 vdd.n1565 185
R17289 vdd.n2297 vdd.n1565 185
R17290 vdd.n2300 vdd.n2299 185
R17291 vdd.n2299 vdd.n2298 185
R17292 vdd.n1569 vdd.n1568 185
R17293 vdd.n1575 vdd.n1569 185
R17294 vdd.n2288 vdd.n2287 185
R17295 vdd.n2289 vdd.n2288 185
R17296 vdd.n1577 vdd.n1576 185
R17297 vdd.n2280 vdd.n1576 185
R17298 vdd.n2283 vdd.n2282 185
R17299 vdd.n2282 vdd.n2281 185
R17300 vdd.n1580 vdd.n1579 185
R17301 vdd.n1581 vdd.n1580 185
R17302 vdd.n2271 vdd.n2270 185
R17303 vdd.n2272 vdd.n2271 185
R17304 vdd.n1589 vdd.n1588 185
R17305 vdd.n1588 vdd.n1587 185
R17306 vdd.n1959 vdd.n1958 185
R17307 vdd.n1958 vdd.n1957 185
R17308 vdd.n1592 vdd.n1591 185
R17309 vdd.n1598 vdd.n1592 185
R17310 vdd.n1948 vdd.n1947 185
R17311 vdd.n1949 vdd.n1948 185
R17312 vdd.n1600 vdd.n1599 185
R17313 vdd.n1940 vdd.n1599 185
R17314 vdd.n1943 vdd.n1942 185
R17315 vdd.n1942 vdd.n1941 185
R17316 vdd.n1603 vdd.n1602 185
R17317 vdd.n1610 vdd.n1603 185
R17318 vdd.n1931 vdd.n1930 185
R17319 vdd.n1932 vdd.n1931 185
R17320 vdd.n1612 vdd.n1611 185
R17321 vdd.n1611 vdd.n1609 185
R17322 vdd.n1926 vdd.n1925 185
R17323 vdd.n1925 vdd.n1924 185
R17324 vdd.n1615 vdd.n1614 185
R17325 vdd.n1616 vdd.n1615 185
R17326 vdd.n1915 vdd.n1914 185
R17327 vdd.n1916 vdd.n1915 185
R17328 vdd.n1623 vdd.n1622 185
R17329 vdd.n1907 vdd.n1622 185
R17330 vdd.n1910 vdd.n1909 185
R17331 vdd.n1909 vdd.n1908 185
R17332 vdd.n1626 vdd.n1625 185
R17333 vdd.n1632 vdd.n1626 185
R17334 vdd.n1898 vdd.n1897 185
R17335 vdd.n1899 vdd.n1898 185
R17336 vdd.n1634 vdd.n1633 185
R17337 vdd.n1890 vdd.n1633 185
R17338 vdd.n1893 vdd.n1892 185
R17339 vdd.n1892 vdd.n1891 185
R17340 vdd.n1637 vdd.n1636 185
R17341 vdd.n1638 vdd.n1637 185
R17342 vdd.n1881 vdd.n1880 185
R17343 vdd.n1882 vdd.n1881 185
R17344 vdd.n1645 vdd.n1644 185
R17345 vdd.n1680 vdd.n1644 185
R17346 vdd.n1876 vdd.n1875 185
R17347 vdd.n1648 vdd.n1647 185
R17348 vdd.n1872 vdd.n1871 185
R17349 vdd.n1873 vdd.n1872 185
R17350 vdd.n1682 vdd.n1681 185
R17351 vdd.n1867 vdd.n1684 185
R17352 vdd.n1866 vdd.n1685 185
R17353 vdd.n1865 vdd.n1686 185
R17354 vdd.n1688 vdd.n1687 185
R17355 vdd.n1861 vdd.n1690 185
R17356 vdd.n1860 vdd.n1691 185
R17357 vdd.n1859 vdd.n1692 185
R17358 vdd.n1694 vdd.n1693 185
R17359 vdd.n1855 vdd.n1696 185
R17360 vdd.n1854 vdd.n1697 185
R17361 vdd.n1853 vdd.n1698 185
R17362 vdd.n1700 vdd.n1699 185
R17363 vdd.n1849 vdd.n1702 185
R17364 vdd.n1848 vdd.n1703 185
R17365 vdd.n1847 vdd.n1704 185
R17366 vdd.n1708 vdd.n1705 185
R17367 vdd.n1843 vdd.n1710 185
R17368 vdd.n1842 vdd.n1711 185
R17369 vdd.n1841 vdd.n1712 185
R17370 vdd.n1714 vdd.n1713 185
R17371 vdd.n1837 vdd.n1716 185
R17372 vdd.n1836 vdd.n1717 185
R17373 vdd.n1835 vdd.n1718 185
R17374 vdd.n1720 vdd.n1719 185
R17375 vdd.n1831 vdd.n1722 185
R17376 vdd.n1830 vdd.n1723 185
R17377 vdd.n1829 vdd.n1724 185
R17378 vdd.n1726 vdd.n1725 185
R17379 vdd.n1825 vdd.n1728 185
R17380 vdd.n1824 vdd.n1729 185
R17381 vdd.n1823 vdd.n1730 185
R17382 vdd.n1732 vdd.n1731 185
R17383 vdd.n1819 vdd.n1734 185
R17384 vdd.n1818 vdd.n1735 185
R17385 vdd.n1817 vdd.n1736 185
R17386 vdd.n1738 vdd.n1737 185
R17387 vdd.n1813 vdd.n1740 185
R17388 vdd.n1812 vdd.n1809 185
R17389 vdd.n1808 vdd.n1741 185
R17390 vdd.n1743 vdd.n1742 185
R17391 vdd.n1804 vdd.n1745 185
R17392 vdd.n1803 vdd.n1746 185
R17393 vdd.n1802 vdd.n1747 185
R17394 vdd.n1749 vdd.n1748 185
R17395 vdd.n1798 vdd.n1751 185
R17396 vdd.n1797 vdd.n1752 185
R17397 vdd.n1796 vdd.n1753 185
R17398 vdd.n1755 vdd.n1754 185
R17399 vdd.n1792 vdd.n1757 185
R17400 vdd.n1791 vdd.n1758 185
R17401 vdd.n1790 vdd.n1759 185
R17402 vdd.n1761 vdd.n1760 185
R17403 vdd.n1786 vdd.n1763 185
R17404 vdd.n1785 vdd.n1764 185
R17405 vdd.n1784 vdd.n1765 185
R17406 vdd.n1767 vdd.n1766 185
R17407 vdd.n1780 vdd.n1769 185
R17408 vdd.n1779 vdd.n1770 185
R17409 vdd.n1778 vdd.n1771 185
R17410 vdd.n1775 vdd.n1679 185
R17411 vdd.n1873 vdd.n1679 185
R17412 vdd.n2361 vdd.n2360 185
R17413 vdd.n2365 vdd.n1525 185
R17414 vdd.n1524 vdd.n1518 185
R17415 vdd.n1522 vdd.n1521 185
R17416 vdd.n1520 vdd.n1279 185
R17417 vdd.n2369 vdd.n1276 185
R17418 vdd.n2371 vdd.n2370 185
R17419 vdd.n2373 vdd.n1274 185
R17420 vdd.n2375 vdd.n2374 185
R17421 vdd.n2376 vdd.n1269 185
R17422 vdd.n2378 vdd.n2377 185
R17423 vdd.n2380 vdd.n1267 185
R17424 vdd.n2382 vdd.n2381 185
R17425 vdd.n2383 vdd.n1262 185
R17426 vdd.n2385 vdd.n2384 185
R17427 vdd.n2387 vdd.n1260 185
R17428 vdd.n2389 vdd.n2388 185
R17429 vdd.n2390 vdd.n1256 185
R17430 vdd.n2392 vdd.n2391 185
R17431 vdd.n2394 vdd.n1253 185
R17432 vdd.n2396 vdd.n2395 185
R17433 vdd.n1254 vdd.n1247 185
R17434 vdd.n2400 vdd.n1251 185
R17435 vdd.n2401 vdd.n1243 185
R17436 vdd.n2403 vdd.n2402 185
R17437 vdd.n2405 vdd.n1241 185
R17438 vdd.n2407 vdd.n2406 185
R17439 vdd.n2408 vdd.n1236 185
R17440 vdd.n2410 vdd.n2409 185
R17441 vdd.n2412 vdd.n1234 185
R17442 vdd.n2414 vdd.n2413 185
R17443 vdd.n2415 vdd.n1229 185
R17444 vdd.n2417 vdd.n2416 185
R17445 vdd.n2419 vdd.n1227 185
R17446 vdd.n2421 vdd.n2420 185
R17447 vdd.n2422 vdd.n1222 185
R17448 vdd.n2424 vdd.n2423 185
R17449 vdd.n2426 vdd.n1220 185
R17450 vdd.n2428 vdd.n2427 185
R17451 vdd.n2429 vdd.n1216 185
R17452 vdd.n2431 vdd.n2430 185
R17453 vdd.n2433 vdd.n1213 185
R17454 vdd.n2435 vdd.n2434 185
R17455 vdd.n1214 vdd.n1207 185
R17456 vdd.n2439 vdd.n1211 185
R17457 vdd.n2440 vdd.n1203 185
R17458 vdd.n2442 vdd.n2441 185
R17459 vdd.n2444 vdd.n1201 185
R17460 vdd.n2446 vdd.n2445 185
R17461 vdd.n2447 vdd.n1196 185
R17462 vdd.n2449 vdd.n2448 185
R17463 vdd.n2451 vdd.n1194 185
R17464 vdd.n2453 vdd.n2452 185
R17465 vdd.n2454 vdd.n1189 185
R17466 vdd.n2456 vdd.n2455 185
R17467 vdd.n2458 vdd.n1187 185
R17468 vdd.n2460 vdd.n2459 185
R17469 vdd.n2461 vdd.n1185 185
R17470 vdd.n2463 vdd.n2462 185
R17471 vdd.n2466 vdd.n2465 185
R17472 vdd.n2468 vdd.n2467 185
R17473 vdd.n2470 vdd.n1183 185
R17474 vdd.n2472 vdd.n2471 185
R17475 vdd.n1530 vdd.n1182 185
R17476 vdd.n2359 vdd.n1528 185
R17477 vdd.n2359 vdd.n2358 185
R17478 vdd.n1538 vdd.n1527 185
R17479 vdd.n2349 vdd.n1527 185
R17480 vdd.n2348 vdd.n2347 185
R17481 vdd.n2350 vdd.n2348 185
R17482 vdd.n1537 vdd.n1536 185
R17483 vdd.n1536 vdd.n1535 185
R17484 vdd.n2341 vdd.n2340 185
R17485 vdd.n2340 vdd.n2339 185
R17486 vdd.n1541 vdd.n1540 185
R17487 vdd.n2330 vdd.n1541 185
R17488 vdd.n2329 vdd.n2328 185
R17489 vdd.n2331 vdd.n2329 185
R17490 vdd.n1548 vdd.n1547 185
R17491 vdd.n1553 vdd.n1547 185
R17492 vdd.n2324 vdd.n2323 185
R17493 vdd.n2323 vdd.n2322 185
R17494 vdd.n1551 vdd.n1550 185
R17495 vdd.n1552 vdd.n1551 185
R17496 vdd.n2313 vdd.n2312 185
R17497 vdd.n2314 vdd.n2313 185
R17498 vdd.n1561 vdd.n1560 185
R17499 vdd.n1560 vdd.n1559 185
R17500 vdd.n2308 vdd.n2307 185
R17501 vdd.n2307 vdd.n2306 185
R17502 vdd.n1564 vdd.n1563 185
R17503 vdd.n2297 vdd.n1564 185
R17504 vdd.n2296 vdd.n2295 185
R17505 vdd.n2298 vdd.n2296 185
R17506 vdd.n1571 vdd.n1570 185
R17507 vdd.n1575 vdd.n1570 185
R17508 vdd.n2291 vdd.n2290 185
R17509 vdd.n2290 vdd.n2289 185
R17510 vdd.n1574 vdd.n1573 185
R17511 vdd.n2280 vdd.n1574 185
R17512 vdd.n2279 vdd.n2278 185
R17513 vdd.n2281 vdd.n2279 185
R17514 vdd.n1583 vdd.n1582 185
R17515 vdd.n1582 vdd.n1581 185
R17516 vdd.n2274 vdd.n2273 185
R17517 vdd.n2273 vdd.n2272 185
R17518 vdd.n1586 vdd.n1585 185
R17519 vdd.n1587 vdd.n1586 185
R17520 vdd.n1956 vdd.n1955 185
R17521 vdd.n1957 vdd.n1956 185
R17522 vdd.n1594 vdd.n1593 185
R17523 vdd.n1598 vdd.n1593 185
R17524 vdd.n1951 vdd.n1950 185
R17525 vdd.n1950 vdd.n1949 185
R17526 vdd.n1597 vdd.n1596 185
R17527 vdd.n1940 vdd.n1597 185
R17528 vdd.n1939 vdd.n1938 185
R17529 vdd.n1941 vdd.n1939 185
R17530 vdd.n1605 vdd.n1604 185
R17531 vdd.n1610 vdd.n1604 185
R17532 vdd.n1934 vdd.n1933 185
R17533 vdd.n1933 vdd.n1932 185
R17534 vdd.n1608 vdd.n1607 185
R17535 vdd.n1609 vdd.n1608 185
R17536 vdd.n1923 vdd.n1922 185
R17537 vdd.n1924 vdd.n1923 185
R17538 vdd.n1618 vdd.n1617 185
R17539 vdd.n1617 vdd.n1616 185
R17540 vdd.n1918 vdd.n1917 185
R17541 vdd.n1917 vdd.n1916 185
R17542 vdd.n1621 vdd.n1620 185
R17543 vdd.n1907 vdd.n1621 185
R17544 vdd.n1906 vdd.n1905 185
R17545 vdd.n1908 vdd.n1906 185
R17546 vdd.n1628 vdd.n1627 185
R17547 vdd.n1632 vdd.n1627 185
R17548 vdd.n1901 vdd.n1900 185
R17549 vdd.n1900 vdd.n1899 185
R17550 vdd.n1631 vdd.n1630 185
R17551 vdd.n1890 vdd.n1631 185
R17552 vdd.n1889 vdd.n1888 185
R17553 vdd.n1891 vdd.n1889 185
R17554 vdd.n1640 vdd.n1639 185
R17555 vdd.n1639 vdd.n1638 185
R17556 vdd.n1884 vdd.n1883 185
R17557 vdd.n1883 vdd.n1882 185
R17558 vdd.n1643 vdd.n1642 185
R17559 vdd.n1680 vdd.n1643 185
R17560 vdd.n1000 vdd.n998 185
R17561 vdd.n2712 vdd.n998 185
R17562 vdd.n2634 vdd.n1018 185
R17563 vdd.n1018 vdd.n1005 185
R17564 vdd.n2636 vdd.n2635 185
R17565 vdd.n2637 vdd.n2636 185
R17566 vdd.n2633 vdd.n1017 185
R17567 vdd.n1399 vdd.n1017 185
R17568 vdd.n2632 vdd.n2631 185
R17569 vdd.n2631 vdd.n2630 185
R17570 vdd.n1020 vdd.n1019 185
R17571 vdd.n1021 vdd.n1020 185
R17572 vdd.n2621 vdd.n2620 185
R17573 vdd.n2622 vdd.n2621 185
R17574 vdd.n2619 vdd.n1031 185
R17575 vdd.n1031 vdd.n1028 185
R17576 vdd.n2618 vdd.n2617 185
R17577 vdd.n2617 vdd.n2616 185
R17578 vdd.n1033 vdd.n1032 185
R17579 vdd.n1425 vdd.n1033 185
R17580 vdd.n2609 vdd.n2608 185
R17581 vdd.n2610 vdd.n2609 185
R17582 vdd.n2607 vdd.n1041 185
R17583 vdd.n1046 vdd.n1041 185
R17584 vdd.n2606 vdd.n2605 185
R17585 vdd.n2605 vdd.n2604 185
R17586 vdd.n1043 vdd.n1042 185
R17587 vdd.n1052 vdd.n1043 185
R17588 vdd.n2597 vdd.n2596 185
R17589 vdd.n2598 vdd.n2597 185
R17590 vdd.n2595 vdd.n1053 185
R17591 vdd.n1437 vdd.n1053 185
R17592 vdd.n2594 vdd.n2593 185
R17593 vdd.n2593 vdd.n2592 185
R17594 vdd.n1055 vdd.n1054 185
R17595 vdd.n1056 vdd.n1055 185
R17596 vdd.n2585 vdd.n2584 185
R17597 vdd.n2586 vdd.n2585 185
R17598 vdd.n2583 vdd.n1065 185
R17599 vdd.n1065 vdd.n1062 185
R17600 vdd.n2582 vdd.n2581 185
R17601 vdd.n2581 vdd.n2580 185
R17602 vdd.n1067 vdd.n1066 185
R17603 vdd.n1076 vdd.n1067 185
R17604 vdd.n2572 vdd.n2571 185
R17605 vdd.n2573 vdd.n2572 185
R17606 vdd.n2570 vdd.n1077 185
R17607 vdd.n1083 vdd.n1077 185
R17608 vdd.n2569 vdd.n2568 185
R17609 vdd.n2568 vdd.n2567 185
R17610 vdd.n1079 vdd.n1078 185
R17611 vdd.n1080 vdd.n1079 185
R17612 vdd.n2560 vdd.n2559 185
R17613 vdd.n2561 vdd.n2560 185
R17614 vdd.n2558 vdd.n1090 185
R17615 vdd.n1090 vdd.n1087 185
R17616 vdd.n2557 vdd.n2556 185
R17617 vdd.n2556 vdd.n2555 185
R17618 vdd.n1092 vdd.n1091 185
R17619 vdd.n1093 vdd.n1092 185
R17620 vdd.n2548 vdd.n2547 185
R17621 vdd.n2549 vdd.n2548 185
R17622 vdd.n2546 vdd.n1101 185
R17623 vdd.n1106 vdd.n1101 185
R17624 vdd.n2545 vdd.n2544 185
R17625 vdd.n2544 vdd.n2543 185
R17626 vdd.n1103 vdd.n1102 185
R17627 vdd.n1112 vdd.n1103 185
R17628 vdd.n2536 vdd.n2535 185
R17629 vdd.n2537 vdd.n2536 185
R17630 vdd.n2534 vdd.n1113 185
R17631 vdd.n1119 vdd.n1113 185
R17632 vdd.n2533 vdd.n2532 185
R17633 vdd.n2532 vdd.n2531 185
R17634 vdd.n1115 vdd.n1114 185
R17635 vdd.n1116 vdd.n1115 185
R17636 vdd.n2524 vdd.n2523 185
R17637 vdd.n2525 vdd.n2524 185
R17638 vdd.n2522 vdd.n1126 185
R17639 vdd.n1126 vdd.n1123 185
R17640 vdd.n2521 vdd.n2520 185
R17641 vdd.n2520 vdd.n2519 185
R17642 vdd.n1128 vdd.n1127 185
R17643 vdd.n1137 vdd.n1128 185
R17644 vdd.n2512 vdd.n2511 185
R17645 vdd.n2513 vdd.n2512 185
R17646 vdd.n2510 vdd.n1138 185
R17647 vdd.n1138 vdd.n1134 185
R17648 vdd.n2509 vdd.n2508 185
R17649 vdd.n1140 vdd.n1139 185
R17650 vdd.n2505 vdd.n2504 185
R17651 vdd.n2506 vdd.n2505 185
R17652 vdd.n2503 vdd.n1176 185
R17653 vdd.n2502 vdd.n2501 185
R17654 vdd.n2500 vdd.n2499 185
R17655 vdd.n2498 vdd.n2497 185
R17656 vdd.n2496 vdd.n2495 185
R17657 vdd.n2494 vdd.n2493 185
R17658 vdd.n2492 vdd.n2491 185
R17659 vdd.n2490 vdd.n2489 185
R17660 vdd.n2488 vdd.n2487 185
R17661 vdd.n2486 vdd.n2485 185
R17662 vdd.n2484 vdd.n2483 185
R17663 vdd.n2482 vdd.n2481 185
R17664 vdd.n2480 vdd.n2479 185
R17665 vdd.n2478 vdd.n2477 185
R17666 vdd.n2476 vdd.n2475 185
R17667 vdd.n1321 vdd.n1177 185
R17668 vdd.n1323 vdd.n1322 185
R17669 vdd.n1325 vdd.n1324 185
R17670 vdd.n1327 vdd.n1326 185
R17671 vdd.n1329 vdd.n1328 185
R17672 vdd.n1331 vdd.n1330 185
R17673 vdd.n1333 vdd.n1332 185
R17674 vdd.n1335 vdd.n1334 185
R17675 vdd.n1337 vdd.n1336 185
R17676 vdd.n1339 vdd.n1338 185
R17677 vdd.n1341 vdd.n1340 185
R17678 vdd.n1343 vdd.n1342 185
R17679 vdd.n1345 vdd.n1344 185
R17680 vdd.n1347 vdd.n1346 185
R17681 vdd.n1350 vdd.n1349 185
R17682 vdd.n1352 vdd.n1351 185
R17683 vdd.n1354 vdd.n1353 185
R17684 vdd.n2715 vdd.n2714 185
R17685 vdd.n2717 vdd.n2716 185
R17686 vdd.n2719 vdd.n2718 185
R17687 vdd.n2722 vdd.n2721 185
R17688 vdd.n2724 vdd.n2723 185
R17689 vdd.n2726 vdd.n2725 185
R17690 vdd.n2728 vdd.n2727 185
R17691 vdd.n2730 vdd.n2729 185
R17692 vdd.n2732 vdd.n2731 185
R17693 vdd.n2734 vdd.n2733 185
R17694 vdd.n2736 vdd.n2735 185
R17695 vdd.n2738 vdd.n2737 185
R17696 vdd.n2740 vdd.n2739 185
R17697 vdd.n2742 vdd.n2741 185
R17698 vdd.n2744 vdd.n2743 185
R17699 vdd.n2746 vdd.n2745 185
R17700 vdd.n2748 vdd.n2747 185
R17701 vdd.n2750 vdd.n2749 185
R17702 vdd.n2752 vdd.n2751 185
R17703 vdd.n2754 vdd.n2753 185
R17704 vdd.n2756 vdd.n2755 185
R17705 vdd.n2758 vdd.n2757 185
R17706 vdd.n2760 vdd.n2759 185
R17707 vdd.n2762 vdd.n2761 185
R17708 vdd.n2764 vdd.n2763 185
R17709 vdd.n2766 vdd.n2765 185
R17710 vdd.n2768 vdd.n2767 185
R17711 vdd.n2770 vdd.n2769 185
R17712 vdd.n2772 vdd.n2771 185
R17713 vdd.n2774 vdd.n2773 185
R17714 vdd.n2776 vdd.n2775 185
R17715 vdd.n2778 vdd.n2777 185
R17716 vdd.n2780 vdd.n2779 185
R17717 vdd.n2781 vdd.n999 185
R17718 vdd.n2783 vdd.n2782 185
R17719 vdd.n2784 vdd.n2783 185
R17720 vdd.n2713 vdd.n1003 185
R17721 vdd.n2713 vdd.n2712 185
R17722 vdd.n1397 vdd.n1004 185
R17723 vdd.n1005 vdd.n1004 185
R17724 vdd.n1398 vdd.n1015 185
R17725 vdd.n2637 vdd.n1015 185
R17726 vdd.n1401 vdd.n1400 185
R17727 vdd.n1400 vdd.n1399 185
R17728 vdd.n1402 vdd.n1022 185
R17729 vdd.n2630 vdd.n1022 185
R17730 vdd.n1404 vdd.n1403 185
R17731 vdd.n1403 vdd.n1021 185
R17732 vdd.n1405 vdd.n1029 185
R17733 vdd.n2622 vdd.n1029 185
R17734 vdd.n1407 vdd.n1406 185
R17735 vdd.n1406 vdd.n1028 185
R17736 vdd.n1408 vdd.n1034 185
R17737 vdd.n2616 vdd.n1034 185
R17738 vdd.n1427 vdd.n1426 185
R17739 vdd.n1426 vdd.n1425 185
R17740 vdd.n1428 vdd.n1039 185
R17741 vdd.n2610 vdd.n1039 185
R17742 vdd.n1430 vdd.n1429 185
R17743 vdd.n1429 vdd.n1046 185
R17744 vdd.n1431 vdd.n1044 185
R17745 vdd.n2604 vdd.n1044 185
R17746 vdd.n1433 vdd.n1432 185
R17747 vdd.n1432 vdd.n1052 185
R17748 vdd.n1434 vdd.n1050 185
R17749 vdd.n2598 vdd.n1050 185
R17750 vdd.n1436 vdd.n1435 185
R17751 vdd.n1437 vdd.n1436 185
R17752 vdd.n1396 vdd.n1057 185
R17753 vdd.n2592 vdd.n1057 185
R17754 vdd.n1395 vdd.n1394 185
R17755 vdd.n1394 vdd.n1056 185
R17756 vdd.n1393 vdd.n1063 185
R17757 vdd.n2586 vdd.n1063 185
R17758 vdd.n1392 vdd.n1391 185
R17759 vdd.n1391 vdd.n1062 185
R17760 vdd.n1390 vdd.n1068 185
R17761 vdd.n2580 vdd.n1068 185
R17762 vdd.n1389 vdd.n1388 185
R17763 vdd.n1388 vdd.n1076 185
R17764 vdd.n1387 vdd.n1074 185
R17765 vdd.n2573 vdd.n1074 185
R17766 vdd.n1386 vdd.n1385 185
R17767 vdd.n1385 vdd.n1083 185
R17768 vdd.n1384 vdd.n1081 185
R17769 vdd.n2567 vdd.n1081 185
R17770 vdd.n1383 vdd.n1382 185
R17771 vdd.n1382 vdd.n1080 185
R17772 vdd.n1381 vdd.n1088 185
R17773 vdd.n2561 vdd.n1088 185
R17774 vdd.n1380 vdd.n1379 185
R17775 vdd.n1379 vdd.n1087 185
R17776 vdd.n1378 vdd.n1094 185
R17777 vdd.n2555 vdd.n1094 185
R17778 vdd.n1377 vdd.n1376 185
R17779 vdd.n1376 vdd.n1093 185
R17780 vdd.n1375 vdd.n1099 185
R17781 vdd.n2549 vdd.n1099 185
R17782 vdd.n1374 vdd.n1373 185
R17783 vdd.n1373 vdd.n1106 185
R17784 vdd.n1372 vdd.n1104 185
R17785 vdd.n2543 vdd.n1104 185
R17786 vdd.n1371 vdd.n1370 185
R17787 vdd.n1370 vdd.n1112 185
R17788 vdd.n1369 vdd.n1110 185
R17789 vdd.n2537 vdd.n1110 185
R17790 vdd.n1368 vdd.n1367 185
R17791 vdd.n1367 vdd.n1119 185
R17792 vdd.n1366 vdd.n1117 185
R17793 vdd.n2531 vdd.n1117 185
R17794 vdd.n1365 vdd.n1364 185
R17795 vdd.n1364 vdd.n1116 185
R17796 vdd.n1363 vdd.n1124 185
R17797 vdd.n2525 vdd.n1124 185
R17798 vdd.n1362 vdd.n1361 185
R17799 vdd.n1361 vdd.n1123 185
R17800 vdd.n1360 vdd.n1129 185
R17801 vdd.n2519 vdd.n1129 185
R17802 vdd.n1359 vdd.n1358 185
R17803 vdd.n1358 vdd.n1137 185
R17804 vdd.n1357 vdd.n1135 185
R17805 vdd.n2513 vdd.n1135 185
R17806 vdd.n1356 vdd.n1355 185
R17807 vdd.n1355 vdd.n1134 185
R17808 vdd.n3629 vdd.n3628 185
R17809 vdd.n3628 vdd.n3627 185
R17810 vdd.n3630 vdd.n387 185
R17811 vdd.n387 vdd.n386 185
R17812 vdd.n3632 vdd.n3631 185
R17813 vdd.n3633 vdd.n3632 185
R17814 vdd.n382 vdd.n381 185
R17815 vdd.n3634 vdd.n382 185
R17816 vdd.n3637 vdd.n3636 185
R17817 vdd.n3636 vdd.n3635 185
R17818 vdd.n3638 vdd.n376 185
R17819 vdd.n376 vdd.n375 185
R17820 vdd.n3640 vdd.n3639 185
R17821 vdd.n3641 vdd.n3640 185
R17822 vdd.n371 vdd.n370 185
R17823 vdd.n3642 vdd.n371 185
R17824 vdd.n3645 vdd.n3644 185
R17825 vdd.n3644 vdd.n3643 185
R17826 vdd.n3646 vdd.n365 185
R17827 vdd.n3603 vdd.n365 185
R17828 vdd.n3648 vdd.n3647 185
R17829 vdd.n3649 vdd.n3648 185
R17830 vdd.n360 vdd.n359 185
R17831 vdd.n3650 vdd.n360 185
R17832 vdd.n3653 vdd.n3652 185
R17833 vdd.n3652 vdd.n3651 185
R17834 vdd.n3654 vdd.n354 185
R17835 vdd.n361 vdd.n354 185
R17836 vdd.n3656 vdd.n3655 185
R17837 vdd.n3657 vdd.n3656 185
R17838 vdd.n350 vdd.n349 185
R17839 vdd.n3658 vdd.n350 185
R17840 vdd.n3661 vdd.n3660 185
R17841 vdd.n3660 vdd.n3659 185
R17842 vdd.n3662 vdd.n345 185
R17843 vdd.n345 vdd.n344 185
R17844 vdd.n3664 vdd.n3663 185
R17845 vdd.n3665 vdd.n3664 185
R17846 vdd.n339 vdd.n337 185
R17847 vdd.n3666 vdd.n339 185
R17848 vdd.n3669 vdd.n3668 185
R17849 vdd.n3668 vdd.n3667 185
R17850 vdd.n338 vdd.n336 185
R17851 vdd.n340 vdd.n338 185
R17852 vdd.n3579 vdd.n3578 185
R17853 vdd.n3580 vdd.n3579 185
R17854 vdd.n635 vdd.n634 185
R17855 vdd.n634 vdd.n633 185
R17856 vdd.n3574 vdd.n3573 185
R17857 vdd.n3573 vdd.n3572 185
R17858 vdd.n638 vdd.n637 185
R17859 vdd.n644 vdd.n638 185
R17860 vdd.n3560 vdd.n3559 185
R17861 vdd.n3561 vdd.n3560 185
R17862 vdd.n646 vdd.n645 185
R17863 vdd.n3552 vdd.n645 185
R17864 vdd.n3555 vdd.n3554 185
R17865 vdd.n3554 vdd.n3553 185
R17866 vdd.n649 vdd.n648 185
R17867 vdd.n656 vdd.n649 185
R17868 vdd.n3543 vdd.n3542 185
R17869 vdd.n3544 vdd.n3543 185
R17870 vdd.n658 vdd.n657 185
R17871 vdd.n657 vdd.n655 185
R17872 vdd.n3538 vdd.n3537 185
R17873 vdd.n3537 vdd.n3536 185
R17874 vdd.n661 vdd.n660 185
R17875 vdd.n662 vdd.n661 185
R17876 vdd.n3527 vdd.n3526 185
R17877 vdd.n3528 vdd.n3527 185
R17878 vdd.n669 vdd.n668 185
R17879 vdd.n3519 vdd.n668 185
R17880 vdd.n3522 vdd.n3521 185
R17881 vdd.n3521 vdd.n3520 185
R17882 vdd.n672 vdd.n671 185
R17883 vdd.n679 vdd.n672 185
R17884 vdd.n3510 vdd.n3509 185
R17885 vdd.n3511 vdd.n3510 185
R17886 vdd.n681 vdd.n680 185
R17887 vdd.n680 vdd.n678 185
R17888 vdd.n3505 vdd.n3504 185
R17889 vdd.n3504 vdd.n3503 185
R17890 vdd.n684 vdd.n683 185
R17891 vdd.n723 vdd.n684 185
R17892 vdd.n3493 vdd.n3492 185
R17893 vdd.n3491 vdd.n725 185
R17894 vdd.n3490 vdd.n724 185
R17895 vdd.n3495 vdd.n724 185
R17896 vdd.n729 vdd.n728 185
R17897 vdd.n733 vdd.n732 185
R17898 vdd.n3486 vdd.n734 185
R17899 vdd.n3485 vdd.n3484 185
R17900 vdd.n3483 vdd.n3482 185
R17901 vdd.n3481 vdd.n3480 185
R17902 vdd.n3479 vdd.n3478 185
R17903 vdd.n3477 vdd.n3476 185
R17904 vdd.n3475 vdd.n3474 185
R17905 vdd.n3473 vdd.n3472 185
R17906 vdd.n3471 vdd.n3470 185
R17907 vdd.n3469 vdd.n3468 185
R17908 vdd.n3467 vdd.n3466 185
R17909 vdd.n3465 vdd.n3464 185
R17910 vdd.n3463 vdd.n3462 185
R17911 vdd.n3461 vdd.n3460 185
R17912 vdd.n3459 vdd.n3458 185
R17913 vdd.n3450 vdd.n747 185
R17914 vdd.n3452 vdd.n3451 185
R17915 vdd.n3449 vdd.n3448 185
R17916 vdd.n3447 vdd.n3446 185
R17917 vdd.n3445 vdd.n3444 185
R17918 vdd.n3443 vdd.n3442 185
R17919 vdd.n3441 vdd.n3440 185
R17920 vdd.n3439 vdd.n3438 185
R17921 vdd.n3437 vdd.n3436 185
R17922 vdd.n3435 vdd.n3434 185
R17923 vdd.n3433 vdd.n3432 185
R17924 vdd.n3431 vdd.n3430 185
R17925 vdd.n3429 vdd.n3428 185
R17926 vdd.n3427 vdd.n3426 185
R17927 vdd.n3425 vdd.n3424 185
R17928 vdd.n3423 vdd.n3422 185
R17929 vdd.n3421 vdd.n3420 185
R17930 vdd.n3419 vdd.n3418 185
R17931 vdd.n3417 vdd.n3416 185
R17932 vdd.n3415 vdd.n3414 185
R17933 vdd.n3413 vdd.n3412 185
R17934 vdd.n3411 vdd.n3410 185
R17935 vdd.n3404 vdd.n767 185
R17936 vdd.n3406 vdd.n3405 185
R17937 vdd.n3403 vdd.n3402 185
R17938 vdd.n3401 vdd.n3400 185
R17939 vdd.n3399 vdd.n3398 185
R17940 vdd.n3397 vdd.n3396 185
R17941 vdd.n3395 vdd.n3394 185
R17942 vdd.n3393 vdd.n3392 185
R17943 vdd.n3391 vdd.n3390 185
R17944 vdd.n3389 vdd.n3388 185
R17945 vdd.n3387 vdd.n3386 185
R17946 vdd.n3385 vdd.n3384 185
R17947 vdd.n3383 vdd.n3382 185
R17948 vdd.n3381 vdd.n3380 185
R17949 vdd.n3379 vdd.n3378 185
R17950 vdd.n3377 vdd.n3376 185
R17951 vdd.n3375 vdd.n3374 185
R17952 vdd.n3373 vdd.n3372 185
R17953 vdd.n3371 vdd.n3370 185
R17954 vdd.n3369 vdd.n3368 185
R17955 vdd.n3367 vdd.n691 185
R17956 vdd.n3497 vdd.n3496 185
R17957 vdd.n3496 vdd.n3495 185
R17958 vdd.n3624 vdd.n3623 185
R17959 vdd.n618 vdd.n425 185
R17960 vdd.n617 vdd.n616 185
R17961 vdd.n615 vdd.n614 185
R17962 vdd.n613 vdd.n430 185
R17963 vdd.n609 vdd.n608 185
R17964 vdd.n607 vdd.n606 185
R17965 vdd.n605 vdd.n604 185
R17966 vdd.n603 vdd.n432 185
R17967 vdd.n599 vdd.n598 185
R17968 vdd.n597 vdd.n596 185
R17969 vdd.n595 vdd.n594 185
R17970 vdd.n593 vdd.n434 185
R17971 vdd.n589 vdd.n588 185
R17972 vdd.n587 vdd.n586 185
R17973 vdd.n585 vdd.n584 185
R17974 vdd.n583 vdd.n436 185
R17975 vdd.n579 vdd.n578 185
R17976 vdd.n577 vdd.n576 185
R17977 vdd.n575 vdd.n574 185
R17978 vdd.n573 vdd.n438 185
R17979 vdd.n569 vdd.n568 185
R17980 vdd.n567 vdd.n566 185
R17981 vdd.n565 vdd.n564 185
R17982 vdd.n563 vdd.n442 185
R17983 vdd.n559 vdd.n558 185
R17984 vdd.n557 vdd.n556 185
R17985 vdd.n555 vdd.n554 185
R17986 vdd.n553 vdd.n444 185
R17987 vdd.n549 vdd.n548 185
R17988 vdd.n547 vdd.n546 185
R17989 vdd.n545 vdd.n544 185
R17990 vdd.n543 vdd.n446 185
R17991 vdd.n539 vdd.n538 185
R17992 vdd.n537 vdd.n536 185
R17993 vdd.n535 vdd.n534 185
R17994 vdd.n533 vdd.n448 185
R17995 vdd.n529 vdd.n528 185
R17996 vdd.n527 vdd.n526 185
R17997 vdd.n525 vdd.n524 185
R17998 vdd.n523 vdd.n450 185
R17999 vdd.n519 vdd.n518 185
R18000 vdd.n517 vdd.n516 185
R18001 vdd.n515 vdd.n514 185
R18002 vdd.n513 vdd.n454 185
R18003 vdd.n509 vdd.n508 185
R18004 vdd.n507 vdd.n506 185
R18005 vdd.n505 vdd.n504 185
R18006 vdd.n503 vdd.n456 185
R18007 vdd.n499 vdd.n498 185
R18008 vdd.n497 vdd.n496 185
R18009 vdd.n495 vdd.n494 185
R18010 vdd.n493 vdd.n458 185
R18011 vdd.n489 vdd.n488 185
R18012 vdd.n487 vdd.n486 185
R18013 vdd.n485 vdd.n484 185
R18014 vdd.n483 vdd.n460 185
R18015 vdd.n479 vdd.n478 185
R18016 vdd.n477 vdd.n476 185
R18017 vdd.n475 vdd.n474 185
R18018 vdd.n473 vdd.n462 185
R18019 vdd.n469 vdd.n468 185
R18020 vdd.n467 vdd.n466 185
R18021 vdd.n465 vdd.n392 185
R18022 vdd.n3620 vdd.n393 185
R18023 vdd.n3627 vdd.n393 185
R18024 vdd.n3619 vdd.n3618 185
R18025 vdd.n3618 vdd.n386 185
R18026 vdd.n3617 vdd.n385 185
R18027 vdd.n3633 vdd.n385 185
R18028 vdd.n621 vdd.n384 185
R18029 vdd.n3634 vdd.n384 185
R18030 vdd.n3613 vdd.n383 185
R18031 vdd.n3635 vdd.n383 185
R18032 vdd.n3612 vdd.n3611 185
R18033 vdd.n3611 vdd.n375 185
R18034 vdd.n3610 vdd.n374 185
R18035 vdd.n3641 vdd.n374 185
R18036 vdd.n623 vdd.n373 185
R18037 vdd.n3642 vdd.n373 185
R18038 vdd.n3606 vdd.n372 185
R18039 vdd.n3643 vdd.n372 185
R18040 vdd.n3605 vdd.n3604 185
R18041 vdd.n3604 vdd.n3603 185
R18042 vdd.n3602 vdd.n364 185
R18043 vdd.n3649 vdd.n364 185
R18044 vdd.n625 vdd.n363 185
R18045 vdd.n3650 vdd.n363 185
R18046 vdd.n3598 vdd.n362 185
R18047 vdd.n3651 vdd.n362 185
R18048 vdd.n3597 vdd.n3596 185
R18049 vdd.n3596 vdd.n361 185
R18050 vdd.n3595 vdd.n353 185
R18051 vdd.n3657 vdd.n353 185
R18052 vdd.n627 vdd.n352 185
R18053 vdd.n3658 vdd.n352 185
R18054 vdd.n3591 vdd.n351 185
R18055 vdd.n3659 vdd.n351 185
R18056 vdd.n3590 vdd.n3589 185
R18057 vdd.n3589 vdd.n344 185
R18058 vdd.n3588 vdd.n343 185
R18059 vdd.n3665 vdd.n343 185
R18060 vdd.n629 vdd.n342 185
R18061 vdd.n3666 vdd.n342 185
R18062 vdd.n3584 vdd.n341 185
R18063 vdd.n3667 vdd.n341 185
R18064 vdd.n3583 vdd.n3582 185
R18065 vdd.n3582 vdd.n340 185
R18066 vdd.n3581 vdd.n631 185
R18067 vdd.n3581 vdd.n3580 185
R18068 vdd.n3569 vdd.n632 185
R18069 vdd.n633 vdd.n632 185
R18070 vdd.n3571 vdd.n3570 185
R18071 vdd.n3572 vdd.n3571 185
R18072 vdd.n640 vdd.n639 185
R18073 vdd.n644 vdd.n639 185
R18074 vdd.n3563 vdd.n3562 185
R18075 vdd.n3562 vdd.n3561 185
R18076 vdd.n643 vdd.n642 185
R18077 vdd.n3552 vdd.n643 185
R18078 vdd.n3551 vdd.n3550 185
R18079 vdd.n3553 vdd.n3551 185
R18080 vdd.n651 vdd.n650 185
R18081 vdd.n656 vdd.n650 185
R18082 vdd.n3546 vdd.n3545 185
R18083 vdd.n3545 vdd.n3544 185
R18084 vdd.n654 vdd.n653 185
R18085 vdd.n655 vdd.n654 185
R18086 vdd.n3535 vdd.n3534 185
R18087 vdd.n3536 vdd.n3535 185
R18088 vdd.n664 vdd.n663 185
R18089 vdd.n663 vdd.n662 185
R18090 vdd.n3530 vdd.n3529 185
R18091 vdd.n3529 vdd.n3528 185
R18092 vdd.n667 vdd.n666 185
R18093 vdd.n3519 vdd.n667 185
R18094 vdd.n3518 vdd.n3517 185
R18095 vdd.n3520 vdd.n3518 185
R18096 vdd.n674 vdd.n673 185
R18097 vdd.n679 vdd.n673 185
R18098 vdd.n3513 vdd.n3512 185
R18099 vdd.n3512 vdd.n3511 185
R18100 vdd.n677 vdd.n676 185
R18101 vdd.n678 vdd.n677 185
R18102 vdd.n3502 vdd.n3501 185
R18103 vdd.n3503 vdd.n3502 185
R18104 vdd.n686 vdd.n685 185
R18105 vdd.n723 vdd.n685 185
R18106 vdd.n3091 vdd.n3090 185
R18107 vdd.n962 vdd.n961 185
R18108 vdd.n3087 vdd.n3086 185
R18109 vdd.n3088 vdd.n3087 185
R18110 vdd.n3085 vdd.n2819 185
R18111 vdd.n3084 vdd.n3083 185
R18112 vdd.n3082 vdd.n3081 185
R18113 vdd.n3080 vdd.n3079 185
R18114 vdd.n3078 vdd.n3077 185
R18115 vdd.n3076 vdd.n3075 185
R18116 vdd.n3074 vdd.n3073 185
R18117 vdd.n3072 vdd.n3071 185
R18118 vdd.n3070 vdd.n3069 185
R18119 vdd.n3068 vdd.n3067 185
R18120 vdd.n3066 vdd.n3065 185
R18121 vdd.n3064 vdd.n3063 185
R18122 vdd.n3062 vdd.n3061 185
R18123 vdd.n3060 vdd.n3059 185
R18124 vdd.n3058 vdd.n3057 185
R18125 vdd.n3056 vdd.n3055 185
R18126 vdd.n3054 vdd.n3053 185
R18127 vdd.n3052 vdd.n3051 185
R18128 vdd.n3050 vdd.n3049 185
R18129 vdd.n3048 vdd.n3047 185
R18130 vdd.n3046 vdd.n3045 185
R18131 vdd.n3044 vdd.n3043 185
R18132 vdd.n3042 vdd.n3041 185
R18133 vdd.n3040 vdd.n3039 185
R18134 vdd.n3038 vdd.n3037 185
R18135 vdd.n3036 vdd.n3035 185
R18136 vdd.n3034 vdd.n3033 185
R18137 vdd.n3032 vdd.n3031 185
R18138 vdd.n3030 vdd.n3029 185
R18139 vdd.n3027 vdd.n3026 185
R18140 vdd.n3025 vdd.n3024 185
R18141 vdd.n3023 vdd.n3022 185
R18142 vdd.n3267 vdd.n3266 185
R18143 vdd.n3269 vdd.n834 185
R18144 vdd.n3271 vdd.n3270 185
R18145 vdd.n3273 vdd.n831 185
R18146 vdd.n3275 vdd.n3274 185
R18147 vdd.n3277 vdd.n829 185
R18148 vdd.n3279 vdd.n3278 185
R18149 vdd.n3280 vdd.n828 185
R18150 vdd.n3282 vdd.n3281 185
R18151 vdd.n3284 vdd.n826 185
R18152 vdd.n3286 vdd.n3285 185
R18153 vdd.n3287 vdd.n825 185
R18154 vdd.n3289 vdd.n3288 185
R18155 vdd.n3291 vdd.n823 185
R18156 vdd.n3293 vdd.n3292 185
R18157 vdd.n3294 vdd.n822 185
R18158 vdd.n3296 vdd.n3295 185
R18159 vdd.n3298 vdd.n731 185
R18160 vdd.n3300 vdd.n3299 185
R18161 vdd.n3302 vdd.n820 185
R18162 vdd.n3304 vdd.n3303 185
R18163 vdd.n3305 vdd.n819 185
R18164 vdd.n3307 vdd.n3306 185
R18165 vdd.n3309 vdd.n817 185
R18166 vdd.n3311 vdd.n3310 185
R18167 vdd.n3312 vdd.n816 185
R18168 vdd.n3314 vdd.n3313 185
R18169 vdd.n3316 vdd.n814 185
R18170 vdd.n3318 vdd.n3317 185
R18171 vdd.n3319 vdd.n813 185
R18172 vdd.n3321 vdd.n3320 185
R18173 vdd.n3323 vdd.n812 185
R18174 vdd.n3324 vdd.n811 185
R18175 vdd.n3327 vdd.n3326 185
R18176 vdd.n3328 vdd.n809 185
R18177 vdd.n809 vdd.n692 185
R18178 vdd.n3265 vdd.n806 185
R18179 vdd.n3331 vdd.n806 185
R18180 vdd.n3264 vdd.n3263 185
R18181 vdd.n3263 vdd.n805 185
R18182 vdd.n3262 vdd.n836 185
R18183 vdd.n3262 vdd.n3261 185
R18184 vdd.n2905 vdd.n837 185
R18185 vdd.n846 vdd.n837 185
R18186 vdd.n2906 vdd.n844 185
R18187 vdd.n3255 vdd.n844 185
R18188 vdd.n2908 vdd.n2907 185
R18189 vdd.n2907 vdd.n843 185
R18190 vdd.n2909 vdd.n852 185
R18191 vdd.n3204 vdd.n852 185
R18192 vdd.n2911 vdd.n2910 185
R18193 vdd.n2910 vdd.n851 185
R18194 vdd.n2912 vdd.n857 185
R18195 vdd.n3198 vdd.n857 185
R18196 vdd.n2914 vdd.n2913 185
R18197 vdd.n2913 vdd.n864 185
R18198 vdd.n2915 vdd.n862 185
R18199 vdd.n3192 vdd.n862 185
R18200 vdd.n2917 vdd.n2916 185
R18201 vdd.n2916 vdd.n870 185
R18202 vdd.n2918 vdd.n868 185
R18203 vdd.n3186 vdd.n868 185
R18204 vdd.n2920 vdd.n2919 185
R18205 vdd.n2919 vdd.n877 185
R18206 vdd.n2921 vdd.n875 185
R18207 vdd.n3180 vdd.n875 185
R18208 vdd.n2923 vdd.n2922 185
R18209 vdd.n2922 vdd.n874 185
R18210 vdd.n2924 vdd.n882 185
R18211 vdd.n3174 vdd.n882 185
R18212 vdd.n2926 vdd.n2925 185
R18213 vdd.n2925 vdd.n881 185
R18214 vdd.n2927 vdd.n888 185
R18215 vdd.n3168 vdd.n888 185
R18216 vdd.n2929 vdd.n2928 185
R18217 vdd.n2928 vdd.n887 185
R18218 vdd.n2930 vdd.n893 185
R18219 vdd.n3162 vdd.n893 185
R18220 vdd.n2932 vdd.n2931 185
R18221 vdd.n2931 vdd.n901 185
R18222 vdd.n2933 vdd.n899 185
R18223 vdd.n3156 vdd.n899 185
R18224 vdd.n2935 vdd.n2934 185
R18225 vdd.n2934 vdd.n908 185
R18226 vdd.n2936 vdd.n906 185
R18227 vdd.n3150 vdd.n906 185
R18228 vdd.n2938 vdd.n2937 185
R18229 vdd.n2937 vdd.n905 185
R18230 vdd.n2939 vdd.n913 185
R18231 vdd.n3143 vdd.n913 185
R18232 vdd.n2941 vdd.n2940 185
R18233 vdd.n2940 vdd.n912 185
R18234 vdd.n2942 vdd.n918 185
R18235 vdd.n3137 vdd.n918 185
R18236 vdd.n2944 vdd.n2943 185
R18237 vdd.n2943 vdd.n925 185
R18238 vdd.n2945 vdd.n923 185
R18239 vdd.n3131 vdd.n923 185
R18240 vdd.n2947 vdd.n2946 185
R18241 vdd.n2946 vdd.n931 185
R18242 vdd.n2948 vdd.n929 185
R18243 vdd.n3125 vdd.n929 185
R18244 vdd.n3000 vdd.n2999 185
R18245 vdd.n2999 vdd.n2998 185
R18246 vdd.n3001 vdd.n935 185
R18247 vdd.n3119 vdd.n935 185
R18248 vdd.n3003 vdd.n3002 185
R18249 vdd.n3004 vdd.n3003 185
R18250 vdd.n2904 vdd.n941 185
R18251 vdd.n3113 vdd.n941 185
R18252 vdd.n2903 vdd.n2902 185
R18253 vdd.n2902 vdd.n940 185
R18254 vdd.n2901 vdd.n947 185
R18255 vdd.n3107 vdd.n947 185
R18256 vdd.n2900 vdd.n2899 185
R18257 vdd.n2899 vdd.n946 185
R18258 vdd.n2822 vdd.n952 185
R18259 vdd.n3101 vdd.n952 185
R18260 vdd.n3018 vdd.n3017 185
R18261 vdd.n3017 vdd.n3016 185
R18262 vdd.n3019 vdd.n958 185
R18263 vdd.n3095 vdd.n958 185
R18264 vdd.n3021 vdd.n3020 185
R18265 vdd.n3021 vdd.n957 185
R18266 vdd.n3092 vdd.n960 185
R18267 vdd.n960 vdd.n957 185
R18268 vdd.n3094 vdd.n3093 185
R18269 vdd.n3095 vdd.n3094 185
R18270 vdd.n951 vdd.n950 185
R18271 vdd.n3016 vdd.n951 185
R18272 vdd.n3103 vdd.n3102 185
R18273 vdd.n3102 vdd.n3101 185
R18274 vdd.n3104 vdd.n949 185
R18275 vdd.n949 vdd.n946 185
R18276 vdd.n3106 vdd.n3105 185
R18277 vdd.n3107 vdd.n3106 185
R18278 vdd.n939 vdd.n938 185
R18279 vdd.n940 vdd.n939 185
R18280 vdd.n3115 vdd.n3114 185
R18281 vdd.n3114 vdd.n3113 185
R18282 vdd.n3116 vdd.n937 185
R18283 vdd.n3004 vdd.n937 185
R18284 vdd.n3118 vdd.n3117 185
R18285 vdd.n3119 vdd.n3118 185
R18286 vdd.n928 vdd.n927 185
R18287 vdd.n2998 vdd.n928 185
R18288 vdd.n3127 vdd.n3126 185
R18289 vdd.n3126 vdd.n3125 185
R18290 vdd.n3128 vdd.n926 185
R18291 vdd.n931 vdd.n926 185
R18292 vdd.n3130 vdd.n3129 185
R18293 vdd.n3131 vdd.n3130 185
R18294 vdd.n917 vdd.n916 185
R18295 vdd.n925 vdd.n917 185
R18296 vdd.n3139 vdd.n3138 185
R18297 vdd.n3138 vdd.n3137 185
R18298 vdd.n3140 vdd.n915 185
R18299 vdd.n915 vdd.n912 185
R18300 vdd.n3142 vdd.n3141 185
R18301 vdd.n3143 vdd.n3142 185
R18302 vdd.n904 vdd.n903 185
R18303 vdd.n905 vdd.n904 185
R18304 vdd.n3152 vdd.n3151 185
R18305 vdd.n3151 vdd.n3150 185
R18306 vdd.n3153 vdd.n902 185
R18307 vdd.n908 vdd.n902 185
R18308 vdd.n3155 vdd.n3154 185
R18309 vdd.n3156 vdd.n3155 185
R18310 vdd.n892 vdd.n891 185
R18311 vdd.n901 vdd.n892 185
R18312 vdd.n3164 vdd.n3163 185
R18313 vdd.n3163 vdd.n3162 185
R18314 vdd.n3165 vdd.n890 185
R18315 vdd.n890 vdd.n887 185
R18316 vdd.n3167 vdd.n3166 185
R18317 vdd.n3168 vdd.n3167 185
R18318 vdd.n880 vdd.n879 185
R18319 vdd.n881 vdd.n880 185
R18320 vdd.n3176 vdd.n3175 185
R18321 vdd.n3175 vdd.n3174 185
R18322 vdd.n3177 vdd.n878 185
R18323 vdd.n878 vdd.n874 185
R18324 vdd.n3179 vdd.n3178 185
R18325 vdd.n3180 vdd.n3179 185
R18326 vdd.n867 vdd.n866 185
R18327 vdd.n877 vdd.n867 185
R18328 vdd.n3188 vdd.n3187 185
R18329 vdd.n3187 vdd.n3186 185
R18330 vdd.n3189 vdd.n865 185
R18331 vdd.n870 vdd.n865 185
R18332 vdd.n3191 vdd.n3190 185
R18333 vdd.n3192 vdd.n3191 185
R18334 vdd.n856 vdd.n855 185
R18335 vdd.n864 vdd.n856 185
R18336 vdd.n3200 vdd.n3199 185
R18337 vdd.n3199 vdd.n3198 185
R18338 vdd.n3201 vdd.n854 185
R18339 vdd.n854 vdd.n851 185
R18340 vdd.n3203 vdd.n3202 185
R18341 vdd.n3204 vdd.n3203 185
R18342 vdd.n842 vdd.n841 185
R18343 vdd.n843 vdd.n842 185
R18344 vdd.n3257 vdd.n3256 185
R18345 vdd.n3256 vdd.n3255 185
R18346 vdd.n3258 vdd.n840 185
R18347 vdd.n846 vdd.n840 185
R18348 vdd.n3260 vdd.n3259 185
R18349 vdd.n3261 vdd.n3260 185
R18350 vdd.n810 vdd.n808 185
R18351 vdd.n808 vdd.n805 185
R18352 vdd.n3330 vdd.n3329 185
R18353 vdd.n3331 vdd.n3330 185
R18354 vdd.n2711 vdd.n2710 185
R18355 vdd.n2712 vdd.n2711 185
R18356 vdd.n1009 vdd.n1007 185
R18357 vdd.n1007 vdd.n1005 185
R18358 vdd.n2626 vdd.n1016 185
R18359 vdd.n2637 vdd.n1016 185
R18360 vdd.n2627 vdd.n1025 185
R18361 vdd.n1399 vdd.n1025 185
R18362 vdd.n2629 vdd.n2628 185
R18363 vdd.n2630 vdd.n2629 185
R18364 vdd.n2625 vdd.n1024 185
R18365 vdd.n1024 vdd.n1021 185
R18366 vdd.n2624 vdd.n2623 185
R18367 vdd.n2623 vdd.n2622 185
R18368 vdd.n1027 vdd.n1026 185
R18369 vdd.n1028 vdd.n1027 185
R18370 vdd.n2615 vdd.n2614 185
R18371 vdd.n2616 vdd.n2615 185
R18372 vdd.n2613 vdd.n1036 185
R18373 vdd.n1425 vdd.n1036 185
R18374 vdd.n2612 vdd.n2611 185
R18375 vdd.n2611 vdd.n2610 185
R18376 vdd.n1038 vdd.n1037 185
R18377 vdd.n1046 vdd.n1038 185
R18378 vdd.n2603 vdd.n2602 185
R18379 vdd.n2604 vdd.n2603 185
R18380 vdd.n2601 vdd.n1047 185
R18381 vdd.n1052 vdd.n1047 185
R18382 vdd.n2600 vdd.n2599 185
R18383 vdd.n2599 vdd.n2598 185
R18384 vdd.n1049 vdd.n1048 185
R18385 vdd.n1437 vdd.n1049 185
R18386 vdd.n2591 vdd.n2590 185
R18387 vdd.n2592 vdd.n2591 185
R18388 vdd.n2589 vdd.n1059 185
R18389 vdd.n1059 vdd.n1056 185
R18390 vdd.n2588 vdd.n2587 185
R18391 vdd.n2587 vdd.n2586 185
R18392 vdd.n1061 vdd.n1060 185
R18393 vdd.n1062 vdd.n1061 185
R18394 vdd.n2579 vdd.n2578 185
R18395 vdd.n2580 vdd.n2579 185
R18396 vdd.n2576 vdd.n1070 185
R18397 vdd.n1076 vdd.n1070 185
R18398 vdd.n2575 vdd.n2574 185
R18399 vdd.n2574 vdd.n2573 185
R18400 vdd.n1073 vdd.n1072 185
R18401 vdd.n1083 vdd.n1073 185
R18402 vdd.n2566 vdd.n2565 185
R18403 vdd.n2567 vdd.n2566 185
R18404 vdd.n2564 vdd.n1084 185
R18405 vdd.n1084 vdd.n1080 185
R18406 vdd.n2563 vdd.n2562 185
R18407 vdd.n2562 vdd.n2561 185
R18408 vdd.n1086 vdd.n1085 185
R18409 vdd.n1087 vdd.n1086 185
R18410 vdd.n2554 vdd.n2553 185
R18411 vdd.n2555 vdd.n2554 185
R18412 vdd.n2552 vdd.n1096 185
R18413 vdd.n1096 vdd.n1093 185
R18414 vdd.n2551 vdd.n2550 185
R18415 vdd.n2550 vdd.n2549 185
R18416 vdd.n1098 vdd.n1097 185
R18417 vdd.n1106 vdd.n1098 185
R18418 vdd.n2542 vdd.n2541 185
R18419 vdd.n2543 vdd.n2542 185
R18420 vdd.n2540 vdd.n1107 185
R18421 vdd.n1112 vdd.n1107 185
R18422 vdd.n2539 vdd.n2538 185
R18423 vdd.n2538 vdd.n2537 185
R18424 vdd.n1109 vdd.n1108 185
R18425 vdd.n1119 vdd.n1109 185
R18426 vdd.n2530 vdd.n2529 185
R18427 vdd.n2531 vdd.n2530 185
R18428 vdd.n2528 vdd.n1120 185
R18429 vdd.n1120 vdd.n1116 185
R18430 vdd.n2527 vdd.n2526 185
R18431 vdd.n2526 vdd.n2525 185
R18432 vdd.n1122 vdd.n1121 185
R18433 vdd.n1123 vdd.n1122 185
R18434 vdd.n2518 vdd.n2517 185
R18435 vdd.n2519 vdd.n2518 185
R18436 vdd.n2516 vdd.n1131 185
R18437 vdd.n1137 vdd.n1131 185
R18438 vdd.n2515 vdd.n2514 185
R18439 vdd.n2514 vdd.n2513 185
R18440 vdd.n1133 vdd.n1132 185
R18441 vdd.n1134 vdd.n1133 185
R18442 vdd.n2642 vdd.n980 185
R18443 vdd.n2784 vdd.n980 185
R18444 vdd.n2644 vdd.n2643 185
R18445 vdd.n2646 vdd.n2645 185
R18446 vdd.n2648 vdd.n2647 185
R18447 vdd.n2650 vdd.n2649 185
R18448 vdd.n2652 vdd.n2651 185
R18449 vdd.n2654 vdd.n2653 185
R18450 vdd.n2656 vdd.n2655 185
R18451 vdd.n2658 vdd.n2657 185
R18452 vdd.n2660 vdd.n2659 185
R18453 vdd.n2662 vdd.n2661 185
R18454 vdd.n2664 vdd.n2663 185
R18455 vdd.n2666 vdd.n2665 185
R18456 vdd.n2668 vdd.n2667 185
R18457 vdd.n2670 vdd.n2669 185
R18458 vdd.n2672 vdd.n2671 185
R18459 vdd.n2674 vdd.n2673 185
R18460 vdd.n2676 vdd.n2675 185
R18461 vdd.n2678 vdd.n2677 185
R18462 vdd.n2680 vdd.n2679 185
R18463 vdd.n2682 vdd.n2681 185
R18464 vdd.n2684 vdd.n2683 185
R18465 vdd.n2686 vdd.n2685 185
R18466 vdd.n2688 vdd.n2687 185
R18467 vdd.n2690 vdd.n2689 185
R18468 vdd.n2692 vdd.n2691 185
R18469 vdd.n2694 vdd.n2693 185
R18470 vdd.n2696 vdd.n2695 185
R18471 vdd.n2698 vdd.n2697 185
R18472 vdd.n2700 vdd.n2699 185
R18473 vdd.n2702 vdd.n2701 185
R18474 vdd.n2704 vdd.n2703 185
R18475 vdd.n2706 vdd.n2705 185
R18476 vdd.n2708 vdd.n2707 185
R18477 vdd.n2709 vdd.n1008 185
R18478 vdd.n2641 vdd.n1006 185
R18479 vdd.n2712 vdd.n1006 185
R18480 vdd.n2640 vdd.n2639 185
R18481 vdd.n2639 vdd.n1005 185
R18482 vdd.n2638 vdd.n1013 185
R18483 vdd.n2638 vdd.n2637 185
R18484 vdd.n1415 vdd.n1014 185
R18485 vdd.n1399 vdd.n1014 185
R18486 vdd.n1416 vdd.n1023 185
R18487 vdd.n2630 vdd.n1023 185
R18488 vdd.n1418 vdd.n1417 185
R18489 vdd.n1417 vdd.n1021 185
R18490 vdd.n1419 vdd.n1030 185
R18491 vdd.n2622 vdd.n1030 185
R18492 vdd.n1421 vdd.n1420 185
R18493 vdd.n1420 vdd.n1028 185
R18494 vdd.n1422 vdd.n1035 185
R18495 vdd.n2616 vdd.n1035 185
R18496 vdd.n1424 vdd.n1423 185
R18497 vdd.n1425 vdd.n1424 185
R18498 vdd.n1414 vdd.n1040 185
R18499 vdd.n2610 vdd.n1040 185
R18500 vdd.n1413 vdd.n1412 185
R18501 vdd.n1412 vdd.n1046 185
R18502 vdd.n1411 vdd.n1045 185
R18503 vdd.n2604 vdd.n1045 185
R18504 vdd.n1410 vdd.n1409 185
R18505 vdd.n1409 vdd.n1052 185
R18506 vdd.n1318 vdd.n1051 185
R18507 vdd.n2598 vdd.n1051 185
R18508 vdd.n1439 vdd.n1438 185
R18509 vdd.n1438 vdd.n1437 185
R18510 vdd.n1440 vdd.n1058 185
R18511 vdd.n2592 vdd.n1058 185
R18512 vdd.n1442 vdd.n1441 185
R18513 vdd.n1441 vdd.n1056 185
R18514 vdd.n1443 vdd.n1064 185
R18515 vdd.n2586 vdd.n1064 185
R18516 vdd.n1445 vdd.n1444 185
R18517 vdd.n1444 vdd.n1062 185
R18518 vdd.n1446 vdd.n1069 185
R18519 vdd.n2580 vdd.n1069 185
R18520 vdd.n1448 vdd.n1447 185
R18521 vdd.n1447 vdd.n1076 185
R18522 vdd.n1449 vdd.n1075 185
R18523 vdd.n2573 vdd.n1075 185
R18524 vdd.n1451 vdd.n1450 185
R18525 vdd.n1450 vdd.n1083 185
R18526 vdd.n1452 vdd.n1082 185
R18527 vdd.n2567 vdd.n1082 185
R18528 vdd.n1454 vdd.n1453 185
R18529 vdd.n1453 vdd.n1080 185
R18530 vdd.n1455 vdd.n1089 185
R18531 vdd.n2561 vdd.n1089 185
R18532 vdd.n1457 vdd.n1456 185
R18533 vdd.n1456 vdd.n1087 185
R18534 vdd.n1458 vdd.n1095 185
R18535 vdd.n2555 vdd.n1095 185
R18536 vdd.n1460 vdd.n1459 185
R18537 vdd.n1459 vdd.n1093 185
R18538 vdd.n1461 vdd.n1100 185
R18539 vdd.n2549 vdd.n1100 185
R18540 vdd.n1463 vdd.n1462 185
R18541 vdd.n1462 vdd.n1106 185
R18542 vdd.n1464 vdd.n1105 185
R18543 vdd.n2543 vdd.n1105 185
R18544 vdd.n1466 vdd.n1465 185
R18545 vdd.n1465 vdd.n1112 185
R18546 vdd.n1467 vdd.n1111 185
R18547 vdd.n2537 vdd.n1111 185
R18548 vdd.n1469 vdd.n1468 185
R18549 vdd.n1468 vdd.n1119 185
R18550 vdd.n1470 vdd.n1118 185
R18551 vdd.n2531 vdd.n1118 185
R18552 vdd.n1472 vdd.n1471 185
R18553 vdd.n1471 vdd.n1116 185
R18554 vdd.n1473 vdd.n1125 185
R18555 vdd.n2525 vdd.n1125 185
R18556 vdd.n1475 vdd.n1474 185
R18557 vdd.n1474 vdd.n1123 185
R18558 vdd.n1476 vdd.n1130 185
R18559 vdd.n2519 vdd.n1130 185
R18560 vdd.n1478 vdd.n1477 185
R18561 vdd.n1477 vdd.n1137 185
R18562 vdd.n1479 vdd.n1136 185
R18563 vdd.n2513 vdd.n1136 185
R18564 vdd.n1481 vdd.n1480 185
R18565 vdd.n1480 vdd.n1134 185
R18566 vdd.n1281 vdd.n1280 185
R18567 vdd.n1283 vdd.n1282 185
R18568 vdd.n1285 vdd.n1284 185
R18569 vdd.n1287 vdd.n1286 185
R18570 vdd.n1289 vdd.n1288 185
R18571 vdd.n1291 vdd.n1290 185
R18572 vdd.n1293 vdd.n1292 185
R18573 vdd.n1295 vdd.n1294 185
R18574 vdd.n1297 vdd.n1296 185
R18575 vdd.n1299 vdd.n1298 185
R18576 vdd.n1301 vdd.n1300 185
R18577 vdd.n1303 vdd.n1302 185
R18578 vdd.n1305 vdd.n1304 185
R18579 vdd.n1307 vdd.n1306 185
R18580 vdd.n1309 vdd.n1308 185
R18581 vdd.n1311 vdd.n1310 185
R18582 vdd.n1313 vdd.n1312 185
R18583 vdd.n1515 vdd.n1314 185
R18584 vdd.n1514 vdd.n1513 185
R18585 vdd.n1512 vdd.n1511 185
R18586 vdd.n1510 vdd.n1509 185
R18587 vdd.n1508 vdd.n1507 185
R18588 vdd.n1506 vdd.n1505 185
R18589 vdd.n1504 vdd.n1503 185
R18590 vdd.n1502 vdd.n1501 185
R18591 vdd.n1500 vdd.n1499 185
R18592 vdd.n1498 vdd.n1497 185
R18593 vdd.n1496 vdd.n1495 185
R18594 vdd.n1494 vdd.n1493 185
R18595 vdd.n1492 vdd.n1491 185
R18596 vdd.n1490 vdd.n1489 185
R18597 vdd.n1488 vdd.n1487 185
R18598 vdd.n1486 vdd.n1485 185
R18599 vdd.n1484 vdd.n1483 185
R18600 vdd.n1482 vdd.n1175 185
R18601 vdd.n2506 vdd.n1175 185
R18602 vdd.n327 vdd.n326 171.744
R18603 vdd.n326 vdd.n325 171.744
R18604 vdd.n325 vdd.n294 171.744
R18605 vdd.n318 vdd.n294 171.744
R18606 vdd.n318 vdd.n317 171.744
R18607 vdd.n317 vdd.n299 171.744
R18608 vdd.n310 vdd.n299 171.744
R18609 vdd.n310 vdd.n309 171.744
R18610 vdd.n309 vdd.n303 171.744
R18611 vdd.n268 vdd.n267 171.744
R18612 vdd.n267 vdd.n266 171.744
R18613 vdd.n266 vdd.n235 171.744
R18614 vdd.n259 vdd.n235 171.744
R18615 vdd.n259 vdd.n258 171.744
R18616 vdd.n258 vdd.n240 171.744
R18617 vdd.n251 vdd.n240 171.744
R18618 vdd.n251 vdd.n250 171.744
R18619 vdd.n250 vdd.n244 171.744
R18620 vdd.n225 vdd.n224 171.744
R18621 vdd.n224 vdd.n223 171.744
R18622 vdd.n223 vdd.n192 171.744
R18623 vdd.n216 vdd.n192 171.744
R18624 vdd.n216 vdd.n215 171.744
R18625 vdd.n215 vdd.n197 171.744
R18626 vdd.n208 vdd.n197 171.744
R18627 vdd.n208 vdd.n207 171.744
R18628 vdd.n207 vdd.n201 171.744
R18629 vdd.n166 vdd.n165 171.744
R18630 vdd.n165 vdd.n164 171.744
R18631 vdd.n164 vdd.n133 171.744
R18632 vdd.n157 vdd.n133 171.744
R18633 vdd.n157 vdd.n156 171.744
R18634 vdd.n156 vdd.n138 171.744
R18635 vdd.n149 vdd.n138 171.744
R18636 vdd.n149 vdd.n148 171.744
R18637 vdd.n148 vdd.n142 171.744
R18638 vdd.n124 vdd.n123 171.744
R18639 vdd.n123 vdd.n122 171.744
R18640 vdd.n122 vdd.n91 171.744
R18641 vdd.n115 vdd.n91 171.744
R18642 vdd.n115 vdd.n114 171.744
R18643 vdd.n114 vdd.n96 171.744
R18644 vdd.n107 vdd.n96 171.744
R18645 vdd.n107 vdd.n106 171.744
R18646 vdd.n106 vdd.n100 171.744
R18647 vdd.n65 vdd.n64 171.744
R18648 vdd.n64 vdd.n63 171.744
R18649 vdd.n63 vdd.n32 171.744
R18650 vdd.n56 vdd.n32 171.744
R18651 vdd.n56 vdd.n55 171.744
R18652 vdd.n55 vdd.n37 171.744
R18653 vdd.n48 vdd.n37 171.744
R18654 vdd.n48 vdd.n47 171.744
R18655 vdd.n47 vdd.n41 171.744
R18656 vdd.n2201 vdd.n2200 171.744
R18657 vdd.n2200 vdd.n2199 171.744
R18658 vdd.n2199 vdd.n2168 171.744
R18659 vdd.n2192 vdd.n2168 171.744
R18660 vdd.n2192 vdd.n2191 171.744
R18661 vdd.n2191 vdd.n2173 171.744
R18662 vdd.n2184 vdd.n2173 171.744
R18663 vdd.n2184 vdd.n2183 171.744
R18664 vdd.n2183 vdd.n2177 171.744
R18665 vdd.n2260 vdd.n2259 171.744
R18666 vdd.n2259 vdd.n2258 171.744
R18667 vdd.n2258 vdd.n2227 171.744
R18668 vdd.n2251 vdd.n2227 171.744
R18669 vdd.n2251 vdd.n2250 171.744
R18670 vdd.n2250 vdd.n2232 171.744
R18671 vdd.n2243 vdd.n2232 171.744
R18672 vdd.n2243 vdd.n2242 171.744
R18673 vdd.n2242 vdd.n2236 171.744
R18674 vdd.n2099 vdd.n2098 171.744
R18675 vdd.n2098 vdd.n2097 171.744
R18676 vdd.n2097 vdd.n2066 171.744
R18677 vdd.n2090 vdd.n2066 171.744
R18678 vdd.n2090 vdd.n2089 171.744
R18679 vdd.n2089 vdd.n2071 171.744
R18680 vdd.n2082 vdd.n2071 171.744
R18681 vdd.n2082 vdd.n2081 171.744
R18682 vdd.n2081 vdd.n2075 171.744
R18683 vdd.n2158 vdd.n2157 171.744
R18684 vdd.n2157 vdd.n2156 171.744
R18685 vdd.n2156 vdd.n2125 171.744
R18686 vdd.n2149 vdd.n2125 171.744
R18687 vdd.n2149 vdd.n2148 171.744
R18688 vdd.n2148 vdd.n2130 171.744
R18689 vdd.n2141 vdd.n2130 171.744
R18690 vdd.n2141 vdd.n2140 171.744
R18691 vdd.n2140 vdd.n2134 171.744
R18692 vdd.n1998 vdd.n1997 171.744
R18693 vdd.n1997 vdd.n1996 171.744
R18694 vdd.n1996 vdd.n1965 171.744
R18695 vdd.n1989 vdd.n1965 171.744
R18696 vdd.n1989 vdd.n1988 171.744
R18697 vdd.n1988 vdd.n1970 171.744
R18698 vdd.n1981 vdd.n1970 171.744
R18699 vdd.n1981 vdd.n1980 171.744
R18700 vdd.n1980 vdd.n1974 171.744
R18701 vdd.n2057 vdd.n2056 171.744
R18702 vdd.n2056 vdd.n2055 171.744
R18703 vdd.n2055 vdd.n2024 171.744
R18704 vdd.n2048 vdd.n2024 171.744
R18705 vdd.n2048 vdd.n2047 171.744
R18706 vdd.n2047 vdd.n2029 171.744
R18707 vdd.n2040 vdd.n2029 171.744
R18708 vdd.n2040 vdd.n2039 171.744
R18709 vdd.n2039 vdd.n2033 171.744
R18710 vdd.n468 vdd.n467 146.341
R18711 vdd.n474 vdd.n473 146.341
R18712 vdd.n478 vdd.n477 146.341
R18713 vdd.n484 vdd.n483 146.341
R18714 vdd.n488 vdd.n487 146.341
R18715 vdd.n494 vdd.n493 146.341
R18716 vdd.n498 vdd.n497 146.341
R18717 vdd.n504 vdd.n503 146.341
R18718 vdd.n508 vdd.n507 146.341
R18719 vdd.n514 vdd.n513 146.341
R18720 vdd.n518 vdd.n517 146.341
R18721 vdd.n524 vdd.n523 146.341
R18722 vdd.n528 vdd.n527 146.341
R18723 vdd.n534 vdd.n533 146.341
R18724 vdd.n538 vdd.n537 146.341
R18725 vdd.n544 vdd.n543 146.341
R18726 vdd.n548 vdd.n547 146.341
R18727 vdd.n554 vdd.n553 146.341
R18728 vdd.n558 vdd.n557 146.341
R18729 vdd.n564 vdd.n563 146.341
R18730 vdd.n568 vdd.n567 146.341
R18731 vdd.n574 vdd.n573 146.341
R18732 vdd.n578 vdd.n577 146.341
R18733 vdd.n584 vdd.n583 146.341
R18734 vdd.n588 vdd.n587 146.341
R18735 vdd.n594 vdd.n593 146.341
R18736 vdd.n598 vdd.n597 146.341
R18737 vdd.n604 vdd.n603 146.341
R18738 vdd.n608 vdd.n607 146.341
R18739 vdd.n614 vdd.n613 146.341
R18740 vdd.n616 vdd.n425 146.341
R18741 vdd.n3502 vdd.n685 146.341
R18742 vdd.n3502 vdd.n677 146.341
R18743 vdd.n3512 vdd.n677 146.341
R18744 vdd.n3512 vdd.n673 146.341
R18745 vdd.n3518 vdd.n673 146.341
R18746 vdd.n3518 vdd.n667 146.341
R18747 vdd.n3529 vdd.n667 146.341
R18748 vdd.n3529 vdd.n663 146.341
R18749 vdd.n3535 vdd.n663 146.341
R18750 vdd.n3535 vdd.n654 146.341
R18751 vdd.n3545 vdd.n654 146.341
R18752 vdd.n3545 vdd.n650 146.341
R18753 vdd.n3551 vdd.n650 146.341
R18754 vdd.n3551 vdd.n643 146.341
R18755 vdd.n3562 vdd.n643 146.341
R18756 vdd.n3562 vdd.n639 146.341
R18757 vdd.n3571 vdd.n639 146.341
R18758 vdd.n3571 vdd.n632 146.341
R18759 vdd.n3581 vdd.n632 146.341
R18760 vdd.n3582 vdd.n3581 146.341
R18761 vdd.n3582 vdd.n341 146.341
R18762 vdd.n342 vdd.n341 146.341
R18763 vdd.n343 vdd.n342 146.341
R18764 vdd.n3589 vdd.n343 146.341
R18765 vdd.n3589 vdd.n351 146.341
R18766 vdd.n352 vdd.n351 146.341
R18767 vdd.n353 vdd.n352 146.341
R18768 vdd.n3596 vdd.n353 146.341
R18769 vdd.n3596 vdd.n362 146.341
R18770 vdd.n363 vdd.n362 146.341
R18771 vdd.n364 vdd.n363 146.341
R18772 vdd.n3604 vdd.n364 146.341
R18773 vdd.n3604 vdd.n372 146.341
R18774 vdd.n373 vdd.n372 146.341
R18775 vdd.n374 vdd.n373 146.341
R18776 vdd.n3611 vdd.n374 146.341
R18777 vdd.n3611 vdd.n383 146.341
R18778 vdd.n384 vdd.n383 146.341
R18779 vdd.n385 vdd.n384 146.341
R18780 vdd.n3618 vdd.n385 146.341
R18781 vdd.n3618 vdd.n393 146.341
R18782 vdd.n725 vdd.n724 146.341
R18783 vdd.n728 vdd.n724 146.341
R18784 vdd.n734 vdd.n733 146.341
R18785 vdd.n3484 vdd.n3483 146.341
R18786 vdd.n3480 vdd.n3479 146.341
R18787 vdd.n3476 vdd.n3475 146.341
R18788 vdd.n3472 vdd.n3471 146.341
R18789 vdd.n3468 vdd.n3467 146.341
R18790 vdd.n3464 vdd.n3463 146.341
R18791 vdd.n3460 vdd.n3459 146.341
R18792 vdd.n3451 vdd.n3450 146.341
R18793 vdd.n3448 vdd.n3447 146.341
R18794 vdd.n3444 vdd.n3443 146.341
R18795 vdd.n3440 vdd.n3439 146.341
R18796 vdd.n3436 vdd.n3435 146.341
R18797 vdd.n3432 vdd.n3431 146.341
R18798 vdd.n3428 vdd.n3427 146.341
R18799 vdd.n3424 vdd.n3423 146.341
R18800 vdd.n3420 vdd.n3419 146.341
R18801 vdd.n3416 vdd.n3415 146.341
R18802 vdd.n3412 vdd.n3411 146.341
R18803 vdd.n3405 vdd.n3404 146.341
R18804 vdd.n3402 vdd.n3401 146.341
R18805 vdd.n3398 vdd.n3397 146.341
R18806 vdd.n3394 vdd.n3393 146.341
R18807 vdd.n3390 vdd.n3389 146.341
R18808 vdd.n3386 vdd.n3385 146.341
R18809 vdd.n3382 vdd.n3381 146.341
R18810 vdd.n3378 vdd.n3377 146.341
R18811 vdd.n3374 vdd.n3373 146.341
R18812 vdd.n3370 vdd.n3369 146.341
R18813 vdd.n3496 vdd.n691 146.341
R18814 vdd.n3504 vdd.n684 146.341
R18815 vdd.n3504 vdd.n680 146.341
R18816 vdd.n3510 vdd.n680 146.341
R18817 vdd.n3510 vdd.n672 146.341
R18818 vdd.n3521 vdd.n672 146.341
R18819 vdd.n3521 vdd.n668 146.341
R18820 vdd.n3527 vdd.n668 146.341
R18821 vdd.n3527 vdd.n661 146.341
R18822 vdd.n3537 vdd.n661 146.341
R18823 vdd.n3537 vdd.n657 146.341
R18824 vdd.n3543 vdd.n657 146.341
R18825 vdd.n3543 vdd.n649 146.341
R18826 vdd.n3554 vdd.n649 146.341
R18827 vdd.n3554 vdd.n645 146.341
R18828 vdd.n3560 vdd.n645 146.341
R18829 vdd.n3560 vdd.n638 146.341
R18830 vdd.n3573 vdd.n638 146.341
R18831 vdd.n3573 vdd.n634 146.341
R18832 vdd.n3579 vdd.n634 146.341
R18833 vdd.n3579 vdd.n338 146.341
R18834 vdd.n3668 vdd.n338 146.341
R18835 vdd.n3668 vdd.n339 146.341
R18836 vdd.n3664 vdd.n339 146.341
R18837 vdd.n3664 vdd.n345 146.341
R18838 vdd.n3660 vdd.n345 146.341
R18839 vdd.n3660 vdd.n350 146.341
R18840 vdd.n3656 vdd.n350 146.341
R18841 vdd.n3656 vdd.n354 146.341
R18842 vdd.n3652 vdd.n354 146.341
R18843 vdd.n3652 vdd.n360 146.341
R18844 vdd.n3648 vdd.n360 146.341
R18845 vdd.n3648 vdd.n365 146.341
R18846 vdd.n3644 vdd.n365 146.341
R18847 vdd.n3644 vdd.n371 146.341
R18848 vdd.n3640 vdd.n371 146.341
R18849 vdd.n3640 vdd.n376 146.341
R18850 vdd.n3636 vdd.n376 146.341
R18851 vdd.n3636 vdd.n382 146.341
R18852 vdd.n3632 vdd.n382 146.341
R18853 vdd.n3632 vdd.n387 146.341
R18854 vdd.n3628 vdd.n387 146.341
R18855 vdd.n2471 vdd.n2470 146.341
R18856 vdd.n2468 vdd.n2465 146.341
R18857 vdd.n2463 vdd.n1185 146.341
R18858 vdd.n2459 vdd.n2458 146.341
R18859 vdd.n2456 vdd.n1189 146.341
R18860 vdd.n2452 vdd.n2451 146.341
R18861 vdd.n2449 vdd.n1196 146.341
R18862 vdd.n2445 vdd.n2444 146.341
R18863 vdd.n2442 vdd.n1203 146.341
R18864 vdd.n1214 vdd.n1211 146.341
R18865 vdd.n2434 vdd.n2433 146.341
R18866 vdd.n2431 vdd.n1216 146.341
R18867 vdd.n2427 vdd.n2426 146.341
R18868 vdd.n2424 vdd.n1222 146.341
R18869 vdd.n2420 vdd.n2419 146.341
R18870 vdd.n2417 vdd.n1229 146.341
R18871 vdd.n2413 vdd.n2412 146.341
R18872 vdd.n2410 vdd.n1236 146.341
R18873 vdd.n2406 vdd.n2405 146.341
R18874 vdd.n2403 vdd.n1243 146.341
R18875 vdd.n1254 vdd.n1251 146.341
R18876 vdd.n2395 vdd.n2394 146.341
R18877 vdd.n2392 vdd.n1256 146.341
R18878 vdd.n2388 vdd.n2387 146.341
R18879 vdd.n2385 vdd.n1262 146.341
R18880 vdd.n2381 vdd.n2380 146.341
R18881 vdd.n2378 vdd.n1269 146.341
R18882 vdd.n2374 vdd.n2373 146.341
R18883 vdd.n2371 vdd.n1276 146.341
R18884 vdd.n1522 vdd.n1520 146.341
R18885 vdd.n1525 vdd.n1524 146.341
R18886 vdd.n1883 vdd.n1643 146.341
R18887 vdd.n1883 vdd.n1639 146.341
R18888 vdd.n1889 vdd.n1639 146.341
R18889 vdd.n1889 vdd.n1631 146.341
R18890 vdd.n1900 vdd.n1631 146.341
R18891 vdd.n1900 vdd.n1627 146.341
R18892 vdd.n1906 vdd.n1627 146.341
R18893 vdd.n1906 vdd.n1621 146.341
R18894 vdd.n1917 vdd.n1621 146.341
R18895 vdd.n1917 vdd.n1617 146.341
R18896 vdd.n1923 vdd.n1617 146.341
R18897 vdd.n1923 vdd.n1608 146.341
R18898 vdd.n1933 vdd.n1608 146.341
R18899 vdd.n1933 vdd.n1604 146.341
R18900 vdd.n1939 vdd.n1604 146.341
R18901 vdd.n1939 vdd.n1597 146.341
R18902 vdd.n1950 vdd.n1597 146.341
R18903 vdd.n1950 vdd.n1593 146.341
R18904 vdd.n1956 vdd.n1593 146.341
R18905 vdd.n1956 vdd.n1586 146.341
R18906 vdd.n2273 vdd.n1586 146.341
R18907 vdd.n2273 vdd.n1582 146.341
R18908 vdd.n2279 vdd.n1582 146.341
R18909 vdd.n2279 vdd.n1574 146.341
R18910 vdd.n2290 vdd.n1574 146.341
R18911 vdd.n2290 vdd.n1570 146.341
R18912 vdd.n2296 vdd.n1570 146.341
R18913 vdd.n2296 vdd.n1564 146.341
R18914 vdd.n2307 vdd.n1564 146.341
R18915 vdd.n2307 vdd.n1560 146.341
R18916 vdd.n2313 vdd.n1560 146.341
R18917 vdd.n2313 vdd.n1551 146.341
R18918 vdd.n2323 vdd.n1551 146.341
R18919 vdd.n2323 vdd.n1547 146.341
R18920 vdd.n2329 vdd.n1547 146.341
R18921 vdd.n2329 vdd.n1541 146.341
R18922 vdd.n2340 vdd.n1541 146.341
R18923 vdd.n2340 vdd.n1536 146.341
R18924 vdd.n2348 vdd.n1536 146.341
R18925 vdd.n2348 vdd.n1527 146.341
R18926 vdd.n2359 vdd.n1527 146.341
R18927 vdd.n1872 vdd.n1648 146.341
R18928 vdd.n1872 vdd.n1681 146.341
R18929 vdd.n1685 vdd.n1684 146.341
R18930 vdd.n1687 vdd.n1686 146.341
R18931 vdd.n1691 vdd.n1690 146.341
R18932 vdd.n1693 vdd.n1692 146.341
R18933 vdd.n1697 vdd.n1696 146.341
R18934 vdd.n1699 vdd.n1698 146.341
R18935 vdd.n1703 vdd.n1702 146.341
R18936 vdd.n1705 vdd.n1704 146.341
R18937 vdd.n1711 vdd.n1710 146.341
R18938 vdd.n1713 vdd.n1712 146.341
R18939 vdd.n1717 vdd.n1716 146.341
R18940 vdd.n1719 vdd.n1718 146.341
R18941 vdd.n1723 vdd.n1722 146.341
R18942 vdd.n1725 vdd.n1724 146.341
R18943 vdd.n1729 vdd.n1728 146.341
R18944 vdd.n1731 vdd.n1730 146.341
R18945 vdd.n1735 vdd.n1734 146.341
R18946 vdd.n1737 vdd.n1736 146.341
R18947 vdd.n1809 vdd.n1740 146.341
R18948 vdd.n1742 vdd.n1741 146.341
R18949 vdd.n1746 vdd.n1745 146.341
R18950 vdd.n1748 vdd.n1747 146.341
R18951 vdd.n1752 vdd.n1751 146.341
R18952 vdd.n1754 vdd.n1753 146.341
R18953 vdd.n1758 vdd.n1757 146.341
R18954 vdd.n1760 vdd.n1759 146.341
R18955 vdd.n1764 vdd.n1763 146.341
R18956 vdd.n1766 vdd.n1765 146.341
R18957 vdd.n1770 vdd.n1769 146.341
R18958 vdd.n1771 vdd.n1679 146.341
R18959 vdd.n1881 vdd.n1644 146.341
R18960 vdd.n1881 vdd.n1637 146.341
R18961 vdd.n1892 vdd.n1637 146.341
R18962 vdd.n1892 vdd.n1633 146.341
R18963 vdd.n1898 vdd.n1633 146.341
R18964 vdd.n1898 vdd.n1626 146.341
R18965 vdd.n1909 vdd.n1626 146.341
R18966 vdd.n1909 vdd.n1622 146.341
R18967 vdd.n1915 vdd.n1622 146.341
R18968 vdd.n1915 vdd.n1615 146.341
R18969 vdd.n1925 vdd.n1615 146.341
R18970 vdd.n1925 vdd.n1611 146.341
R18971 vdd.n1931 vdd.n1611 146.341
R18972 vdd.n1931 vdd.n1603 146.341
R18973 vdd.n1942 vdd.n1603 146.341
R18974 vdd.n1942 vdd.n1599 146.341
R18975 vdd.n1948 vdd.n1599 146.341
R18976 vdd.n1948 vdd.n1592 146.341
R18977 vdd.n1958 vdd.n1592 146.341
R18978 vdd.n1958 vdd.n1588 146.341
R18979 vdd.n2271 vdd.n1588 146.341
R18980 vdd.n2271 vdd.n1580 146.341
R18981 vdd.n2282 vdd.n1580 146.341
R18982 vdd.n2282 vdd.n1576 146.341
R18983 vdd.n2288 vdd.n1576 146.341
R18984 vdd.n2288 vdd.n1569 146.341
R18985 vdd.n2299 vdd.n1569 146.341
R18986 vdd.n2299 vdd.n1565 146.341
R18987 vdd.n2305 vdd.n1565 146.341
R18988 vdd.n2305 vdd.n1558 146.341
R18989 vdd.n2315 vdd.n1558 146.341
R18990 vdd.n2315 vdd.n1554 146.341
R18991 vdd.n2321 vdd.n1554 146.341
R18992 vdd.n2321 vdd.n1546 146.341
R18993 vdd.n2332 vdd.n1546 146.341
R18994 vdd.n2332 vdd.n1542 146.341
R18995 vdd.n2338 vdd.n1542 146.341
R18996 vdd.n2338 vdd.n1534 146.341
R18997 vdd.n2351 vdd.n1534 146.341
R18998 vdd.n2351 vdd.n1529 146.341
R18999 vdd.n2357 vdd.n1529 146.341
R19000 vdd.n1315 vdd.t167 127.284
R19001 vdd.n1010 vdd.t207 127.284
R19002 vdd.n1319 vdd.t204 127.284
R19003 vdd.n1001 vdd.t228 127.284
R19004 vdd.n896 vdd.t191 127.284
R19005 vdd.n896 vdd.t192 127.284
R19006 vdd.n2823 vdd.t222 127.284
R19007 vdd.n832 vdd.t183 127.284
R19008 vdd.n2820 vdd.t215 127.284
R19009 vdd.n799 vdd.t162 127.284
R19010 vdd.n1071 vdd.t218 127.284
R19011 vdd.n1071 vdd.t219 127.284
R19012 vdd.n22 vdd.n20 117.314
R19013 vdd.n17 vdd.n15 117.314
R19014 vdd.n27 vdd.n26 116.927
R19015 vdd.n24 vdd.n23 116.927
R19016 vdd.n22 vdd.n21 116.927
R19017 vdd.n17 vdd.n16 116.927
R19018 vdd.n19 vdd.n18 116.927
R19019 vdd.n27 vdd.n25 116.927
R19020 vdd.n1316 vdd.t166 111.188
R19021 vdd.n1011 vdd.t208 111.188
R19022 vdd.n1320 vdd.t203 111.188
R19023 vdd.n1002 vdd.t229 111.188
R19024 vdd.n2824 vdd.t221 111.188
R19025 vdd.n833 vdd.t184 111.188
R19026 vdd.n2821 vdd.t214 111.188
R19027 vdd.n800 vdd.t163 111.188
R19028 vdd.n3094 vdd.n960 99.5127
R19029 vdd.n3094 vdd.n951 99.5127
R19030 vdd.n3102 vdd.n951 99.5127
R19031 vdd.n3102 vdd.n949 99.5127
R19032 vdd.n3106 vdd.n949 99.5127
R19033 vdd.n3106 vdd.n939 99.5127
R19034 vdd.n3114 vdd.n939 99.5127
R19035 vdd.n3114 vdd.n937 99.5127
R19036 vdd.n3118 vdd.n937 99.5127
R19037 vdd.n3118 vdd.n928 99.5127
R19038 vdd.n3126 vdd.n928 99.5127
R19039 vdd.n3126 vdd.n926 99.5127
R19040 vdd.n3130 vdd.n926 99.5127
R19041 vdd.n3130 vdd.n917 99.5127
R19042 vdd.n3138 vdd.n917 99.5127
R19043 vdd.n3138 vdd.n915 99.5127
R19044 vdd.n3142 vdd.n915 99.5127
R19045 vdd.n3142 vdd.n904 99.5127
R19046 vdd.n3151 vdd.n904 99.5127
R19047 vdd.n3151 vdd.n902 99.5127
R19048 vdd.n3155 vdd.n902 99.5127
R19049 vdd.n3155 vdd.n892 99.5127
R19050 vdd.n3163 vdd.n892 99.5127
R19051 vdd.n3163 vdd.n890 99.5127
R19052 vdd.n3167 vdd.n890 99.5127
R19053 vdd.n3167 vdd.n880 99.5127
R19054 vdd.n3175 vdd.n880 99.5127
R19055 vdd.n3175 vdd.n878 99.5127
R19056 vdd.n3179 vdd.n878 99.5127
R19057 vdd.n3179 vdd.n867 99.5127
R19058 vdd.n3187 vdd.n867 99.5127
R19059 vdd.n3187 vdd.n865 99.5127
R19060 vdd.n3191 vdd.n865 99.5127
R19061 vdd.n3191 vdd.n856 99.5127
R19062 vdd.n3199 vdd.n856 99.5127
R19063 vdd.n3199 vdd.n854 99.5127
R19064 vdd.n3203 vdd.n854 99.5127
R19065 vdd.n3203 vdd.n842 99.5127
R19066 vdd.n3256 vdd.n842 99.5127
R19067 vdd.n3256 vdd.n840 99.5127
R19068 vdd.n3260 vdd.n840 99.5127
R19069 vdd.n3260 vdd.n808 99.5127
R19070 vdd.n3330 vdd.n808 99.5127
R19071 vdd.n3326 vdd.n809 99.5127
R19072 vdd.n3324 vdd.n3323 99.5127
R19073 vdd.n3321 vdd.n813 99.5127
R19074 vdd.n3317 vdd.n3316 99.5127
R19075 vdd.n3314 vdd.n816 99.5127
R19076 vdd.n3310 vdd.n3309 99.5127
R19077 vdd.n3307 vdd.n819 99.5127
R19078 vdd.n3303 vdd.n3302 99.5127
R19079 vdd.n3300 vdd.n3298 99.5127
R19080 vdd.n3296 vdd.n822 99.5127
R19081 vdd.n3292 vdd.n3291 99.5127
R19082 vdd.n3289 vdd.n825 99.5127
R19083 vdd.n3285 vdd.n3284 99.5127
R19084 vdd.n3282 vdd.n828 99.5127
R19085 vdd.n3278 vdd.n3277 99.5127
R19086 vdd.n3275 vdd.n831 99.5127
R19087 vdd.n3270 vdd.n3269 99.5127
R19088 vdd.n3021 vdd.n958 99.5127
R19089 vdd.n3017 vdd.n958 99.5127
R19090 vdd.n3017 vdd.n952 99.5127
R19091 vdd.n2899 vdd.n952 99.5127
R19092 vdd.n2899 vdd.n947 99.5127
R19093 vdd.n2902 vdd.n947 99.5127
R19094 vdd.n2902 vdd.n941 99.5127
R19095 vdd.n3003 vdd.n941 99.5127
R19096 vdd.n3003 vdd.n935 99.5127
R19097 vdd.n2999 vdd.n935 99.5127
R19098 vdd.n2999 vdd.n929 99.5127
R19099 vdd.n2946 vdd.n929 99.5127
R19100 vdd.n2946 vdd.n923 99.5127
R19101 vdd.n2943 vdd.n923 99.5127
R19102 vdd.n2943 vdd.n918 99.5127
R19103 vdd.n2940 vdd.n918 99.5127
R19104 vdd.n2940 vdd.n913 99.5127
R19105 vdd.n2937 vdd.n913 99.5127
R19106 vdd.n2937 vdd.n906 99.5127
R19107 vdd.n2934 vdd.n906 99.5127
R19108 vdd.n2934 vdd.n899 99.5127
R19109 vdd.n2931 vdd.n899 99.5127
R19110 vdd.n2931 vdd.n893 99.5127
R19111 vdd.n2928 vdd.n893 99.5127
R19112 vdd.n2928 vdd.n888 99.5127
R19113 vdd.n2925 vdd.n888 99.5127
R19114 vdd.n2925 vdd.n882 99.5127
R19115 vdd.n2922 vdd.n882 99.5127
R19116 vdd.n2922 vdd.n875 99.5127
R19117 vdd.n2919 vdd.n875 99.5127
R19118 vdd.n2919 vdd.n868 99.5127
R19119 vdd.n2916 vdd.n868 99.5127
R19120 vdd.n2916 vdd.n862 99.5127
R19121 vdd.n2913 vdd.n862 99.5127
R19122 vdd.n2913 vdd.n857 99.5127
R19123 vdd.n2910 vdd.n857 99.5127
R19124 vdd.n2910 vdd.n852 99.5127
R19125 vdd.n2907 vdd.n852 99.5127
R19126 vdd.n2907 vdd.n844 99.5127
R19127 vdd.n844 vdd.n837 99.5127
R19128 vdd.n3262 vdd.n837 99.5127
R19129 vdd.n3263 vdd.n3262 99.5127
R19130 vdd.n3263 vdd.n806 99.5127
R19131 vdd.n3087 vdd.n962 99.5127
R19132 vdd.n3087 vdd.n2819 99.5127
R19133 vdd.n3083 vdd.n3082 99.5127
R19134 vdd.n3079 vdd.n3078 99.5127
R19135 vdd.n3075 vdd.n3074 99.5127
R19136 vdd.n3071 vdd.n3070 99.5127
R19137 vdd.n3067 vdd.n3066 99.5127
R19138 vdd.n3063 vdd.n3062 99.5127
R19139 vdd.n3059 vdd.n3058 99.5127
R19140 vdd.n3055 vdd.n3054 99.5127
R19141 vdd.n3051 vdd.n3050 99.5127
R19142 vdd.n3047 vdd.n3046 99.5127
R19143 vdd.n3043 vdd.n3042 99.5127
R19144 vdd.n3039 vdd.n3038 99.5127
R19145 vdd.n3035 vdd.n3034 99.5127
R19146 vdd.n3031 vdd.n3030 99.5127
R19147 vdd.n3026 vdd.n3025 99.5127
R19148 vdd.n2783 vdd.n999 99.5127
R19149 vdd.n2779 vdd.n2778 99.5127
R19150 vdd.n2775 vdd.n2774 99.5127
R19151 vdd.n2771 vdd.n2770 99.5127
R19152 vdd.n2767 vdd.n2766 99.5127
R19153 vdd.n2763 vdd.n2762 99.5127
R19154 vdd.n2759 vdd.n2758 99.5127
R19155 vdd.n2755 vdd.n2754 99.5127
R19156 vdd.n2751 vdd.n2750 99.5127
R19157 vdd.n2747 vdd.n2746 99.5127
R19158 vdd.n2743 vdd.n2742 99.5127
R19159 vdd.n2739 vdd.n2738 99.5127
R19160 vdd.n2735 vdd.n2734 99.5127
R19161 vdd.n2731 vdd.n2730 99.5127
R19162 vdd.n2727 vdd.n2726 99.5127
R19163 vdd.n2723 vdd.n2722 99.5127
R19164 vdd.n2718 vdd.n2717 99.5127
R19165 vdd.n1355 vdd.n1135 99.5127
R19166 vdd.n1358 vdd.n1135 99.5127
R19167 vdd.n1358 vdd.n1129 99.5127
R19168 vdd.n1361 vdd.n1129 99.5127
R19169 vdd.n1361 vdd.n1124 99.5127
R19170 vdd.n1364 vdd.n1124 99.5127
R19171 vdd.n1364 vdd.n1117 99.5127
R19172 vdd.n1367 vdd.n1117 99.5127
R19173 vdd.n1367 vdd.n1110 99.5127
R19174 vdd.n1370 vdd.n1110 99.5127
R19175 vdd.n1370 vdd.n1104 99.5127
R19176 vdd.n1373 vdd.n1104 99.5127
R19177 vdd.n1373 vdd.n1099 99.5127
R19178 vdd.n1376 vdd.n1099 99.5127
R19179 vdd.n1376 vdd.n1094 99.5127
R19180 vdd.n1379 vdd.n1094 99.5127
R19181 vdd.n1379 vdd.n1088 99.5127
R19182 vdd.n1382 vdd.n1088 99.5127
R19183 vdd.n1382 vdd.n1081 99.5127
R19184 vdd.n1385 vdd.n1081 99.5127
R19185 vdd.n1385 vdd.n1074 99.5127
R19186 vdd.n1388 vdd.n1074 99.5127
R19187 vdd.n1388 vdd.n1068 99.5127
R19188 vdd.n1391 vdd.n1068 99.5127
R19189 vdd.n1391 vdd.n1063 99.5127
R19190 vdd.n1394 vdd.n1063 99.5127
R19191 vdd.n1394 vdd.n1057 99.5127
R19192 vdd.n1436 vdd.n1057 99.5127
R19193 vdd.n1436 vdd.n1050 99.5127
R19194 vdd.n1432 vdd.n1050 99.5127
R19195 vdd.n1432 vdd.n1044 99.5127
R19196 vdd.n1429 vdd.n1044 99.5127
R19197 vdd.n1429 vdd.n1039 99.5127
R19198 vdd.n1426 vdd.n1039 99.5127
R19199 vdd.n1426 vdd.n1034 99.5127
R19200 vdd.n1406 vdd.n1034 99.5127
R19201 vdd.n1406 vdd.n1029 99.5127
R19202 vdd.n1403 vdd.n1029 99.5127
R19203 vdd.n1403 vdd.n1022 99.5127
R19204 vdd.n1400 vdd.n1022 99.5127
R19205 vdd.n1400 vdd.n1015 99.5127
R19206 vdd.n1015 vdd.n1004 99.5127
R19207 vdd.n2713 vdd.n1004 99.5127
R19208 vdd.n2505 vdd.n1140 99.5127
R19209 vdd.n2505 vdd.n1176 99.5127
R19210 vdd.n2501 vdd.n2500 99.5127
R19211 vdd.n2497 vdd.n2496 99.5127
R19212 vdd.n2493 vdd.n2492 99.5127
R19213 vdd.n2489 vdd.n2488 99.5127
R19214 vdd.n2485 vdd.n2484 99.5127
R19215 vdd.n2481 vdd.n2480 99.5127
R19216 vdd.n2477 vdd.n2476 99.5127
R19217 vdd.n1322 vdd.n1321 99.5127
R19218 vdd.n1326 vdd.n1325 99.5127
R19219 vdd.n1330 vdd.n1329 99.5127
R19220 vdd.n1334 vdd.n1333 99.5127
R19221 vdd.n1338 vdd.n1337 99.5127
R19222 vdd.n1342 vdd.n1341 99.5127
R19223 vdd.n1346 vdd.n1345 99.5127
R19224 vdd.n1351 vdd.n1350 99.5127
R19225 vdd.n2512 vdd.n1138 99.5127
R19226 vdd.n2512 vdd.n1128 99.5127
R19227 vdd.n2520 vdd.n1128 99.5127
R19228 vdd.n2520 vdd.n1126 99.5127
R19229 vdd.n2524 vdd.n1126 99.5127
R19230 vdd.n2524 vdd.n1115 99.5127
R19231 vdd.n2532 vdd.n1115 99.5127
R19232 vdd.n2532 vdd.n1113 99.5127
R19233 vdd.n2536 vdd.n1113 99.5127
R19234 vdd.n2536 vdd.n1103 99.5127
R19235 vdd.n2544 vdd.n1103 99.5127
R19236 vdd.n2544 vdd.n1101 99.5127
R19237 vdd.n2548 vdd.n1101 99.5127
R19238 vdd.n2548 vdd.n1092 99.5127
R19239 vdd.n2556 vdd.n1092 99.5127
R19240 vdd.n2556 vdd.n1090 99.5127
R19241 vdd.n2560 vdd.n1090 99.5127
R19242 vdd.n2560 vdd.n1079 99.5127
R19243 vdd.n2568 vdd.n1079 99.5127
R19244 vdd.n2568 vdd.n1077 99.5127
R19245 vdd.n2572 vdd.n1077 99.5127
R19246 vdd.n2572 vdd.n1067 99.5127
R19247 vdd.n2581 vdd.n1067 99.5127
R19248 vdd.n2581 vdd.n1065 99.5127
R19249 vdd.n2585 vdd.n1065 99.5127
R19250 vdd.n2585 vdd.n1055 99.5127
R19251 vdd.n2593 vdd.n1055 99.5127
R19252 vdd.n2593 vdd.n1053 99.5127
R19253 vdd.n2597 vdd.n1053 99.5127
R19254 vdd.n2597 vdd.n1043 99.5127
R19255 vdd.n2605 vdd.n1043 99.5127
R19256 vdd.n2605 vdd.n1041 99.5127
R19257 vdd.n2609 vdd.n1041 99.5127
R19258 vdd.n2609 vdd.n1033 99.5127
R19259 vdd.n2617 vdd.n1033 99.5127
R19260 vdd.n2617 vdd.n1031 99.5127
R19261 vdd.n2621 vdd.n1031 99.5127
R19262 vdd.n2621 vdd.n1020 99.5127
R19263 vdd.n2631 vdd.n1020 99.5127
R19264 vdd.n2631 vdd.n1017 99.5127
R19265 vdd.n2636 vdd.n1017 99.5127
R19266 vdd.n2636 vdd.n1018 99.5127
R19267 vdd.n1018 vdd.n998 99.5127
R19268 vdd.n3246 vdd.n3245 99.5127
R19269 vdd.n3243 vdd.n3209 99.5127
R19270 vdd.n3239 vdd.n3238 99.5127
R19271 vdd.n3236 vdd.n3212 99.5127
R19272 vdd.n3232 vdd.n3231 99.5127
R19273 vdd.n3229 vdd.n3215 99.5127
R19274 vdd.n3225 vdd.n3224 99.5127
R19275 vdd.n3222 vdd.n3219 99.5127
R19276 vdd.n3363 vdd.n787 99.5127
R19277 vdd.n3361 vdd.n3360 99.5127
R19278 vdd.n3358 vdd.n789 99.5127
R19279 vdd.n3354 vdd.n3353 99.5127
R19280 vdd.n3351 vdd.n792 99.5127
R19281 vdd.n3347 vdd.n3346 99.5127
R19282 vdd.n3344 vdd.n795 99.5127
R19283 vdd.n3340 vdd.n3339 99.5127
R19284 vdd.n3337 vdd.n798 99.5127
R19285 vdd.n2895 vdd.n959 99.5127
R19286 vdd.n3015 vdd.n959 99.5127
R19287 vdd.n3015 vdd.n953 99.5127
R19288 vdd.n3011 vdd.n953 99.5127
R19289 vdd.n3011 vdd.n948 99.5127
R19290 vdd.n3008 vdd.n948 99.5127
R19291 vdd.n3008 vdd.n942 99.5127
R19292 vdd.n3005 vdd.n942 99.5127
R19293 vdd.n3005 vdd.n936 99.5127
R19294 vdd.n2997 vdd.n936 99.5127
R19295 vdd.n2997 vdd.n930 99.5127
R19296 vdd.n2993 vdd.n930 99.5127
R19297 vdd.n2993 vdd.n924 99.5127
R19298 vdd.n2990 vdd.n924 99.5127
R19299 vdd.n2990 vdd.n919 99.5127
R19300 vdd.n2987 vdd.n919 99.5127
R19301 vdd.n2987 vdd.n914 99.5127
R19302 vdd.n2984 vdd.n914 99.5127
R19303 vdd.n2984 vdd.n907 99.5127
R19304 vdd.n2981 vdd.n907 99.5127
R19305 vdd.n2981 vdd.n900 99.5127
R19306 vdd.n2978 vdd.n900 99.5127
R19307 vdd.n2978 vdd.n894 99.5127
R19308 vdd.n2975 vdd.n894 99.5127
R19309 vdd.n2975 vdd.n889 99.5127
R19310 vdd.n2972 vdd.n889 99.5127
R19311 vdd.n2972 vdd.n883 99.5127
R19312 vdd.n2969 vdd.n883 99.5127
R19313 vdd.n2969 vdd.n876 99.5127
R19314 vdd.n2966 vdd.n876 99.5127
R19315 vdd.n2966 vdd.n869 99.5127
R19316 vdd.n2963 vdd.n869 99.5127
R19317 vdd.n2963 vdd.n863 99.5127
R19318 vdd.n2960 vdd.n863 99.5127
R19319 vdd.n2960 vdd.n858 99.5127
R19320 vdd.n2957 vdd.n858 99.5127
R19321 vdd.n2957 vdd.n853 99.5127
R19322 vdd.n2954 vdd.n853 99.5127
R19323 vdd.n2954 vdd.n845 99.5127
R19324 vdd.n2951 vdd.n845 99.5127
R19325 vdd.n2951 vdd.n838 99.5127
R19326 vdd.n838 vdd.n804 99.5127
R19327 vdd.n3332 vdd.n804 99.5127
R19328 vdd.n2830 vdd.n2829 99.5127
R19329 vdd.n2834 vdd.n2833 99.5127
R19330 vdd.n2838 vdd.n2837 99.5127
R19331 vdd.n2842 vdd.n2841 99.5127
R19332 vdd.n2846 vdd.n2845 99.5127
R19333 vdd.n2850 vdd.n2849 99.5127
R19334 vdd.n2854 vdd.n2853 99.5127
R19335 vdd.n2858 vdd.n2857 99.5127
R19336 vdd.n2862 vdd.n2861 99.5127
R19337 vdd.n2866 vdd.n2865 99.5127
R19338 vdd.n2870 vdd.n2869 99.5127
R19339 vdd.n2874 vdd.n2873 99.5127
R19340 vdd.n2878 vdd.n2877 99.5127
R19341 vdd.n2882 vdd.n2881 99.5127
R19342 vdd.n2886 vdd.n2885 99.5127
R19343 vdd.n2890 vdd.n2889 99.5127
R19344 vdd.n2892 vdd.n2818 99.5127
R19345 vdd.n3096 vdd.n956 99.5127
R19346 vdd.n3096 vdd.n954 99.5127
R19347 vdd.n3100 vdd.n954 99.5127
R19348 vdd.n3100 vdd.n945 99.5127
R19349 vdd.n3108 vdd.n945 99.5127
R19350 vdd.n3108 vdd.n943 99.5127
R19351 vdd.n3112 vdd.n943 99.5127
R19352 vdd.n3112 vdd.n934 99.5127
R19353 vdd.n3120 vdd.n934 99.5127
R19354 vdd.n3120 vdd.n932 99.5127
R19355 vdd.n3124 vdd.n932 99.5127
R19356 vdd.n3124 vdd.n922 99.5127
R19357 vdd.n3132 vdd.n922 99.5127
R19358 vdd.n3132 vdd.n920 99.5127
R19359 vdd.n3136 vdd.n920 99.5127
R19360 vdd.n3136 vdd.n911 99.5127
R19361 vdd.n3144 vdd.n911 99.5127
R19362 vdd.n3144 vdd.n909 99.5127
R19363 vdd.n3149 vdd.n909 99.5127
R19364 vdd.n3149 vdd.n898 99.5127
R19365 vdd.n3157 vdd.n898 99.5127
R19366 vdd.n3157 vdd.n895 99.5127
R19367 vdd.n3161 vdd.n895 99.5127
R19368 vdd.n3161 vdd.n886 99.5127
R19369 vdd.n3169 vdd.n886 99.5127
R19370 vdd.n3169 vdd.n884 99.5127
R19371 vdd.n3173 vdd.n884 99.5127
R19372 vdd.n3173 vdd.n873 99.5127
R19373 vdd.n3181 vdd.n873 99.5127
R19374 vdd.n3181 vdd.n871 99.5127
R19375 vdd.n3185 vdd.n871 99.5127
R19376 vdd.n3185 vdd.n861 99.5127
R19377 vdd.n3193 vdd.n861 99.5127
R19378 vdd.n3193 vdd.n859 99.5127
R19379 vdd.n3197 vdd.n859 99.5127
R19380 vdd.n3197 vdd.n850 99.5127
R19381 vdd.n3205 vdd.n850 99.5127
R19382 vdd.n3205 vdd.n847 99.5127
R19383 vdd.n3254 vdd.n847 99.5127
R19384 vdd.n3254 vdd.n848 99.5127
R19385 vdd.n848 vdd.n839 99.5127
R19386 vdd.n3249 vdd.n839 99.5127
R19387 vdd.n3249 vdd.n807 99.5127
R19388 vdd.n2707 vdd.n2706 99.5127
R19389 vdd.n2703 vdd.n2702 99.5127
R19390 vdd.n2699 vdd.n2698 99.5127
R19391 vdd.n2695 vdd.n2694 99.5127
R19392 vdd.n2691 vdd.n2690 99.5127
R19393 vdd.n2687 vdd.n2686 99.5127
R19394 vdd.n2683 vdd.n2682 99.5127
R19395 vdd.n2679 vdd.n2678 99.5127
R19396 vdd.n2675 vdd.n2674 99.5127
R19397 vdd.n2671 vdd.n2670 99.5127
R19398 vdd.n2667 vdd.n2666 99.5127
R19399 vdd.n2663 vdd.n2662 99.5127
R19400 vdd.n2659 vdd.n2658 99.5127
R19401 vdd.n2655 vdd.n2654 99.5127
R19402 vdd.n2651 vdd.n2650 99.5127
R19403 vdd.n2647 vdd.n2646 99.5127
R19404 vdd.n2643 vdd.n980 99.5127
R19405 vdd.n1480 vdd.n1136 99.5127
R19406 vdd.n1477 vdd.n1136 99.5127
R19407 vdd.n1477 vdd.n1130 99.5127
R19408 vdd.n1474 vdd.n1130 99.5127
R19409 vdd.n1474 vdd.n1125 99.5127
R19410 vdd.n1471 vdd.n1125 99.5127
R19411 vdd.n1471 vdd.n1118 99.5127
R19412 vdd.n1468 vdd.n1118 99.5127
R19413 vdd.n1468 vdd.n1111 99.5127
R19414 vdd.n1465 vdd.n1111 99.5127
R19415 vdd.n1465 vdd.n1105 99.5127
R19416 vdd.n1462 vdd.n1105 99.5127
R19417 vdd.n1462 vdd.n1100 99.5127
R19418 vdd.n1459 vdd.n1100 99.5127
R19419 vdd.n1459 vdd.n1095 99.5127
R19420 vdd.n1456 vdd.n1095 99.5127
R19421 vdd.n1456 vdd.n1089 99.5127
R19422 vdd.n1453 vdd.n1089 99.5127
R19423 vdd.n1453 vdd.n1082 99.5127
R19424 vdd.n1450 vdd.n1082 99.5127
R19425 vdd.n1450 vdd.n1075 99.5127
R19426 vdd.n1447 vdd.n1075 99.5127
R19427 vdd.n1447 vdd.n1069 99.5127
R19428 vdd.n1444 vdd.n1069 99.5127
R19429 vdd.n1444 vdd.n1064 99.5127
R19430 vdd.n1441 vdd.n1064 99.5127
R19431 vdd.n1441 vdd.n1058 99.5127
R19432 vdd.n1438 vdd.n1058 99.5127
R19433 vdd.n1438 vdd.n1051 99.5127
R19434 vdd.n1409 vdd.n1051 99.5127
R19435 vdd.n1409 vdd.n1045 99.5127
R19436 vdd.n1412 vdd.n1045 99.5127
R19437 vdd.n1412 vdd.n1040 99.5127
R19438 vdd.n1424 vdd.n1040 99.5127
R19439 vdd.n1424 vdd.n1035 99.5127
R19440 vdd.n1420 vdd.n1035 99.5127
R19441 vdd.n1420 vdd.n1030 99.5127
R19442 vdd.n1417 vdd.n1030 99.5127
R19443 vdd.n1417 vdd.n1023 99.5127
R19444 vdd.n1023 vdd.n1014 99.5127
R19445 vdd.n2638 vdd.n1014 99.5127
R19446 vdd.n2639 vdd.n2638 99.5127
R19447 vdd.n2639 vdd.n1006 99.5127
R19448 vdd.n1284 vdd.n1283 99.5127
R19449 vdd.n1288 vdd.n1287 99.5127
R19450 vdd.n1292 vdd.n1291 99.5127
R19451 vdd.n1296 vdd.n1295 99.5127
R19452 vdd.n1300 vdd.n1299 99.5127
R19453 vdd.n1304 vdd.n1303 99.5127
R19454 vdd.n1308 vdd.n1307 99.5127
R19455 vdd.n1312 vdd.n1311 99.5127
R19456 vdd.n1513 vdd.n1314 99.5127
R19457 vdd.n1511 vdd.n1510 99.5127
R19458 vdd.n1507 vdd.n1506 99.5127
R19459 vdd.n1503 vdd.n1502 99.5127
R19460 vdd.n1499 vdd.n1498 99.5127
R19461 vdd.n1495 vdd.n1494 99.5127
R19462 vdd.n1491 vdd.n1490 99.5127
R19463 vdd.n1487 vdd.n1486 99.5127
R19464 vdd.n1483 vdd.n1175 99.5127
R19465 vdd.n2514 vdd.n1133 99.5127
R19466 vdd.n2514 vdd.n1131 99.5127
R19467 vdd.n2518 vdd.n1131 99.5127
R19468 vdd.n2518 vdd.n1122 99.5127
R19469 vdd.n2526 vdd.n1122 99.5127
R19470 vdd.n2526 vdd.n1120 99.5127
R19471 vdd.n2530 vdd.n1120 99.5127
R19472 vdd.n2530 vdd.n1109 99.5127
R19473 vdd.n2538 vdd.n1109 99.5127
R19474 vdd.n2538 vdd.n1107 99.5127
R19475 vdd.n2542 vdd.n1107 99.5127
R19476 vdd.n2542 vdd.n1098 99.5127
R19477 vdd.n2550 vdd.n1098 99.5127
R19478 vdd.n2550 vdd.n1096 99.5127
R19479 vdd.n2554 vdd.n1096 99.5127
R19480 vdd.n2554 vdd.n1086 99.5127
R19481 vdd.n2562 vdd.n1086 99.5127
R19482 vdd.n2562 vdd.n1084 99.5127
R19483 vdd.n2566 vdd.n1084 99.5127
R19484 vdd.n2566 vdd.n1073 99.5127
R19485 vdd.n2574 vdd.n1073 99.5127
R19486 vdd.n2574 vdd.n1070 99.5127
R19487 vdd.n2579 vdd.n1070 99.5127
R19488 vdd.n2579 vdd.n1061 99.5127
R19489 vdd.n2587 vdd.n1061 99.5127
R19490 vdd.n2587 vdd.n1059 99.5127
R19491 vdd.n2591 vdd.n1059 99.5127
R19492 vdd.n2591 vdd.n1049 99.5127
R19493 vdd.n2599 vdd.n1049 99.5127
R19494 vdd.n2599 vdd.n1047 99.5127
R19495 vdd.n2603 vdd.n1047 99.5127
R19496 vdd.n2603 vdd.n1038 99.5127
R19497 vdd.n2611 vdd.n1038 99.5127
R19498 vdd.n2611 vdd.n1036 99.5127
R19499 vdd.n2615 vdd.n1036 99.5127
R19500 vdd.n2615 vdd.n1027 99.5127
R19501 vdd.n2623 vdd.n1027 99.5127
R19502 vdd.n2623 vdd.n1024 99.5127
R19503 vdd.n2629 vdd.n1024 99.5127
R19504 vdd.n2629 vdd.n1025 99.5127
R19505 vdd.n1025 vdd.n1016 99.5127
R19506 vdd.n1016 vdd.n1007 99.5127
R19507 vdd.n2711 vdd.n1007 99.5127
R19508 vdd.n9 vdd.n7 98.9633
R19509 vdd.n2 vdd.n0 98.9633
R19510 vdd.n9 vdd.n8 98.6055
R19511 vdd.n11 vdd.n10 98.6055
R19512 vdd.n13 vdd.n12 98.6055
R19513 vdd.n6 vdd.n5 98.6055
R19514 vdd.n4 vdd.n3 98.6055
R19515 vdd.n2 vdd.n1 98.6055
R19516 vdd.t36 vdd.n303 85.8723
R19517 vdd.t152 vdd.n244 85.8723
R19518 vdd.t15 vdd.n201 85.8723
R19519 vdd.t141 vdd.n142 85.8723
R19520 vdd.t122 vdd.n100 85.8723
R19521 vdd.t82 vdd.n41 85.8723
R19522 vdd.t62 vdd.n2177 85.8723
R19523 vdd.t105 vdd.n2236 85.8723
R19524 vdd.t43 vdd.n2075 85.8723
R19525 vdd.t88 vdd.n2134 85.8723
R19526 vdd.t83 vdd.n1974 85.8723
R19527 vdd.t124 vdd.n2033 85.8723
R19528 vdd.n897 vdd.n896 78.546
R19529 vdd.n2577 vdd.n1071 78.546
R19530 vdd.n290 vdd.n289 75.1835
R19531 vdd.n288 vdd.n287 75.1835
R19532 vdd.n286 vdd.n285 75.1835
R19533 vdd.n284 vdd.n283 75.1835
R19534 vdd.n282 vdd.n281 75.1835
R19535 vdd.n280 vdd.n279 75.1835
R19536 vdd.n278 vdd.n277 75.1835
R19537 vdd.n276 vdd.n275 75.1835
R19538 vdd.n274 vdd.n273 75.1835
R19539 vdd.n188 vdd.n187 75.1835
R19540 vdd.n186 vdd.n185 75.1835
R19541 vdd.n184 vdd.n183 75.1835
R19542 vdd.n182 vdd.n181 75.1835
R19543 vdd.n180 vdd.n179 75.1835
R19544 vdd.n178 vdd.n177 75.1835
R19545 vdd.n176 vdd.n175 75.1835
R19546 vdd.n174 vdd.n173 75.1835
R19547 vdd.n172 vdd.n171 75.1835
R19548 vdd.n87 vdd.n86 75.1835
R19549 vdd.n85 vdd.n84 75.1835
R19550 vdd.n83 vdd.n82 75.1835
R19551 vdd.n81 vdd.n80 75.1835
R19552 vdd.n79 vdd.n78 75.1835
R19553 vdd.n77 vdd.n76 75.1835
R19554 vdd.n75 vdd.n74 75.1835
R19555 vdd.n73 vdd.n72 75.1835
R19556 vdd.n71 vdd.n70 75.1835
R19557 vdd.n2207 vdd.n2206 75.1835
R19558 vdd.n2209 vdd.n2208 75.1835
R19559 vdd.n2211 vdd.n2210 75.1835
R19560 vdd.n2213 vdd.n2212 75.1835
R19561 vdd.n2215 vdd.n2214 75.1835
R19562 vdd.n2217 vdd.n2216 75.1835
R19563 vdd.n2219 vdd.n2218 75.1835
R19564 vdd.n2221 vdd.n2220 75.1835
R19565 vdd.n2223 vdd.n2222 75.1835
R19566 vdd.n2105 vdd.n2104 75.1835
R19567 vdd.n2107 vdd.n2106 75.1835
R19568 vdd.n2109 vdd.n2108 75.1835
R19569 vdd.n2111 vdd.n2110 75.1835
R19570 vdd.n2113 vdd.n2112 75.1835
R19571 vdd.n2115 vdd.n2114 75.1835
R19572 vdd.n2117 vdd.n2116 75.1835
R19573 vdd.n2119 vdd.n2118 75.1835
R19574 vdd.n2121 vdd.n2120 75.1835
R19575 vdd.n2004 vdd.n2003 75.1835
R19576 vdd.n2006 vdd.n2005 75.1835
R19577 vdd.n2008 vdd.n2007 75.1835
R19578 vdd.n2010 vdd.n2009 75.1835
R19579 vdd.n2012 vdd.n2011 75.1835
R19580 vdd.n2014 vdd.n2013 75.1835
R19581 vdd.n2016 vdd.n2015 75.1835
R19582 vdd.n2018 vdd.n2017 75.1835
R19583 vdd.n2020 vdd.n2019 75.1835
R19584 vdd.n3088 vdd.n2801 72.8958
R19585 vdd.n3088 vdd.n2802 72.8958
R19586 vdd.n3088 vdd.n2803 72.8958
R19587 vdd.n3088 vdd.n2804 72.8958
R19588 vdd.n3088 vdd.n2805 72.8958
R19589 vdd.n3088 vdd.n2806 72.8958
R19590 vdd.n3088 vdd.n2807 72.8958
R19591 vdd.n3088 vdd.n2808 72.8958
R19592 vdd.n3088 vdd.n2809 72.8958
R19593 vdd.n3088 vdd.n2810 72.8958
R19594 vdd.n3088 vdd.n2811 72.8958
R19595 vdd.n3088 vdd.n2812 72.8958
R19596 vdd.n3088 vdd.n2813 72.8958
R19597 vdd.n3088 vdd.n2814 72.8958
R19598 vdd.n3088 vdd.n2815 72.8958
R19599 vdd.n3088 vdd.n2816 72.8958
R19600 vdd.n3088 vdd.n2817 72.8958
R19601 vdd.n803 vdd.n692 72.8958
R19602 vdd.n3338 vdd.n692 72.8958
R19603 vdd.n797 vdd.n692 72.8958
R19604 vdd.n3345 vdd.n692 72.8958
R19605 vdd.n794 vdd.n692 72.8958
R19606 vdd.n3352 vdd.n692 72.8958
R19607 vdd.n791 vdd.n692 72.8958
R19608 vdd.n3359 vdd.n692 72.8958
R19609 vdd.n3362 vdd.n692 72.8958
R19610 vdd.n3218 vdd.n692 72.8958
R19611 vdd.n3223 vdd.n692 72.8958
R19612 vdd.n3217 vdd.n692 72.8958
R19613 vdd.n3230 vdd.n692 72.8958
R19614 vdd.n3214 vdd.n692 72.8958
R19615 vdd.n3237 vdd.n692 72.8958
R19616 vdd.n3211 vdd.n692 72.8958
R19617 vdd.n3244 vdd.n692 72.8958
R19618 vdd.n2507 vdd.n2506 72.8958
R19619 vdd.n2506 vdd.n1142 72.8958
R19620 vdd.n2506 vdd.n1143 72.8958
R19621 vdd.n2506 vdd.n1144 72.8958
R19622 vdd.n2506 vdd.n1145 72.8958
R19623 vdd.n2506 vdd.n1146 72.8958
R19624 vdd.n2506 vdd.n1147 72.8958
R19625 vdd.n2506 vdd.n1148 72.8958
R19626 vdd.n2506 vdd.n1149 72.8958
R19627 vdd.n2506 vdd.n1150 72.8958
R19628 vdd.n2506 vdd.n1151 72.8958
R19629 vdd.n2506 vdd.n1152 72.8958
R19630 vdd.n2506 vdd.n1153 72.8958
R19631 vdd.n2506 vdd.n1154 72.8958
R19632 vdd.n2506 vdd.n1155 72.8958
R19633 vdd.n2506 vdd.n1156 72.8958
R19634 vdd.n2506 vdd.n1157 72.8958
R19635 vdd.n2784 vdd.n981 72.8958
R19636 vdd.n2784 vdd.n982 72.8958
R19637 vdd.n2784 vdd.n983 72.8958
R19638 vdd.n2784 vdd.n984 72.8958
R19639 vdd.n2784 vdd.n985 72.8958
R19640 vdd.n2784 vdd.n986 72.8958
R19641 vdd.n2784 vdd.n987 72.8958
R19642 vdd.n2784 vdd.n988 72.8958
R19643 vdd.n2784 vdd.n989 72.8958
R19644 vdd.n2784 vdd.n990 72.8958
R19645 vdd.n2784 vdd.n991 72.8958
R19646 vdd.n2784 vdd.n992 72.8958
R19647 vdd.n2784 vdd.n993 72.8958
R19648 vdd.n2784 vdd.n994 72.8958
R19649 vdd.n2784 vdd.n995 72.8958
R19650 vdd.n2784 vdd.n996 72.8958
R19651 vdd.n2784 vdd.n997 72.8958
R19652 vdd.n3089 vdd.n3088 72.8958
R19653 vdd.n3088 vdd.n2785 72.8958
R19654 vdd.n3088 vdd.n2786 72.8958
R19655 vdd.n3088 vdd.n2787 72.8958
R19656 vdd.n3088 vdd.n2788 72.8958
R19657 vdd.n3088 vdd.n2789 72.8958
R19658 vdd.n3088 vdd.n2790 72.8958
R19659 vdd.n3088 vdd.n2791 72.8958
R19660 vdd.n3088 vdd.n2792 72.8958
R19661 vdd.n3088 vdd.n2793 72.8958
R19662 vdd.n3088 vdd.n2794 72.8958
R19663 vdd.n3088 vdd.n2795 72.8958
R19664 vdd.n3088 vdd.n2796 72.8958
R19665 vdd.n3088 vdd.n2797 72.8958
R19666 vdd.n3088 vdd.n2798 72.8958
R19667 vdd.n3088 vdd.n2799 72.8958
R19668 vdd.n3088 vdd.n2800 72.8958
R19669 vdd.n3268 vdd.n692 72.8958
R19670 vdd.n835 vdd.n692 72.8958
R19671 vdd.n3276 vdd.n692 72.8958
R19672 vdd.n830 vdd.n692 72.8958
R19673 vdd.n3283 vdd.n692 72.8958
R19674 vdd.n827 vdd.n692 72.8958
R19675 vdd.n3290 vdd.n692 72.8958
R19676 vdd.n824 vdd.n692 72.8958
R19677 vdd.n3297 vdd.n692 72.8958
R19678 vdd.n3301 vdd.n692 72.8958
R19679 vdd.n821 vdd.n692 72.8958
R19680 vdd.n3308 vdd.n692 72.8958
R19681 vdd.n818 vdd.n692 72.8958
R19682 vdd.n3315 vdd.n692 72.8958
R19683 vdd.n815 vdd.n692 72.8958
R19684 vdd.n3322 vdd.n692 72.8958
R19685 vdd.n3325 vdd.n692 72.8958
R19686 vdd.n2784 vdd.n979 72.8958
R19687 vdd.n2784 vdd.n978 72.8958
R19688 vdd.n2784 vdd.n977 72.8958
R19689 vdd.n2784 vdd.n976 72.8958
R19690 vdd.n2784 vdd.n975 72.8958
R19691 vdd.n2784 vdd.n974 72.8958
R19692 vdd.n2784 vdd.n973 72.8958
R19693 vdd.n2784 vdd.n972 72.8958
R19694 vdd.n2784 vdd.n971 72.8958
R19695 vdd.n2784 vdd.n970 72.8958
R19696 vdd.n2784 vdd.n969 72.8958
R19697 vdd.n2784 vdd.n968 72.8958
R19698 vdd.n2784 vdd.n967 72.8958
R19699 vdd.n2784 vdd.n966 72.8958
R19700 vdd.n2784 vdd.n965 72.8958
R19701 vdd.n2784 vdd.n964 72.8958
R19702 vdd.n2784 vdd.n963 72.8958
R19703 vdd.n2506 vdd.n1158 72.8958
R19704 vdd.n2506 vdd.n1159 72.8958
R19705 vdd.n2506 vdd.n1160 72.8958
R19706 vdd.n2506 vdd.n1161 72.8958
R19707 vdd.n2506 vdd.n1162 72.8958
R19708 vdd.n2506 vdd.n1163 72.8958
R19709 vdd.n2506 vdd.n1164 72.8958
R19710 vdd.n2506 vdd.n1165 72.8958
R19711 vdd.n2506 vdd.n1166 72.8958
R19712 vdd.n2506 vdd.n1167 72.8958
R19713 vdd.n2506 vdd.n1168 72.8958
R19714 vdd.n2506 vdd.n1169 72.8958
R19715 vdd.n2506 vdd.n1170 72.8958
R19716 vdd.n2506 vdd.n1171 72.8958
R19717 vdd.n2506 vdd.n1172 72.8958
R19718 vdd.n2506 vdd.n1173 72.8958
R19719 vdd.n2506 vdd.n1174 72.8958
R19720 vdd.n1874 vdd.n1873 66.2847
R19721 vdd.n1873 vdd.n1649 66.2847
R19722 vdd.n1873 vdd.n1650 66.2847
R19723 vdd.n1873 vdd.n1651 66.2847
R19724 vdd.n1873 vdd.n1652 66.2847
R19725 vdd.n1873 vdd.n1653 66.2847
R19726 vdd.n1873 vdd.n1654 66.2847
R19727 vdd.n1873 vdd.n1655 66.2847
R19728 vdd.n1873 vdd.n1656 66.2847
R19729 vdd.n1873 vdd.n1657 66.2847
R19730 vdd.n1873 vdd.n1658 66.2847
R19731 vdd.n1873 vdd.n1659 66.2847
R19732 vdd.n1873 vdd.n1660 66.2847
R19733 vdd.n1873 vdd.n1661 66.2847
R19734 vdd.n1873 vdd.n1662 66.2847
R19735 vdd.n1873 vdd.n1663 66.2847
R19736 vdd.n1873 vdd.n1664 66.2847
R19737 vdd.n1873 vdd.n1665 66.2847
R19738 vdd.n1873 vdd.n1666 66.2847
R19739 vdd.n1873 vdd.n1667 66.2847
R19740 vdd.n1873 vdd.n1668 66.2847
R19741 vdd.n1873 vdd.n1669 66.2847
R19742 vdd.n1873 vdd.n1670 66.2847
R19743 vdd.n1873 vdd.n1671 66.2847
R19744 vdd.n1873 vdd.n1672 66.2847
R19745 vdd.n1873 vdd.n1673 66.2847
R19746 vdd.n1873 vdd.n1674 66.2847
R19747 vdd.n1873 vdd.n1675 66.2847
R19748 vdd.n1873 vdd.n1676 66.2847
R19749 vdd.n1873 vdd.n1677 66.2847
R19750 vdd.n1873 vdd.n1678 66.2847
R19751 vdd.n1526 vdd.n1141 66.2847
R19752 vdd.n1523 vdd.n1141 66.2847
R19753 vdd.n1519 vdd.n1141 66.2847
R19754 vdd.n2372 vdd.n1141 66.2847
R19755 vdd.n1275 vdd.n1141 66.2847
R19756 vdd.n2379 vdd.n1141 66.2847
R19757 vdd.n1268 vdd.n1141 66.2847
R19758 vdd.n2386 vdd.n1141 66.2847
R19759 vdd.n1261 vdd.n1141 66.2847
R19760 vdd.n2393 vdd.n1141 66.2847
R19761 vdd.n1255 vdd.n1141 66.2847
R19762 vdd.n1250 vdd.n1141 66.2847
R19763 vdd.n2404 vdd.n1141 66.2847
R19764 vdd.n1242 vdd.n1141 66.2847
R19765 vdd.n2411 vdd.n1141 66.2847
R19766 vdd.n1235 vdd.n1141 66.2847
R19767 vdd.n2418 vdd.n1141 66.2847
R19768 vdd.n1228 vdd.n1141 66.2847
R19769 vdd.n2425 vdd.n1141 66.2847
R19770 vdd.n1221 vdd.n1141 66.2847
R19771 vdd.n2432 vdd.n1141 66.2847
R19772 vdd.n1215 vdd.n1141 66.2847
R19773 vdd.n1210 vdd.n1141 66.2847
R19774 vdd.n2443 vdd.n1141 66.2847
R19775 vdd.n1202 vdd.n1141 66.2847
R19776 vdd.n2450 vdd.n1141 66.2847
R19777 vdd.n1195 vdd.n1141 66.2847
R19778 vdd.n2457 vdd.n1141 66.2847
R19779 vdd.n1188 vdd.n1141 66.2847
R19780 vdd.n2464 vdd.n1141 66.2847
R19781 vdd.n2469 vdd.n1141 66.2847
R19782 vdd.n1184 vdd.n1141 66.2847
R19783 vdd.n3495 vdd.n3494 66.2847
R19784 vdd.n3495 vdd.n693 66.2847
R19785 vdd.n3495 vdd.n694 66.2847
R19786 vdd.n3495 vdd.n695 66.2847
R19787 vdd.n3495 vdd.n696 66.2847
R19788 vdd.n3495 vdd.n697 66.2847
R19789 vdd.n3495 vdd.n698 66.2847
R19790 vdd.n3495 vdd.n699 66.2847
R19791 vdd.n3495 vdd.n700 66.2847
R19792 vdd.n3495 vdd.n701 66.2847
R19793 vdd.n3495 vdd.n702 66.2847
R19794 vdd.n3495 vdd.n703 66.2847
R19795 vdd.n3495 vdd.n704 66.2847
R19796 vdd.n3495 vdd.n705 66.2847
R19797 vdd.n3495 vdd.n706 66.2847
R19798 vdd.n3495 vdd.n707 66.2847
R19799 vdd.n3495 vdd.n708 66.2847
R19800 vdd.n3495 vdd.n709 66.2847
R19801 vdd.n3495 vdd.n710 66.2847
R19802 vdd.n3495 vdd.n711 66.2847
R19803 vdd.n3495 vdd.n712 66.2847
R19804 vdd.n3495 vdd.n713 66.2847
R19805 vdd.n3495 vdd.n714 66.2847
R19806 vdd.n3495 vdd.n715 66.2847
R19807 vdd.n3495 vdd.n716 66.2847
R19808 vdd.n3495 vdd.n717 66.2847
R19809 vdd.n3495 vdd.n718 66.2847
R19810 vdd.n3495 vdd.n719 66.2847
R19811 vdd.n3495 vdd.n720 66.2847
R19812 vdd.n3495 vdd.n721 66.2847
R19813 vdd.n3495 vdd.n722 66.2847
R19814 vdd.n3626 vdd.n3625 66.2847
R19815 vdd.n3626 vdd.n424 66.2847
R19816 vdd.n3626 vdd.n423 66.2847
R19817 vdd.n3626 vdd.n422 66.2847
R19818 vdd.n3626 vdd.n421 66.2847
R19819 vdd.n3626 vdd.n420 66.2847
R19820 vdd.n3626 vdd.n419 66.2847
R19821 vdd.n3626 vdd.n418 66.2847
R19822 vdd.n3626 vdd.n417 66.2847
R19823 vdd.n3626 vdd.n416 66.2847
R19824 vdd.n3626 vdd.n415 66.2847
R19825 vdd.n3626 vdd.n414 66.2847
R19826 vdd.n3626 vdd.n413 66.2847
R19827 vdd.n3626 vdd.n412 66.2847
R19828 vdd.n3626 vdd.n411 66.2847
R19829 vdd.n3626 vdd.n410 66.2847
R19830 vdd.n3626 vdd.n409 66.2847
R19831 vdd.n3626 vdd.n408 66.2847
R19832 vdd.n3626 vdd.n407 66.2847
R19833 vdd.n3626 vdd.n406 66.2847
R19834 vdd.n3626 vdd.n405 66.2847
R19835 vdd.n3626 vdd.n404 66.2847
R19836 vdd.n3626 vdd.n403 66.2847
R19837 vdd.n3626 vdd.n402 66.2847
R19838 vdd.n3626 vdd.n401 66.2847
R19839 vdd.n3626 vdd.n400 66.2847
R19840 vdd.n3626 vdd.n399 66.2847
R19841 vdd.n3626 vdd.n398 66.2847
R19842 vdd.n3626 vdd.n397 66.2847
R19843 vdd.n3626 vdd.n396 66.2847
R19844 vdd.n3626 vdd.n395 66.2847
R19845 vdd.n3626 vdd.n394 66.2847
R19846 vdd.n467 vdd.n394 52.4337
R19847 vdd.n473 vdd.n395 52.4337
R19848 vdd.n477 vdd.n396 52.4337
R19849 vdd.n483 vdd.n397 52.4337
R19850 vdd.n487 vdd.n398 52.4337
R19851 vdd.n493 vdd.n399 52.4337
R19852 vdd.n497 vdd.n400 52.4337
R19853 vdd.n503 vdd.n401 52.4337
R19854 vdd.n507 vdd.n402 52.4337
R19855 vdd.n513 vdd.n403 52.4337
R19856 vdd.n517 vdd.n404 52.4337
R19857 vdd.n523 vdd.n405 52.4337
R19858 vdd.n527 vdd.n406 52.4337
R19859 vdd.n533 vdd.n407 52.4337
R19860 vdd.n537 vdd.n408 52.4337
R19861 vdd.n543 vdd.n409 52.4337
R19862 vdd.n547 vdd.n410 52.4337
R19863 vdd.n553 vdd.n411 52.4337
R19864 vdd.n557 vdd.n412 52.4337
R19865 vdd.n563 vdd.n413 52.4337
R19866 vdd.n567 vdd.n414 52.4337
R19867 vdd.n573 vdd.n415 52.4337
R19868 vdd.n577 vdd.n416 52.4337
R19869 vdd.n583 vdd.n417 52.4337
R19870 vdd.n587 vdd.n418 52.4337
R19871 vdd.n593 vdd.n419 52.4337
R19872 vdd.n597 vdd.n420 52.4337
R19873 vdd.n603 vdd.n421 52.4337
R19874 vdd.n607 vdd.n422 52.4337
R19875 vdd.n613 vdd.n423 52.4337
R19876 vdd.n616 vdd.n424 52.4337
R19877 vdd.n3625 vdd.n3624 52.4337
R19878 vdd.n3494 vdd.n3493 52.4337
R19879 vdd.n728 vdd.n693 52.4337
R19880 vdd.n734 vdd.n694 52.4337
R19881 vdd.n3483 vdd.n695 52.4337
R19882 vdd.n3479 vdd.n696 52.4337
R19883 vdd.n3475 vdd.n697 52.4337
R19884 vdd.n3471 vdd.n698 52.4337
R19885 vdd.n3467 vdd.n699 52.4337
R19886 vdd.n3463 vdd.n700 52.4337
R19887 vdd.n3459 vdd.n701 52.4337
R19888 vdd.n3451 vdd.n702 52.4337
R19889 vdd.n3447 vdd.n703 52.4337
R19890 vdd.n3443 vdd.n704 52.4337
R19891 vdd.n3439 vdd.n705 52.4337
R19892 vdd.n3435 vdd.n706 52.4337
R19893 vdd.n3431 vdd.n707 52.4337
R19894 vdd.n3427 vdd.n708 52.4337
R19895 vdd.n3423 vdd.n709 52.4337
R19896 vdd.n3419 vdd.n710 52.4337
R19897 vdd.n3415 vdd.n711 52.4337
R19898 vdd.n3411 vdd.n712 52.4337
R19899 vdd.n3405 vdd.n713 52.4337
R19900 vdd.n3401 vdd.n714 52.4337
R19901 vdd.n3397 vdd.n715 52.4337
R19902 vdd.n3393 vdd.n716 52.4337
R19903 vdd.n3389 vdd.n717 52.4337
R19904 vdd.n3385 vdd.n718 52.4337
R19905 vdd.n3381 vdd.n719 52.4337
R19906 vdd.n3377 vdd.n720 52.4337
R19907 vdd.n3373 vdd.n721 52.4337
R19908 vdd.n3369 vdd.n722 52.4337
R19909 vdd.n2471 vdd.n1184 52.4337
R19910 vdd.n2469 vdd.n2468 52.4337
R19911 vdd.n2464 vdd.n2463 52.4337
R19912 vdd.n2459 vdd.n1188 52.4337
R19913 vdd.n2457 vdd.n2456 52.4337
R19914 vdd.n2452 vdd.n1195 52.4337
R19915 vdd.n2450 vdd.n2449 52.4337
R19916 vdd.n2445 vdd.n1202 52.4337
R19917 vdd.n2443 vdd.n2442 52.4337
R19918 vdd.n1211 vdd.n1210 52.4337
R19919 vdd.n2434 vdd.n1215 52.4337
R19920 vdd.n2432 vdd.n2431 52.4337
R19921 vdd.n2427 vdd.n1221 52.4337
R19922 vdd.n2425 vdd.n2424 52.4337
R19923 vdd.n2420 vdd.n1228 52.4337
R19924 vdd.n2418 vdd.n2417 52.4337
R19925 vdd.n2413 vdd.n1235 52.4337
R19926 vdd.n2411 vdd.n2410 52.4337
R19927 vdd.n2406 vdd.n1242 52.4337
R19928 vdd.n2404 vdd.n2403 52.4337
R19929 vdd.n1251 vdd.n1250 52.4337
R19930 vdd.n2395 vdd.n1255 52.4337
R19931 vdd.n2393 vdd.n2392 52.4337
R19932 vdd.n2388 vdd.n1261 52.4337
R19933 vdd.n2386 vdd.n2385 52.4337
R19934 vdd.n2381 vdd.n1268 52.4337
R19935 vdd.n2379 vdd.n2378 52.4337
R19936 vdd.n2374 vdd.n1275 52.4337
R19937 vdd.n2372 vdd.n2371 52.4337
R19938 vdd.n1520 vdd.n1519 52.4337
R19939 vdd.n1524 vdd.n1523 52.4337
R19940 vdd.n2360 vdd.n1526 52.4337
R19941 vdd.n1875 vdd.n1874 52.4337
R19942 vdd.n1681 vdd.n1649 52.4337
R19943 vdd.n1685 vdd.n1650 52.4337
R19944 vdd.n1687 vdd.n1651 52.4337
R19945 vdd.n1691 vdd.n1652 52.4337
R19946 vdd.n1693 vdd.n1653 52.4337
R19947 vdd.n1697 vdd.n1654 52.4337
R19948 vdd.n1699 vdd.n1655 52.4337
R19949 vdd.n1703 vdd.n1656 52.4337
R19950 vdd.n1705 vdd.n1657 52.4337
R19951 vdd.n1711 vdd.n1658 52.4337
R19952 vdd.n1713 vdd.n1659 52.4337
R19953 vdd.n1717 vdd.n1660 52.4337
R19954 vdd.n1719 vdd.n1661 52.4337
R19955 vdd.n1723 vdd.n1662 52.4337
R19956 vdd.n1725 vdd.n1663 52.4337
R19957 vdd.n1729 vdd.n1664 52.4337
R19958 vdd.n1731 vdd.n1665 52.4337
R19959 vdd.n1735 vdd.n1666 52.4337
R19960 vdd.n1737 vdd.n1667 52.4337
R19961 vdd.n1809 vdd.n1668 52.4337
R19962 vdd.n1742 vdd.n1669 52.4337
R19963 vdd.n1746 vdd.n1670 52.4337
R19964 vdd.n1748 vdd.n1671 52.4337
R19965 vdd.n1752 vdd.n1672 52.4337
R19966 vdd.n1754 vdd.n1673 52.4337
R19967 vdd.n1758 vdd.n1674 52.4337
R19968 vdd.n1760 vdd.n1675 52.4337
R19969 vdd.n1764 vdd.n1676 52.4337
R19970 vdd.n1766 vdd.n1677 52.4337
R19971 vdd.n1770 vdd.n1678 52.4337
R19972 vdd.n1874 vdd.n1648 52.4337
R19973 vdd.n1684 vdd.n1649 52.4337
R19974 vdd.n1686 vdd.n1650 52.4337
R19975 vdd.n1690 vdd.n1651 52.4337
R19976 vdd.n1692 vdd.n1652 52.4337
R19977 vdd.n1696 vdd.n1653 52.4337
R19978 vdd.n1698 vdd.n1654 52.4337
R19979 vdd.n1702 vdd.n1655 52.4337
R19980 vdd.n1704 vdd.n1656 52.4337
R19981 vdd.n1710 vdd.n1657 52.4337
R19982 vdd.n1712 vdd.n1658 52.4337
R19983 vdd.n1716 vdd.n1659 52.4337
R19984 vdd.n1718 vdd.n1660 52.4337
R19985 vdd.n1722 vdd.n1661 52.4337
R19986 vdd.n1724 vdd.n1662 52.4337
R19987 vdd.n1728 vdd.n1663 52.4337
R19988 vdd.n1730 vdd.n1664 52.4337
R19989 vdd.n1734 vdd.n1665 52.4337
R19990 vdd.n1736 vdd.n1666 52.4337
R19991 vdd.n1740 vdd.n1667 52.4337
R19992 vdd.n1741 vdd.n1668 52.4337
R19993 vdd.n1745 vdd.n1669 52.4337
R19994 vdd.n1747 vdd.n1670 52.4337
R19995 vdd.n1751 vdd.n1671 52.4337
R19996 vdd.n1753 vdd.n1672 52.4337
R19997 vdd.n1757 vdd.n1673 52.4337
R19998 vdd.n1759 vdd.n1674 52.4337
R19999 vdd.n1763 vdd.n1675 52.4337
R20000 vdd.n1765 vdd.n1676 52.4337
R20001 vdd.n1769 vdd.n1677 52.4337
R20002 vdd.n1771 vdd.n1678 52.4337
R20003 vdd.n1526 vdd.n1525 52.4337
R20004 vdd.n1523 vdd.n1522 52.4337
R20005 vdd.n1519 vdd.n1276 52.4337
R20006 vdd.n2373 vdd.n2372 52.4337
R20007 vdd.n1275 vdd.n1269 52.4337
R20008 vdd.n2380 vdd.n2379 52.4337
R20009 vdd.n1268 vdd.n1262 52.4337
R20010 vdd.n2387 vdd.n2386 52.4337
R20011 vdd.n1261 vdd.n1256 52.4337
R20012 vdd.n2394 vdd.n2393 52.4337
R20013 vdd.n1255 vdd.n1254 52.4337
R20014 vdd.n1250 vdd.n1243 52.4337
R20015 vdd.n2405 vdd.n2404 52.4337
R20016 vdd.n1242 vdd.n1236 52.4337
R20017 vdd.n2412 vdd.n2411 52.4337
R20018 vdd.n1235 vdd.n1229 52.4337
R20019 vdd.n2419 vdd.n2418 52.4337
R20020 vdd.n1228 vdd.n1222 52.4337
R20021 vdd.n2426 vdd.n2425 52.4337
R20022 vdd.n1221 vdd.n1216 52.4337
R20023 vdd.n2433 vdd.n2432 52.4337
R20024 vdd.n1215 vdd.n1214 52.4337
R20025 vdd.n1210 vdd.n1203 52.4337
R20026 vdd.n2444 vdd.n2443 52.4337
R20027 vdd.n1202 vdd.n1196 52.4337
R20028 vdd.n2451 vdd.n2450 52.4337
R20029 vdd.n1195 vdd.n1189 52.4337
R20030 vdd.n2458 vdd.n2457 52.4337
R20031 vdd.n1188 vdd.n1185 52.4337
R20032 vdd.n2465 vdd.n2464 52.4337
R20033 vdd.n2470 vdd.n2469 52.4337
R20034 vdd.n1530 vdd.n1184 52.4337
R20035 vdd.n3494 vdd.n725 52.4337
R20036 vdd.n733 vdd.n693 52.4337
R20037 vdd.n3484 vdd.n694 52.4337
R20038 vdd.n3480 vdd.n695 52.4337
R20039 vdd.n3476 vdd.n696 52.4337
R20040 vdd.n3472 vdd.n697 52.4337
R20041 vdd.n3468 vdd.n698 52.4337
R20042 vdd.n3464 vdd.n699 52.4337
R20043 vdd.n3460 vdd.n700 52.4337
R20044 vdd.n3450 vdd.n701 52.4337
R20045 vdd.n3448 vdd.n702 52.4337
R20046 vdd.n3444 vdd.n703 52.4337
R20047 vdd.n3440 vdd.n704 52.4337
R20048 vdd.n3436 vdd.n705 52.4337
R20049 vdd.n3432 vdd.n706 52.4337
R20050 vdd.n3428 vdd.n707 52.4337
R20051 vdd.n3424 vdd.n708 52.4337
R20052 vdd.n3420 vdd.n709 52.4337
R20053 vdd.n3416 vdd.n710 52.4337
R20054 vdd.n3412 vdd.n711 52.4337
R20055 vdd.n3404 vdd.n712 52.4337
R20056 vdd.n3402 vdd.n713 52.4337
R20057 vdd.n3398 vdd.n714 52.4337
R20058 vdd.n3394 vdd.n715 52.4337
R20059 vdd.n3390 vdd.n716 52.4337
R20060 vdd.n3386 vdd.n717 52.4337
R20061 vdd.n3382 vdd.n718 52.4337
R20062 vdd.n3378 vdd.n719 52.4337
R20063 vdd.n3374 vdd.n720 52.4337
R20064 vdd.n3370 vdd.n721 52.4337
R20065 vdd.n722 vdd.n691 52.4337
R20066 vdd.n3625 vdd.n425 52.4337
R20067 vdd.n614 vdd.n424 52.4337
R20068 vdd.n608 vdd.n423 52.4337
R20069 vdd.n604 vdd.n422 52.4337
R20070 vdd.n598 vdd.n421 52.4337
R20071 vdd.n594 vdd.n420 52.4337
R20072 vdd.n588 vdd.n419 52.4337
R20073 vdd.n584 vdd.n418 52.4337
R20074 vdd.n578 vdd.n417 52.4337
R20075 vdd.n574 vdd.n416 52.4337
R20076 vdd.n568 vdd.n415 52.4337
R20077 vdd.n564 vdd.n414 52.4337
R20078 vdd.n558 vdd.n413 52.4337
R20079 vdd.n554 vdd.n412 52.4337
R20080 vdd.n548 vdd.n411 52.4337
R20081 vdd.n544 vdd.n410 52.4337
R20082 vdd.n538 vdd.n409 52.4337
R20083 vdd.n534 vdd.n408 52.4337
R20084 vdd.n528 vdd.n407 52.4337
R20085 vdd.n524 vdd.n406 52.4337
R20086 vdd.n518 vdd.n405 52.4337
R20087 vdd.n514 vdd.n404 52.4337
R20088 vdd.n508 vdd.n403 52.4337
R20089 vdd.n504 vdd.n402 52.4337
R20090 vdd.n498 vdd.n401 52.4337
R20091 vdd.n494 vdd.n400 52.4337
R20092 vdd.n488 vdd.n399 52.4337
R20093 vdd.n484 vdd.n398 52.4337
R20094 vdd.n478 vdd.n397 52.4337
R20095 vdd.n474 vdd.n396 52.4337
R20096 vdd.n468 vdd.n395 52.4337
R20097 vdd.n394 vdd.n392 52.4337
R20098 vdd.t251 vdd.t264 51.4683
R20099 vdd.n274 vdd.n272 42.0461
R20100 vdd.n172 vdd.n170 42.0461
R20101 vdd.n71 vdd.n69 42.0461
R20102 vdd.n2207 vdd.n2205 42.0461
R20103 vdd.n2105 vdd.n2103 42.0461
R20104 vdd.n2004 vdd.n2002 42.0461
R20105 vdd.n332 vdd.n331 41.6884
R20106 vdd.n230 vdd.n229 41.6884
R20107 vdd.n129 vdd.n128 41.6884
R20108 vdd.n2265 vdd.n2264 41.6884
R20109 vdd.n2163 vdd.n2162 41.6884
R20110 vdd.n2062 vdd.n2061 41.6884
R20111 vdd.n1774 vdd.n1773 41.1157
R20112 vdd.n1812 vdd.n1811 41.1157
R20113 vdd.n1708 vdd.n1707 41.1157
R20114 vdd.n428 vdd.n427 41.1157
R20115 vdd.n566 vdd.n441 41.1157
R20116 vdd.n454 vdd.n453 41.1157
R20117 vdd.n3325 vdd.n3324 39.2114
R20118 vdd.n3322 vdd.n3321 39.2114
R20119 vdd.n3317 vdd.n815 39.2114
R20120 vdd.n3315 vdd.n3314 39.2114
R20121 vdd.n3310 vdd.n818 39.2114
R20122 vdd.n3308 vdd.n3307 39.2114
R20123 vdd.n3303 vdd.n821 39.2114
R20124 vdd.n3301 vdd.n3300 39.2114
R20125 vdd.n3297 vdd.n3296 39.2114
R20126 vdd.n3292 vdd.n824 39.2114
R20127 vdd.n3290 vdd.n3289 39.2114
R20128 vdd.n3285 vdd.n827 39.2114
R20129 vdd.n3283 vdd.n3282 39.2114
R20130 vdd.n3278 vdd.n830 39.2114
R20131 vdd.n3276 vdd.n3275 39.2114
R20132 vdd.n3270 vdd.n835 39.2114
R20133 vdd.n3268 vdd.n3267 39.2114
R20134 vdd.n3090 vdd.n3089 39.2114
R20135 vdd.n2819 vdd.n2785 39.2114
R20136 vdd.n3082 vdd.n2786 39.2114
R20137 vdd.n3078 vdd.n2787 39.2114
R20138 vdd.n3074 vdd.n2788 39.2114
R20139 vdd.n3070 vdd.n2789 39.2114
R20140 vdd.n3066 vdd.n2790 39.2114
R20141 vdd.n3062 vdd.n2791 39.2114
R20142 vdd.n3058 vdd.n2792 39.2114
R20143 vdd.n3054 vdd.n2793 39.2114
R20144 vdd.n3050 vdd.n2794 39.2114
R20145 vdd.n3046 vdd.n2795 39.2114
R20146 vdd.n3042 vdd.n2796 39.2114
R20147 vdd.n3038 vdd.n2797 39.2114
R20148 vdd.n3034 vdd.n2798 39.2114
R20149 vdd.n3030 vdd.n2799 39.2114
R20150 vdd.n3025 vdd.n2800 39.2114
R20151 vdd.n2779 vdd.n997 39.2114
R20152 vdd.n2775 vdd.n996 39.2114
R20153 vdd.n2771 vdd.n995 39.2114
R20154 vdd.n2767 vdd.n994 39.2114
R20155 vdd.n2763 vdd.n993 39.2114
R20156 vdd.n2759 vdd.n992 39.2114
R20157 vdd.n2755 vdd.n991 39.2114
R20158 vdd.n2751 vdd.n990 39.2114
R20159 vdd.n2747 vdd.n989 39.2114
R20160 vdd.n2743 vdd.n988 39.2114
R20161 vdd.n2739 vdd.n987 39.2114
R20162 vdd.n2735 vdd.n986 39.2114
R20163 vdd.n2731 vdd.n985 39.2114
R20164 vdd.n2727 vdd.n984 39.2114
R20165 vdd.n2723 vdd.n983 39.2114
R20166 vdd.n2718 vdd.n982 39.2114
R20167 vdd.n2714 vdd.n981 39.2114
R20168 vdd.n2508 vdd.n2507 39.2114
R20169 vdd.n1176 vdd.n1142 39.2114
R20170 vdd.n2500 vdd.n1143 39.2114
R20171 vdd.n2496 vdd.n1144 39.2114
R20172 vdd.n2492 vdd.n1145 39.2114
R20173 vdd.n2488 vdd.n1146 39.2114
R20174 vdd.n2484 vdd.n1147 39.2114
R20175 vdd.n2480 vdd.n1148 39.2114
R20176 vdd.n2476 vdd.n1149 39.2114
R20177 vdd.n1322 vdd.n1150 39.2114
R20178 vdd.n1326 vdd.n1151 39.2114
R20179 vdd.n1330 vdd.n1152 39.2114
R20180 vdd.n1334 vdd.n1153 39.2114
R20181 vdd.n1338 vdd.n1154 39.2114
R20182 vdd.n1342 vdd.n1155 39.2114
R20183 vdd.n1346 vdd.n1156 39.2114
R20184 vdd.n1351 vdd.n1157 39.2114
R20185 vdd.n3244 vdd.n3243 39.2114
R20186 vdd.n3239 vdd.n3211 39.2114
R20187 vdd.n3237 vdd.n3236 39.2114
R20188 vdd.n3232 vdd.n3214 39.2114
R20189 vdd.n3230 vdd.n3229 39.2114
R20190 vdd.n3225 vdd.n3217 39.2114
R20191 vdd.n3223 vdd.n3222 39.2114
R20192 vdd.n3218 vdd.n787 39.2114
R20193 vdd.n3362 vdd.n3361 39.2114
R20194 vdd.n3359 vdd.n3358 39.2114
R20195 vdd.n3354 vdd.n791 39.2114
R20196 vdd.n3352 vdd.n3351 39.2114
R20197 vdd.n3347 vdd.n794 39.2114
R20198 vdd.n3345 vdd.n3344 39.2114
R20199 vdd.n3340 vdd.n797 39.2114
R20200 vdd.n3338 vdd.n3337 39.2114
R20201 vdd.n3333 vdd.n803 39.2114
R20202 vdd.n2826 vdd.n2801 39.2114
R20203 vdd.n2830 vdd.n2802 39.2114
R20204 vdd.n2834 vdd.n2803 39.2114
R20205 vdd.n2838 vdd.n2804 39.2114
R20206 vdd.n2842 vdd.n2805 39.2114
R20207 vdd.n2846 vdd.n2806 39.2114
R20208 vdd.n2850 vdd.n2807 39.2114
R20209 vdd.n2854 vdd.n2808 39.2114
R20210 vdd.n2858 vdd.n2809 39.2114
R20211 vdd.n2862 vdd.n2810 39.2114
R20212 vdd.n2866 vdd.n2811 39.2114
R20213 vdd.n2870 vdd.n2812 39.2114
R20214 vdd.n2874 vdd.n2813 39.2114
R20215 vdd.n2878 vdd.n2814 39.2114
R20216 vdd.n2882 vdd.n2815 39.2114
R20217 vdd.n2886 vdd.n2816 39.2114
R20218 vdd.n2890 vdd.n2817 39.2114
R20219 vdd.n2829 vdd.n2801 39.2114
R20220 vdd.n2833 vdd.n2802 39.2114
R20221 vdd.n2837 vdd.n2803 39.2114
R20222 vdd.n2841 vdd.n2804 39.2114
R20223 vdd.n2845 vdd.n2805 39.2114
R20224 vdd.n2849 vdd.n2806 39.2114
R20225 vdd.n2853 vdd.n2807 39.2114
R20226 vdd.n2857 vdd.n2808 39.2114
R20227 vdd.n2861 vdd.n2809 39.2114
R20228 vdd.n2865 vdd.n2810 39.2114
R20229 vdd.n2869 vdd.n2811 39.2114
R20230 vdd.n2873 vdd.n2812 39.2114
R20231 vdd.n2877 vdd.n2813 39.2114
R20232 vdd.n2881 vdd.n2814 39.2114
R20233 vdd.n2885 vdd.n2815 39.2114
R20234 vdd.n2889 vdd.n2816 39.2114
R20235 vdd.n2892 vdd.n2817 39.2114
R20236 vdd.n803 vdd.n798 39.2114
R20237 vdd.n3339 vdd.n3338 39.2114
R20238 vdd.n797 vdd.n795 39.2114
R20239 vdd.n3346 vdd.n3345 39.2114
R20240 vdd.n794 vdd.n792 39.2114
R20241 vdd.n3353 vdd.n3352 39.2114
R20242 vdd.n791 vdd.n789 39.2114
R20243 vdd.n3360 vdd.n3359 39.2114
R20244 vdd.n3363 vdd.n3362 39.2114
R20245 vdd.n3219 vdd.n3218 39.2114
R20246 vdd.n3224 vdd.n3223 39.2114
R20247 vdd.n3217 vdd.n3215 39.2114
R20248 vdd.n3231 vdd.n3230 39.2114
R20249 vdd.n3214 vdd.n3212 39.2114
R20250 vdd.n3238 vdd.n3237 39.2114
R20251 vdd.n3211 vdd.n3209 39.2114
R20252 vdd.n3245 vdd.n3244 39.2114
R20253 vdd.n2507 vdd.n1140 39.2114
R20254 vdd.n2501 vdd.n1142 39.2114
R20255 vdd.n2497 vdd.n1143 39.2114
R20256 vdd.n2493 vdd.n1144 39.2114
R20257 vdd.n2489 vdd.n1145 39.2114
R20258 vdd.n2485 vdd.n1146 39.2114
R20259 vdd.n2481 vdd.n1147 39.2114
R20260 vdd.n2477 vdd.n1148 39.2114
R20261 vdd.n1321 vdd.n1149 39.2114
R20262 vdd.n1325 vdd.n1150 39.2114
R20263 vdd.n1329 vdd.n1151 39.2114
R20264 vdd.n1333 vdd.n1152 39.2114
R20265 vdd.n1337 vdd.n1153 39.2114
R20266 vdd.n1341 vdd.n1154 39.2114
R20267 vdd.n1345 vdd.n1155 39.2114
R20268 vdd.n1350 vdd.n1156 39.2114
R20269 vdd.n1354 vdd.n1157 39.2114
R20270 vdd.n2717 vdd.n981 39.2114
R20271 vdd.n2722 vdd.n982 39.2114
R20272 vdd.n2726 vdd.n983 39.2114
R20273 vdd.n2730 vdd.n984 39.2114
R20274 vdd.n2734 vdd.n985 39.2114
R20275 vdd.n2738 vdd.n986 39.2114
R20276 vdd.n2742 vdd.n987 39.2114
R20277 vdd.n2746 vdd.n988 39.2114
R20278 vdd.n2750 vdd.n989 39.2114
R20279 vdd.n2754 vdd.n990 39.2114
R20280 vdd.n2758 vdd.n991 39.2114
R20281 vdd.n2762 vdd.n992 39.2114
R20282 vdd.n2766 vdd.n993 39.2114
R20283 vdd.n2770 vdd.n994 39.2114
R20284 vdd.n2774 vdd.n995 39.2114
R20285 vdd.n2778 vdd.n996 39.2114
R20286 vdd.n999 vdd.n997 39.2114
R20287 vdd.n3089 vdd.n962 39.2114
R20288 vdd.n3083 vdd.n2785 39.2114
R20289 vdd.n3079 vdd.n2786 39.2114
R20290 vdd.n3075 vdd.n2787 39.2114
R20291 vdd.n3071 vdd.n2788 39.2114
R20292 vdd.n3067 vdd.n2789 39.2114
R20293 vdd.n3063 vdd.n2790 39.2114
R20294 vdd.n3059 vdd.n2791 39.2114
R20295 vdd.n3055 vdd.n2792 39.2114
R20296 vdd.n3051 vdd.n2793 39.2114
R20297 vdd.n3047 vdd.n2794 39.2114
R20298 vdd.n3043 vdd.n2795 39.2114
R20299 vdd.n3039 vdd.n2796 39.2114
R20300 vdd.n3035 vdd.n2797 39.2114
R20301 vdd.n3031 vdd.n2798 39.2114
R20302 vdd.n3026 vdd.n2799 39.2114
R20303 vdd.n3022 vdd.n2800 39.2114
R20304 vdd.n3269 vdd.n3268 39.2114
R20305 vdd.n835 vdd.n831 39.2114
R20306 vdd.n3277 vdd.n3276 39.2114
R20307 vdd.n830 vdd.n828 39.2114
R20308 vdd.n3284 vdd.n3283 39.2114
R20309 vdd.n827 vdd.n825 39.2114
R20310 vdd.n3291 vdd.n3290 39.2114
R20311 vdd.n824 vdd.n822 39.2114
R20312 vdd.n3298 vdd.n3297 39.2114
R20313 vdd.n3302 vdd.n3301 39.2114
R20314 vdd.n821 vdd.n819 39.2114
R20315 vdd.n3309 vdd.n3308 39.2114
R20316 vdd.n818 vdd.n816 39.2114
R20317 vdd.n3316 vdd.n3315 39.2114
R20318 vdd.n815 vdd.n813 39.2114
R20319 vdd.n3323 vdd.n3322 39.2114
R20320 vdd.n3326 vdd.n3325 39.2114
R20321 vdd.n1008 vdd.n963 39.2114
R20322 vdd.n2706 vdd.n964 39.2114
R20323 vdd.n2702 vdd.n965 39.2114
R20324 vdd.n2698 vdd.n966 39.2114
R20325 vdd.n2694 vdd.n967 39.2114
R20326 vdd.n2690 vdd.n968 39.2114
R20327 vdd.n2686 vdd.n969 39.2114
R20328 vdd.n2682 vdd.n970 39.2114
R20329 vdd.n2678 vdd.n971 39.2114
R20330 vdd.n2674 vdd.n972 39.2114
R20331 vdd.n2670 vdd.n973 39.2114
R20332 vdd.n2666 vdd.n974 39.2114
R20333 vdd.n2662 vdd.n975 39.2114
R20334 vdd.n2658 vdd.n976 39.2114
R20335 vdd.n2654 vdd.n977 39.2114
R20336 vdd.n2650 vdd.n978 39.2114
R20337 vdd.n2646 vdd.n979 39.2114
R20338 vdd.n1280 vdd.n1158 39.2114
R20339 vdd.n1284 vdd.n1159 39.2114
R20340 vdd.n1288 vdd.n1160 39.2114
R20341 vdd.n1292 vdd.n1161 39.2114
R20342 vdd.n1296 vdd.n1162 39.2114
R20343 vdd.n1300 vdd.n1163 39.2114
R20344 vdd.n1304 vdd.n1164 39.2114
R20345 vdd.n1308 vdd.n1165 39.2114
R20346 vdd.n1312 vdd.n1166 39.2114
R20347 vdd.n1513 vdd.n1167 39.2114
R20348 vdd.n1510 vdd.n1168 39.2114
R20349 vdd.n1506 vdd.n1169 39.2114
R20350 vdd.n1502 vdd.n1170 39.2114
R20351 vdd.n1498 vdd.n1171 39.2114
R20352 vdd.n1494 vdd.n1172 39.2114
R20353 vdd.n1490 vdd.n1173 39.2114
R20354 vdd.n1486 vdd.n1174 39.2114
R20355 vdd.n2643 vdd.n979 39.2114
R20356 vdd.n2647 vdd.n978 39.2114
R20357 vdd.n2651 vdd.n977 39.2114
R20358 vdd.n2655 vdd.n976 39.2114
R20359 vdd.n2659 vdd.n975 39.2114
R20360 vdd.n2663 vdd.n974 39.2114
R20361 vdd.n2667 vdd.n973 39.2114
R20362 vdd.n2671 vdd.n972 39.2114
R20363 vdd.n2675 vdd.n971 39.2114
R20364 vdd.n2679 vdd.n970 39.2114
R20365 vdd.n2683 vdd.n969 39.2114
R20366 vdd.n2687 vdd.n968 39.2114
R20367 vdd.n2691 vdd.n967 39.2114
R20368 vdd.n2695 vdd.n966 39.2114
R20369 vdd.n2699 vdd.n965 39.2114
R20370 vdd.n2703 vdd.n964 39.2114
R20371 vdd.n2707 vdd.n963 39.2114
R20372 vdd.n1283 vdd.n1158 39.2114
R20373 vdd.n1287 vdd.n1159 39.2114
R20374 vdd.n1291 vdd.n1160 39.2114
R20375 vdd.n1295 vdd.n1161 39.2114
R20376 vdd.n1299 vdd.n1162 39.2114
R20377 vdd.n1303 vdd.n1163 39.2114
R20378 vdd.n1307 vdd.n1164 39.2114
R20379 vdd.n1311 vdd.n1165 39.2114
R20380 vdd.n1314 vdd.n1166 39.2114
R20381 vdd.n1511 vdd.n1167 39.2114
R20382 vdd.n1507 vdd.n1168 39.2114
R20383 vdd.n1503 vdd.n1169 39.2114
R20384 vdd.n1499 vdd.n1170 39.2114
R20385 vdd.n1495 vdd.n1171 39.2114
R20386 vdd.n1491 vdd.n1172 39.2114
R20387 vdd.n1487 vdd.n1173 39.2114
R20388 vdd.n1483 vdd.n1174 39.2114
R20389 vdd.n2364 vdd.n2363 37.2369
R20390 vdd.n2400 vdd.n1249 37.2369
R20391 vdd.n2439 vdd.n1209 37.2369
R20392 vdd.n3410 vdd.n769 37.2369
R20393 vdd.n3458 vdd.n3457 37.2369
R20394 vdd.n690 vdd.n689 37.2369
R20395 vdd.n1317 vdd.n1316 30.449
R20396 vdd.n1012 vdd.n1011 30.449
R20397 vdd.n1348 vdd.n1320 30.449
R20398 vdd.n2720 vdd.n1002 30.449
R20399 vdd.n2825 vdd.n2824 30.449
R20400 vdd.n3272 vdd.n833 30.449
R20401 vdd.n3028 vdd.n2821 30.449
R20402 vdd.n801 vdd.n800 30.449
R20403 vdd.n2510 vdd.n2509 29.8151
R20404 vdd.n2782 vdd.n1000 29.8151
R20405 vdd.n2715 vdd.n1003 29.8151
R20406 vdd.n1356 vdd.n1353 29.8151
R20407 vdd.n3023 vdd.n3020 29.8151
R20408 vdd.n3266 vdd.n3265 29.8151
R20409 vdd.n3092 vdd.n3091 29.8151
R20410 vdd.n3329 vdd.n3328 29.8151
R20411 vdd.n3248 vdd.n3247 29.8151
R20412 vdd.n3334 vdd.n802 29.8151
R20413 vdd.n2896 vdd.n2894 29.8151
R20414 vdd.n2827 vdd.n955 29.8151
R20415 vdd.n1281 vdd.n1132 29.8151
R20416 vdd.n2710 vdd.n2709 29.8151
R20417 vdd.n2642 vdd.n2641 29.8151
R20418 vdd.n1482 vdd.n1481 29.8151
R20419 vdd.n1873 vdd.n1680 22.2201
R20420 vdd.n2358 vdd.n1141 22.2201
R20421 vdd.n3495 vdd.n723 22.2201
R20422 vdd.n3627 vdd.n3626 22.2201
R20423 vdd.n1884 vdd.n1642 19.3944
R20424 vdd.n1884 vdd.n1640 19.3944
R20425 vdd.n1888 vdd.n1640 19.3944
R20426 vdd.n1888 vdd.n1630 19.3944
R20427 vdd.n1901 vdd.n1630 19.3944
R20428 vdd.n1901 vdd.n1628 19.3944
R20429 vdd.n1905 vdd.n1628 19.3944
R20430 vdd.n1905 vdd.n1620 19.3944
R20431 vdd.n1918 vdd.n1620 19.3944
R20432 vdd.n1918 vdd.n1618 19.3944
R20433 vdd.n1922 vdd.n1618 19.3944
R20434 vdd.n1922 vdd.n1607 19.3944
R20435 vdd.n1934 vdd.n1607 19.3944
R20436 vdd.n1934 vdd.n1605 19.3944
R20437 vdd.n1938 vdd.n1605 19.3944
R20438 vdd.n1938 vdd.n1596 19.3944
R20439 vdd.n1951 vdd.n1596 19.3944
R20440 vdd.n1951 vdd.n1594 19.3944
R20441 vdd.n1955 vdd.n1594 19.3944
R20442 vdd.n1955 vdd.n1585 19.3944
R20443 vdd.n2274 vdd.n1585 19.3944
R20444 vdd.n2274 vdd.n1583 19.3944
R20445 vdd.n2278 vdd.n1583 19.3944
R20446 vdd.n2278 vdd.n1573 19.3944
R20447 vdd.n2291 vdd.n1573 19.3944
R20448 vdd.n2291 vdd.n1571 19.3944
R20449 vdd.n2295 vdd.n1571 19.3944
R20450 vdd.n2295 vdd.n1563 19.3944
R20451 vdd.n2308 vdd.n1563 19.3944
R20452 vdd.n2308 vdd.n1561 19.3944
R20453 vdd.n2312 vdd.n1561 19.3944
R20454 vdd.n2312 vdd.n1550 19.3944
R20455 vdd.n2324 vdd.n1550 19.3944
R20456 vdd.n2324 vdd.n1548 19.3944
R20457 vdd.n2328 vdd.n1548 19.3944
R20458 vdd.n2328 vdd.n1540 19.3944
R20459 vdd.n2341 vdd.n1540 19.3944
R20460 vdd.n2341 vdd.n1537 19.3944
R20461 vdd.n2347 vdd.n1537 19.3944
R20462 vdd.n2347 vdd.n1538 19.3944
R20463 vdd.n1538 vdd.n1528 19.3944
R20464 vdd.n1808 vdd.n1743 19.3944
R20465 vdd.n1804 vdd.n1743 19.3944
R20466 vdd.n1804 vdd.n1803 19.3944
R20467 vdd.n1803 vdd.n1802 19.3944
R20468 vdd.n1802 vdd.n1749 19.3944
R20469 vdd.n1798 vdd.n1749 19.3944
R20470 vdd.n1798 vdd.n1797 19.3944
R20471 vdd.n1797 vdd.n1796 19.3944
R20472 vdd.n1796 vdd.n1755 19.3944
R20473 vdd.n1792 vdd.n1755 19.3944
R20474 vdd.n1792 vdd.n1791 19.3944
R20475 vdd.n1791 vdd.n1790 19.3944
R20476 vdd.n1790 vdd.n1761 19.3944
R20477 vdd.n1786 vdd.n1761 19.3944
R20478 vdd.n1786 vdd.n1785 19.3944
R20479 vdd.n1785 vdd.n1784 19.3944
R20480 vdd.n1784 vdd.n1767 19.3944
R20481 vdd.n1780 vdd.n1767 19.3944
R20482 vdd.n1780 vdd.n1779 19.3944
R20483 vdd.n1779 vdd.n1778 19.3944
R20484 vdd.n1843 vdd.n1842 19.3944
R20485 vdd.n1842 vdd.n1841 19.3944
R20486 vdd.n1841 vdd.n1714 19.3944
R20487 vdd.n1837 vdd.n1714 19.3944
R20488 vdd.n1837 vdd.n1836 19.3944
R20489 vdd.n1836 vdd.n1835 19.3944
R20490 vdd.n1835 vdd.n1720 19.3944
R20491 vdd.n1831 vdd.n1720 19.3944
R20492 vdd.n1831 vdd.n1830 19.3944
R20493 vdd.n1830 vdd.n1829 19.3944
R20494 vdd.n1829 vdd.n1726 19.3944
R20495 vdd.n1825 vdd.n1726 19.3944
R20496 vdd.n1825 vdd.n1824 19.3944
R20497 vdd.n1824 vdd.n1823 19.3944
R20498 vdd.n1823 vdd.n1732 19.3944
R20499 vdd.n1819 vdd.n1732 19.3944
R20500 vdd.n1819 vdd.n1818 19.3944
R20501 vdd.n1818 vdd.n1817 19.3944
R20502 vdd.n1817 vdd.n1738 19.3944
R20503 vdd.n1813 vdd.n1738 19.3944
R20504 vdd.n1876 vdd.n1647 19.3944
R20505 vdd.n1871 vdd.n1647 19.3944
R20506 vdd.n1871 vdd.n1682 19.3944
R20507 vdd.n1867 vdd.n1682 19.3944
R20508 vdd.n1867 vdd.n1866 19.3944
R20509 vdd.n1866 vdd.n1865 19.3944
R20510 vdd.n1865 vdd.n1688 19.3944
R20511 vdd.n1861 vdd.n1688 19.3944
R20512 vdd.n1861 vdd.n1860 19.3944
R20513 vdd.n1860 vdd.n1859 19.3944
R20514 vdd.n1859 vdd.n1694 19.3944
R20515 vdd.n1855 vdd.n1694 19.3944
R20516 vdd.n1855 vdd.n1854 19.3944
R20517 vdd.n1854 vdd.n1853 19.3944
R20518 vdd.n1853 vdd.n1700 19.3944
R20519 vdd.n1849 vdd.n1700 19.3944
R20520 vdd.n1849 vdd.n1848 19.3944
R20521 vdd.n1848 vdd.n1847 19.3944
R20522 vdd.n2396 vdd.n1247 19.3944
R20523 vdd.n2396 vdd.n1253 19.3944
R20524 vdd.n2391 vdd.n1253 19.3944
R20525 vdd.n2391 vdd.n2390 19.3944
R20526 vdd.n2390 vdd.n2389 19.3944
R20527 vdd.n2389 vdd.n1260 19.3944
R20528 vdd.n2384 vdd.n1260 19.3944
R20529 vdd.n2384 vdd.n2383 19.3944
R20530 vdd.n2383 vdd.n2382 19.3944
R20531 vdd.n2382 vdd.n1267 19.3944
R20532 vdd.n2377 vdd.n1267 19.3944
R20533 vdd.n2377 vdd.n2376 19.3944
R20534 vdd.n2376 vdd.n2375 19.3944
R20535 vdd.n2375 vdd.n1274 19.3944
R20536 vdd.n2370 vdd.n1274 19.3944
R20537 vdd.n2370 vdd.n2369 19.3944
R20538 vdd.n1521 vdd.n1279 19.3944
R20539 vdd.n2365 vdd.n1518 19.3944
R20540 vdd.n2435 vdd.n1207 19.3944
R20541 vdd.n2435 vdd.n1213 19.3944
R20542 vdd.n2430 vdd.n1213 19.3944
R20543 vdd.n2430 vdd.n2429 19.3944
R20544 vdd.n2429 vdd.n2428 19.3944
R20545 vdd.n2428 vdd.n1220 19.3944
R20546 vdd.n2423 vdd.n1220 19.3944
R20547 vdd.n2423 vdd.n2422 19.3944
R20548 vdd.n2422 vdd.n2421 19.3944
R20549 vdd.n2421 vdd.n1227 19.3944
R20550 vdd.n2416 vdd.n1227 19.3944
R20551 vdd.n2416 vdd.n2415 19.3944
R20552 vdd.n2415 vdd.n2414 19.3944
R20553 vdd.n2414 vdd.n1234 19.3944
R20554 vdd.n2409 vdd.n1234 19.3944
R20555 vdd.n2409 vdd.n2408 19.3944
R20556 vdd.n2408 vdd.n2407 19.3944
R20557 vdd.n2407 vdd.n1241 19.3944
R20558 vdd.n2402 vdd.n1241 19.3944
R20559 vdd.n2402 vdd.n2401 19.3944
R20560 vdd.n2472 vdd.n1182 19.3944
R20561 vdd.n2472 vdd.n1183 19.3944
R20562 vdd.n2467 vdd.n2466 19.3944
R20563 vdd.n2462 vdd.n2461 19.3944
R20564 vdd.n2461 vdd.n2460 19.3944
R20565 vdd.n2460 vdd.n1187 19.3944
R20566 vdd.n2455 vdd.n1187 19.3944
R20567 vdd.n2455 vdd.n2454 19.3944
R20568 vdd.n2454 vdd.n2453 19.3944
R20569 vdd.n2453 vdd.n1194 19.3944
R20570 vdd.n2448 vdd.n1194 19.3944
R20571 vdd.n2448 vdd.n2447 19.3944
R20572 vdd.n2447 vdd.n2446 19.3944
R20573 vdd.n2446 vdd.n1201 19.3944
R20574 vdd.n2441 vdd.n1201 19.3944
R20575 vdd.n2441 vdd.n2440 19.3944
R20576 vdd.n1880 vdd.n1645 19.3944
R20577 vdd.n1880 vdd.n1636 19.3944
R20578 vdd.n1893 vdd.n1636 19.3944
R20579 vdd.n1893 vdd.n1634 19.3944
R20580 vdd.n1897 vdd.n1634 19.3944
R20581 vdd.n1897 vdd.n1625 19.3944
R20582 vdd.n1910 vdd.n1625 19.3944
R20583 vdd.n1910 vdd.n1623 19.3944
R20584 vdd.n1914 vdd.n1623 19.3944
R20585 vdd.n1914 vdd.n1614 19.3944
R20586 vdd.n1926 vdd.n1614 19.3944
R20587 vdd.n1926 vdd.n1612 19.3944
R20588 vdd.n1930 vdd.n1612 19.3944
R20589 vdd.n1930 vdd.n1602 19.3944
R20590 vdd.n1943 vdd.n1602 19.3944
R20591 vdd.n1943 vdd.n1600 19.3944
R20592 vdd.n1947 vdd.n1600 19.3944
R20593 vdd.n1947 vdd.n1591 19.3944
R20594 vdd.n1959 vdd.n1591 19.3944
R20595 vdd.n1959 vdd.n1589 19.3944
R20596 vdd.n2270 vdd.n1589 19.3944
R20597 vdd.n2270 vdd.n1579 19.3944
R20598 vdd.n2283 vdd.n1579 19.3944
R20599 vdd.n2283 vdd.n1577 19.3944
R20600 vdd.n2287 vdd.n1577 19.3944
R20601 vdd.n2287 vdd.n1568 19.3944
R20602 vdd.n2300 vdd.n1568 19.3944
R20603 vdd.n2300 vdd.n1566 19.3944
R20604 vdd.n2304 vdd.n1566 19.3944
R20605 vdd.n2304 vdd.n1557 19.3944
R20606 vdd.n2316 vdd.n1557 19.3944
R20607 vdd.n2316 vdd.n1555 19.3944
R20608 vdd.n2320 vdd.n1555 19.3944
R20609 vdd.n2320 vdd.n1545 19.3944
R20610 vdd.n2333 vdd.n1545 19.3944
R20611 vdd.n2333 vdd.n1543 19.3944
R20612 vdd.n2337 vdd.n1543 19.3944
R20613 vdd.n2337 vdd.n1533 19.3944
R20614 vdd.n2352 vdd.n1533 19.3944
R20615 vdd.n2352 vdd.n1531 19.3944
R20616 vdd.n2356 vdd.n1531 19.3944
R20617 vdd.n3501 vdd.n686 19.3944
R20618 vdd.n3501 vdd.n676 19.3944
R20619 vdd.n3513 vdd.n676 19.3944
R20620 vdd.n3513 vdd.n674 19.3944
R20621 vdd.n3517 vdd.n674 19.3944
R20622 vdd.n3517 vdd.n666 19.3944
R20623 vdd.n3530 vdd.n666 19.3944
R20624 vdd.n3530 vdd.n664 19.3944
R20625 vdd.n3534 vdd.n664 19.3944
R20626 vdd.n3534 vdd.n653 19.3944
R20627 vdd.n3546 vdd.n653 19.3944
R20628 vdd.n3546 vdd.n651 19.3944
R20629 vdd.n3550 vdd.n651 19.3944
R20630 vdd.n3550 vdd.n642 19.3944
R20631 vdd.n3563 vdd.n642 19.3944
R20632 vdd.n3563 vdd.n640 19.3944
R20633 vdd.n3570 vdd.n640 19.3944
R20634 vdd.n3570 vdd.n3569 19.3944
R20635 vdd.n3569 vdd.n631 19.3944
R20636 vdd.n3583 vdd.n631 19.3944
R20637 vdd.n3584 vdd.n3583 19.3944
R20638 vdd.n3584 vdd.n629 19.3944
R20639 vdd.n3588 vdd.n629 19.3944
R20640 vdd.n3590 vdd.n3588 19.3944
R20641 vdd.n3591 vdd.n3590 19.3944
R20642 vdd.n3591 vdd.n627 19.3944
R20643 vdd.n3595 vdd.n627 19.3944
R20644 vdd.n3597 vdd.n3595 19.3944
R20645 vdd.n3598 vdd.n3597 19.3944
R20646 vdd.n3598 vdd.n625 19.3944
R20647 vdd.n3602 vdd.n625 19.3944
R20648 vdd.n3605 vdd.n3602 19.3944
R20649 vdd.n3606 vdd.n3605 19.3944
R20650 vdd.n3606 vdd.n623 19.3944
R20651 vdd.n3610 vdd.n623 19.3944
R20652 vdd.n3612 vdd.n3610 19.3944
R20653 vdd.n3613 vdd.n3612 19.3944
R20654 vdd.n3613 vdd.n621 19.3944
R20655 vdd.n3617 vdd.n621 19.3944
R20656 vdd.n3619 vdd.n3617 19.3944
R20657 vdd.n3620 vdd.n3619 19.3944
R20658 vdd.n569 vdd.n438 19.3944
R20659 vdd.n575 vdd.n438 19.3944
R20660 vdd.n576 vdd.n575 19.3944
R20661 vdd.n579 vdd.n576 19.3944
R20662 vdd.n579 vdd.n436 19.3944
R20663 vdd.n585 vdd.n436 19.3944
R20664 vdd.n586 vdd.n585 19.3944
R20665 vdd.n589 vdd.n586 19.3944
R20666 vdd.n589 vdd.n434 19.3944
R20667 vdd.n595 vdd.n434 19.3944
R20668 vdd.n596 vdd.n595 19.3944
R20669 vdd.n599 vdd.n596 19.3944
R20670 vdd.n599 vdd.n432 19.3944
R20671 vdd.n605 vdd.n432 19.3944
R20672 vdd.n606 vdd.n605 19.3944
R20673 vdd.n609 vdd.n606 19.3944
R20674 vdd.n609 vdd.n430 19.3944
R20675 vdd.n615 vdd.n430 19.3944
R20676 vdd.n617 vdd.n615 19.3944
R20677 vdd.n618 vdd.n617 19.3944
R20678 vdd.n516 vdd.n515 19.3944
R20679 vdd.n519 vdd.n516 19.3944
R20680 vdd.n519 vdd.n450 19.3944
R20681 vdd.n525 vdd.n450 19.3944
R20682 vdd.n526 vdd.n525 19.3944
R20683 vdd.n529 vdd.n526 19.3944
R20684 vdd.n529 vdd.n448 19.3944
R20685 vdd.n535 vdd.n448 19.3944
R20686 vdd.n536 vdd.n535 19.3944
R20687 vdd.n539 vdd.n536 19.3944
R20688 vdd.n539 vdd.n446 19.3944
R20689 vdd.n545 vdd.n446 19.3944
R20690 vdd.n546 vdd.n545 19.3944
R20691 vdd.n549 vdd.n546 19.3944
R20692 vdd.n549 vdd.n444 19.3944
R20693 vdd.n555 vdd.n444 19.3944
R20694 vdd.n556 vdd.n555 19.3944
R20695 vdd.n559 vdd.n556 19.3944
R20696 vdd.n559 vdd.n442 19.3944
R20697 vdd.n565 vdd.n442 19.3944
R20698 vdd.n466 vdd.n465 19.3944
R20699 vdd.n469 vdd.n466 19.3944
R20700 vdd.n469 vdd.n462 19.3944
R20701 vdd.n475 vdd.n462 19.3944
R20702 vdd.n476 vdd.n475 19.3944
R20703 vdd.n479 vdd.n476 19.3944
R20704 vdd.n479 vdd.n460 19.3944
R20705 vdd.n485 vdd.n460 19.3944
R20706 vdd.n486 vdd.n485 19.3944
R20707 vdd.n489 vdd.n486 19.3944
R20708 vdd.n489 vdd.n458 19.3944
R20709 vdd.n495 vdd.n458 19.3944
R20710 vdd.n496 vdd.n495 19.3944
R20711 vdd.n499 vdd.n496 19.3944
R20712 vdd.n499 vdd.n456 19.3944
R20713 vdd.n505 vdd.n456 19.3944
R20714 vdd.n506 vdd.n505 19.3944
R20715 vdd.n509 vdd.n506 19.3944
R20716 vdd.n3505 vdd.n683 19.3944
R20717 vdd.n3505 vdd.n681 19.3944
R20718 vdd.n3509 vdd.n681 19.3944
R20719 vdd.n3509 vdd.n671 19.3944
R20720 vdd.n3522 vdd.n671 19.3944
R20721 vdd.n3522 vdd.n669 19.3944
R20722 vdd.n3526 vdd.n669 19.3944
R20723 vdd.n3526 vdd.n660 19.3944
R20724 vdd.n3538 vdd.n660 19.3944
R20725 vdd.n3538 vdd.n658 19.3944
R20726 vdd.n3542 vdd.n658 19.3944
R20727 vdd.n3542 vdd.n648 19.3944
R20728 vdd.n3555 vdd.n648 19.3944
R20729 vdd.n3555 vdd.n646 19.3944
R20730 vdd.n3559 vdd.n646 19.3944
R20731 vdd.n3559 vdd.n637 19.3944
R20732 vdd.n3574 vdd.n637 19.3944
R20733 vdd.n3574 vdd.n635 19.3944
R20734 vdd.n3578 vdd.n635 19.3944
R20735 vdd.n3578 vdd.n336 19.3944
R20736 vdd.n3669 vdd.n336 19.3944
R20737 vdd.n3669 vdd.n337 19.3944
R20738 vdd.n3663 vdd.n337 19.3944
R20739 vdd.n3663 vdd.n3662 19.3944
R20740 vdd.n3662 vdd.n3661 19.3944
R20741 vdd.n3661 vdd.n349 19.3944
R20742 vdd.n3655 vdd.n349 19.3944
R20743 vdd.n3655 vdd.n3654 19.3944
R20744 vdd.n3654 vdd.n3653 19.3944
R20745 vdd.n3653 vdd.n359 19.3944
R20746 vdd.n3647 vdd.n359 19.3944
R20747 vdd.n3647 vdd.n3646 19.3944
R20748 vdd.n3646 vdd.n3645 19.3944
R20749 vdd.n3645 vdd.n370 19.3944
R20750 vdd.n3639 vdd.n370 19.3944
R20751 vdd.n3639 vdd.n3638 19.3944
R20752 vdd.n3638 vdd.n3637 19.3944
R20753 vdd.n3637 vdd.n381 19.3944
R20754 vdd.n3631 vdd.n381 19.3944
R20755 vdd.n3631 vdd.n3630 19.3944
R20756 vdd.n3630 vdd.n3629 19.3944
R20757 vdd.n3452 vdd.n747 19.3944
R20758 vdd.n3452 vdd.n3449 19.3944
R20759 vdd.n3449 vdd.n3446 19.3944
R20760 vdd.n3446 vdd.n3445 19.3944
R20761 vdd.n3445 vdd.n3442 19.3944
R20762 vdd.n3442 vdd.n3441 19.3944
R20763 vdd.n3441 vdd.n3438 19.3944
R20764 vdd.n3438 vdd.n3437 19.3944
R20765 vdd.n3437 vdd.n3434 19.3944
R20766 vdd.n3434 vdd.n3433 19.3944
R20767 vdd.n3433 vdd.n3430 19.3944
R20768 vdd.n3430 vdd.n3429 19.3944
R20769 vdd.n3429 vdd.n3426 19.3944
R20770 vdd.n3426 vdd.n3425 19.3944
R20771 vdd.n3425 vdd.n3422 19.3944
R20772 vdd.n3422 vdd.n3421 19.3944
R20773 vdd.n3421 vdd.n3418 19.3944
R20774 vdd.n3418 vdd.n3417 19.3944
R20775 vdd.n3417 vdd.n3414 19.3944
R20776 vdd.n3414 vdd.n3413 19.3944
R20777 vdd.n3492 vdd.n3491 19.3944
R20778 vdd.n3491 vdd.n3490 19.3944
R20779 vdd.n732 vdd.n729 19.3944
R20780 vdd.n3486 vdd.n3485 19.3944
R20781 vdd.n3485 vdd.n3482 19.3944
R20782 vdd.n3482 vdd.n3481 19.3944
R20783 vdd.n3481 vdd.n3478 19.3944
R20784 vdd.n3478 vdd.n3477 19.3944
R20785 vdd.n3477 vdd.n3474 19.3944
R20786 vdd.n3474 vdd.n3473 19.3944
R20787 vdd.n3473 vdd.n3470 19.3944
R20788 vdd.n3470 vdd.n3469 19.3944
R20789 vdd.n3469 vdd.n3466 19.3944
R20790 vdd.n3466 vdd.n3465 19.3944
R20791 vdd.n3465 vdd.n3462 19.3944
R20792 vdd.n3462 vdd.n3461 19.3944
R20793 vdd.n3406 vdd.n767 19.3944
R20794 vdd.n3406 vdd.n3403 19.3944
R20795 vdd.n3403 vdd.n3400 19.3944
R20796 vdd.n3400 vdd.n3399 19.3944
R20797 vdd.n3399 vdd.n3396 19.3944
R20798 vdd.n3396 vdd.n3395 19.3944
R20799 vdd.n3395 vdd.n3392 19.3944
R20800 vdd.n3392 vdd.n3391 19.3944
R20801 vdd.n3391 vdd.n3388 19.3944
R20802 vdd.n3388 vdd.n3387 19.3944
R20803 vdd.n3387 vdd.n3384 19.3944
R20804 vdd.n3384 vdd.n3383 19.3944
R20805 vdd.n3383 vdd.n3380 19.3944
R20806 vdd.n3380 vdd.n3379 19.3944
R20807 vdd.n3379 vdd.n3376 19.3944
R20808 vdd.n3376 vdd.n3375 19.3944
R20809 vdd.n3372 vdd.n3371 19.3944
R20810 vdd.n3368 vdd.n3367 19.3944
R20811 vdd.n1812 vdd.n1808 19.0066
R20812 vdd.n2400 vdd.n1247 19.0066
R20813 vdd.n569 vdd.n566 19.0066
R20814 vdd.n3410 vdd.n767 19.0066
R20815 vdd.n1316 vdd.n1315 16.0975
R20816 vdd.n1011 vdd.n1010 16.0975
R20817 vdd.n1773 vdd.n1772 16.0975
R20818 vdd.n1811 vdd.n1810 16.0975
R20819 vdd.n1707 vdd.n1706 16.0975
R20820 vdd.n2363 vdd.n2362 16.0975
R20821 vdd.n1249 vdd.n1248 16.0975
R20822 vdd.n1209 vdd.n1208 16.0975
R20823 vdd.n1320 vdd.n1319 16.0975
R20824 vdd.n1002 vdd.n1001 16.0975
R20825 vdd.n2824 vdd.n2823 16.0975
R20826 vdd.n427 vdd.n426 16.0975
R20827 vdd.n441 vdd.n440 16.0975
R20828 vdd.n453 vdd.n452 16.0975
R20829 vdd.n769 vdd.n768 16.0975
R20830 vdd.n3457 vdd.n3456 16.0975
R20831 vdd.n833 vdd.n832 16.0975
R20832 vdd.n2821 vdd.n2820 16.0975
R20833 vdd.n689 vdd.n688 16.0975
R20834 vdd.n800 vdd.n799 16.0975
R20835 vdd.t264 vdd.n2784 15.4182
R20836 vdd.n3088 vdd.t251 15.4182
R20837 vdd.n28 vdd.n27 14.6072
R20838 vdd.n328 vdd.n293 13.1884
R20839 vdd.n269 vdd.n234 13.1884
R20840 vdd.n226 vdd.n191 13.1884
R20841 vdd.n167 vdd.n132 13.1884
R20842 vdd.n125 vdd.n90 13.1884
R20843 vdd.n66 vdd.n31 13.1884
R20844 vdd.n2202 vdd.n2167 13.1884
R20845 vdd.n2261 vdd.n2226 13.1884
R20846 vdd.n2100 vdd.n2065 13.1884
R20847 vdd.n2159 vdd.n2124 13.1884
R20848 vdd.n1999 vdd.n1964 13.1884
R20849 vdd.n2058 vdd.n2023 13.1884
R20850 vdd.n2506 vdd.n1134 13.1509
R20851 vdd.n3331 vdd.n692 13.1509
R20852 vdd.n1843 vdd.n1708 12.9944
R20853 vdd.n1847 vdd.n1708 12.9944
R20854 vdd.n2439 vdd.n1207 12.9944
R20855 vdd.n2440 vdd.n2439 12.9944
R20856 vdd.n515 vdd.n454 12.9944
R20857 vdd.n509 vdd.n454 12.9944
R20858 vdd.n3458 vdd.n747 12.9944
R20859 vdd.n3461 vdd.n3458 12.9944
R20860 vdd.n329 vdd.n291 12.8005
R20861 vdd.n324 vdd.n295 12.8005
R20862 vdd.n270 vdd.n232 12.8005
R20863 vdd.n265 vdd.n236 12.8005
R20864 vdd.n227 vdd.n189 12.8005
R20865 vdd.n222 vdd.n193 12.8005
R20866 vdd.n168 vdd.n130 12.8005
R20867 vdd.n163 vdd.n134 12.8005
R20868 vdd.n126 vdd.n88 12.8005
R20869 vdd.n121 vdd.n92 12.8005
R20870 vdd.n67 vdd.n29 12.8005
R20871 vdd.n62 vdd.n33 12.8005
R20872 vdd.n2203 vdd.n2165 12.8005
R20873 vdd.n2198 vdd.n2169 12.8005
R20874 vdd.n2262 vdd.n2224 12.8005
R20875 vdd.n2257 vdd.n2228 12.8005
R20876 vdd.n2101 vdd.n2063 12.8005
R20877 vdd.n2096 vdd.n2067 12.8005
R20878 vdd.n2160 vdd.n2122 12.8005
R20879 vdd.n2155 vdd.n2126 12.8005
R20880 vdd.n2000 vdd.n1962 12.8005
R20881 vdd.n1995 vdd.n1966 12.8005
R20882 vdd.n2059 vdd.n2021 12.8005
R20883 vdd.n2054 vdd.n2025 12.8005
R20884 vdd.n323 vdd.n296 12.0247
R20885 vdd.n264 vdd.n237 12.0247
R20886 vdd.n221 vdd.n194 12.0247
R20887 vdd.n162 vdd.n135 12.0247
R20888 vdd.n120 vdd.n93 12.0247
R20889 vdd.n61 vdd.n34 12.0247
R20890 vdd.n2197 vdd.n2170 12.0247
R20891 vdd.n2256 vdd.n2229 12.0247
R20892 vdd.n2095 vdd.n2068 12.0247
R20893 vdd.n2154 vdd.n2127 12.0247
R20894 vdd.n1994 vdd.n1967 12.0247
R20895 vdd.n2053 vdd.n2026 12.0247
R20896 vdd.n1882 vdd.n1638 11.337
R20897 vdd.n1891 vdd.n1638 11.337
R20898 vdd.n1891 vdd.n1890 11.337
R20899 vdd.n1899 vdd.n1632 11.337
R20900 vdd.n1908 vdd.n1907 11.337
R20901 vdd.n1924 vdd.n1616 11.337
R20902 vdd.n1932 vdd.n1609 11.337
R20903 vdd.n1941 vdd.n1940 11.337
R20904 vdd.n1949 vdd.n1598 11.337
R20905 vdd.n2272 vdd.n1587 11.337
R20906 vdd.n2281 vdd.n1581 11.337
R20907 vdd.n2289 vdd.n1575 11.337
R20908 vdd.n2298 vdd.n2297 11.337
R20909 vdd.n2314 vdd.n1559 11.337
R20910 vdd.n2322 vdd.n1552 11.337
R20911 vdd.n2331 vdd.n2330 11.337
R20912 vdd.n2339 vdd.n1535 11.337
R20913 vdd.n2350 vdd.n1535 11.337
R20914 vdd.n2350 vdd.n2349 11.337
R20915 vdd.n3503 vdd.n678 11.337
R20916 vdd.n3511 vdd.n678 11.337
R20917 vdd.n3511 vdd.n679 11.337
R20918 vdd.n3520 vdd.n3519 11.337
R20919 vdd.n3536 vdd.n662 11.337
R20920 vdd.n3544 vdd.n655 11.337
R20921 vdd.n3553 vdd.n3552 11.337
R20922 vdd.n3561 vdd.n644 11.337
R20923 vdd.n3580 vdd.n633 11.337
R20924 vdd.n3667 vdd.n340 11.337
R20925 vdd.n3665 vdd.n344 11.337
R20926 vdd.n3659 vdd.n3658 11.337
R20927 vdd.n3651 vdd.n361 11.337
R20928 vdd.n3650 vdd.n3649 11.337
R20929 vdd.n3643 vdd.n3642 11.337
R20930 vdd.n3641 vdd.n375 11.337
R20931 vdd.n3635 vdd.n3634 11.337
R20932 vdd.n3634 vdd.n3633 11.337
R20933 vdd.n3633 vdd.n386 11.337
R20934 vdd.n320 vdd.n319 11.249
R20935 vdd.n261 vdd.n260 11.249
R20936 vdd.n218 vdd.n217 11.249
R20937 vdd.n159 vdd.n158 11.249
R20938 vdd.n117 vdd.n116 11.249
R20939 vdd.n58 vdd.n57 11.249
R20940 vdd.n2194 vdd.n2193 11.249
R20941 vdd.n2253 vdd.n2252 11.249
R20942 vdd.n2092 vdd.n2091 11.249
R20943 vdd.n2151 vdd.n2150 11.249
R20944 vdd.n1991 vdd.n1990 11.249
R20945 vdd.n2050 vdd.n2049 11.249
R20946 vdd.n1680 vdd.t224 11.2237
R20947 vdd.n3627 vdd.t173 11.2237
R20948 vdd.t96 vdd.n1553 10.7702
R20949 vdd.n3528 vdd.t22 10.7702
R20950 vdd.n305 vdd.n304 10.7238
R20951 vdd.n246 vdd.n245 10.7238
R20952 vdd.n203 vdd.n202 10.7238
R20953 vdd.n144 vdd.n143 10.7238
R20954 vdd.n102 vdd.n101 10.7238
R20955 vdd.n43 vdd.n42 10.7238
R20956 vdd.n2179 vdd.n2178 10.7238
R20957 vdd.n2238 vdd.n2237 10.7238
R20958 vdd.n2077 vdd.n2076 10.7238
R20959 vdd.n2136 vdd.n2135 10.7238
R20960 vdd.n1976 vdd.n1975 10.7238
R20961 vdd.n2035 vdd.n2034 10.7238
R20962 vdd.n2511 vdd.n2510 10.6151
R20963 vdd.n2511 vdd.n1127 10.6151
R20964 vdd.n2521 vdd.n1127 10.6151
R20965 vdd.n2522 vdd.n2521 10.6151
R20966 vdd.n2523 vdd.n2522 10.6151
R20967 vdd.n2523 vdd.n1114 10.6151
R20968 vdd.n2533 vdd.n1114 10.6151
R20969 vdd.n2534 vdd.n2533 10.6151
R20970 vdd.n2535 vdd.n2534 10.6151
R20971 vdd.n2535 vdd.n1102 10.6151
R20972 vdd.n2545 vdd.n1102 10.6151
R20973 vdd.n2546 vdd.n2545 10.6151
R20974 vdd.n2547 vdd.n2546 10.6151
R20975 vdd.n2547 vdd.n1091 10.6151
R20976 vdd.n2557 vdd.n1091 10.6151
R20977 vdd.n2558 vdd.n2557 10.6151
R20978 vdd.n2559 vdd.n2558 10.6151
R20979 vdd.n2559 vdd.n1078 10.6151
R20980 vdd.n2569 vdd.n1078 10.6151
R20981 vdd.n2570 vdd.n2569 10.6151
R20982 vdd.n2571 vdd.n2570 10.6151
R20983 vdd.n2571 vdd.n1066 10.6151
R20984 vdd.n2582 vdd.n1066 10.6151
R20985 vdd.n2583 vdd.n2582 10.6151
R20986 vdd.n2584 vdd.n2583 10.6151
R20987 vdd.n2584 vdd.n1054 10.6151
R20988 vdd.n2594 vdd.n1054 10.6151
R20989 vdd.n2595 vdd.n2594 10.6151
R20990 vdd.n2596 vdd.n2595 10.6151
R20991 vdd.n2596 vdd.n1042 10.6151
R20992 vdd.n2606 vdd.n1042 10.6151
R20993 vdd.n2607 vdd.n2606 10.6151
R20994 vdd.n2608 vdd.n2607 10.6151
R20995 vdd.n2608 vdd.n1032 10.6151
R20996 vdd.n2618 vdd.n1032 10.6151
R20997 vdd.n2619 vdd.n2618 10.6151
R20998 vdd.n2620 vdd.n2619 10.6151
R20999 vdd.n2620 vdd.n1019 10.6151
R21000 vdd.n2632 vdd.n1019 10.6151
R21001 vdd.n2633 vdd.n2632 10.6151
R21002 vdd.n2635 vdd.n2633 10.6151
R21003 vdd.n2635 vdd.n2634 10.6151
R21004 vdd.n2634 vdd.n1000 10.6151
R21005 vdd.n2782 vdd.n2781 10.6151
R21006 vdd.n2781 vdd.n2780 10.6151
R21007 vdd.n2780 vdd.n2777 10.6151
R21008 vdd.n2777 vdd.n2776 10.6151
R21009 vdd.n2776 vdd.n2773 10.6151
R21010 vdd.n2773 vdd.n2772 10.6151
R21011 vdd.n2772 vdd.n2769 10.6151
R21012 vdd.n2769 vdd.n2768 10.6151
R21013 vdd.n2768 vdd.n2765 10.6151
R21014 vdd.n2765 vdd.n2764 10.6151
R21015 vdd.n2764 vdd.n2761 10.6151
R21016 vdd.n2761 vdd.n2760 10.6151
R21017 vdd.n2760 vdd.n2757 10.6151
R21018 vdd.n2757 vdd.n2756 10.6151
R21019 vdd.n2756 vdd.n2753 10.6151
R21020 vdd.n2753 vdd.n2752 10.6151
R21021 vdd.n2752 vdd.n2749 10.6151
R21022 vdd.n2749 vdd.n2748 10.6151
R21023 vdd.n2748 vdd.n2745 10.6151
R21024 vdd.n2745 vdd.n2744 10.6151
R21025 vdd.n2744 vdd.n2741 10.6151
R21026 vdd.n2741 vdd.n2740 10.6151
R21027 vdd.n2740 vdd.n2737 10.6151
R21028 vdd.n2737 vdd.n2736 10.6151
R21029 vdd.n2736 vdd.n2733 10.6151
R21030 vdd.n2733 vdd.n2732 10.6151
R21031 vdd.n2732 vdd.n2729 10.6151
R21032 vdd.n2729 vdd.n2728 10.6151
R21033 vdd.n2728 vdd.n2725 10.6151
R21034 vdd.n2725 vdd.n2724 10.6151
R21035 vdd.n2724 vdd.n2721 10.6151
R21036 vdd.n2719 vdd.n2716 10.6151
R21037 vdd.n2716 vdd.n2715 10.6151
R21038 vdd.n1357 vdd.n1356 10.6151
R21039 vdd.n1359 vdd.n1357 10.6151
R21040 vdd.n1360 vdd.n1359 10.6151
R21041 vdd.n1362 vdd.n1360 10.6151
R21042 vdd.n1363 vdd.n1362 10.6151
R21043 vdd.n1365 vdd.n1363 10.6151
R21044 vdd.n1366 vdd.n1365 10.6151
R21045 vdd.n1368 vdd.n1366 10.6151
R21046 vdd.n1369 vdd.n1368 10.6151
R21047 vdd.n1371 vdd.n1369 10.6151
R21048 vdd.n1372 vdd.n1371 10.6151
R21049 vdd.n1374 vdd.n1372 10.6151
R21050 vdd.n1375 vdd.n1374 10.6151
R21051 vdd.n1377 vdd.n1375 10.6151
R21052 vdd.n1378 vdd.n1377 10.6151
R21053 vdd.n1380 vdd.n1378 10.6151
R21054 vdd.n1381 vdd.n1380 10.6151
R21055 vdd.n1383 vdd.n1381 10.6151
R21056 vdd.n1384 vdd.n1383 10.6151
R21057 vdd.n1386 vdd.n1384 10.6151
R21058 vdd.n1387 vdd.n1386 10.6151
R21059 vdd.n1389 vdd.n1387 10.6151
R21060 vdd.n1390 vdd.n1389 10.6151
R21061 vdd.n1392 vdd.n1390 10.6151
R21062 vdd.n1393 vdd.n1392 10.6151
R21063 vdd.n1395 vdd.n1393 10.6151
R21064 vdd.n1396 vdd.n1395 10.6151
R21065 vdd.n1435 vdd.n1396 10.6151
R21066 vdd.n1435 vdd.n1434 10.6151
R21067 vdd.n1434 vdd.n1433 10.6151
R21068 vdd.n1433 vdd.n1431 10.6151
R21069 vdd.n1431 vdd.n1430 10.6151
R21070 vdd.n1430 vdd.n1428 10.6151
R21071 vdd.n1428 vdd.n1427 10.6151
R21072 vdd.n1427 vdd.n1408 10.6151
R21073 vdd.n1408 vdd.n1407 10.6151
R21074 vdd.n1407 vdd.n1405 10.6151
R21075 vdd.n1405 vdd.n1404 10.6151
R21076 vdd.n1404 vdd.n1402 10.6151
R21077 vdd.n1402 vdd.n1401 10.6151
R21078 vdd.n1401 vdd.n1398 10.6151
R21079 vdd.n1398 vdd.n1397 10.6151
R21080 vdd.n1397 vdd.n1003 10.6151
R21081 vdd.n2509 vdd.n1139 10.6151
R21082 vdd.n2504 vdd.n1139 10.6151
R21083 vdd.n2504 vdd.n2503 10.6151
R21084 vdd.n2503 vdd.n2502 10.6151
R21085 vdd.n2502 vdd.n2499 10.6151
R21086 vdd.n2499 vdd.n2498 10.6151
R21087 vdd.n2498 vdd.n2495 10.6151
R21088 vdd.n2495 vdd.n2494 10.6151
R21089 vdd.n2494 vdd.n2491 10.6151
R21090 vdd.n2491 vdd.n2490 10.6151
R21091 vdd.n2490 vdd.n2487 10.6151
R21092 vdd.n2487 vdd.n2486 10.6151
R21093 vdd.n2486 vdd.n2483 10.6151
R21094 vdd.n2483 vdd.n2482 10.6151
R21095 vdd.n2482 vdd.n2479 10.6151
R21096 vdd.n2479 vdd.n2478 10.6151
R21097 vdd.n2478 vdd.n2475 10.6151
R21098 vdd.n2475 vdd.n1177 10.6151
R21099 vdd.n1323 vdd.n1177 10.6151
R21100 vdd.n1324 vdd.n1323 10.6151
R21101 vdd.n1327 vdd.n1324 10.6151
R21102 vdd.n1328 vdd.n1327 10.6151
R21103 vdd.n1331 vdd.n1328 10.6151
R21104 vdd.n1332 vdd.n1331 10.6151
R21105 vdd.n1335 vdd.n1332 10.6151
R21106 vdd.n1336 vdd.n1335 10.6151
R21107 vdd.n1339 vdd.n1336 10.6151
R21108 vdd.n1340 vdd.n1339 10.6151
R21109 vdd.n1343 vdd.n1340 10.6151
R21110 vdd.n1344 vdd.n1343 10.6151
R21111 vdd.n1347 vdd.n1344 10.6151
R21112 vdd.n1352 vdd.n1349 10.6151
R21113 vdd.n1353 vdd.n1352 10.6151
R21114 vdd.n3020 vdd.n3019 10.6151
R21115 vdd.n3019 vdd.n3018 10.6151
R21116 vdd.n3018 vdd.n2822 10.6151
R21117 vdd.n2900 vdd.n2822 10.6151
R21118 vdd.n2901 vdd.n2900 10.6151
R21119 vdd.n2903 vdd.n2901 10.6151
R21120 vdd.n2904 vdd.n2903 10.6151
R21121 vdd.n3002 vdd.n2904 10.6151
R21122 vdd.n3002 vdd.n3001 10.6151
R21123 vdd.n3001 vdd.n3000 10.6151
R21124 vdd.n3000 vdd.n2948 10.6151
R21125 vdd.n2948 vdd.n2947 10.6151
R21126 vdd.n2947 vdd.n2945 10.6151
R21127 vdd.n2945 vdd.n2944 10.6151
R21128 vdd.n2944 vdd.n2942 10.6151
R21129 vdd.n2942 vdd.n2941 10.6151
R21130 vdd.n2941 vdd.n2939 10.6151
R21131 vdd.n2939 vdd.n2938 10.6151
R21132 vdd.n2938 vdd.n2936 10.6151
R21133 vdd.n2936 vdd.n2935 10.6151
R21134 vdd.n2935 vdd.n2933 10.6151
R21135 vdd.n2933 vdd.n2932 10.6151
R21136 vdd.n2932 vdd.n2930 10.6151
R21137 vdd.n2930 vdd.n2929 10.6151
R21138 vdd.n2929 vdd.n2927 10.6151
R21139 vdd.n2927 vdd.n2926 10.6151
R21140 vdd.n2926 vdd.n2924 10.6151
R21141 vdd.n2924 vdd.n2923 10.6151
R21142 vdd.n2923 vdd.n2921 10.6151
R21143 vdd.n2921 vdd.n2920 10.6151
R21144 vdd.n2920 vdd.n2918 10.6151
R21145 vdd.n2918 vdd.n2917 10.6151
R21146 vdd.n2917 vdd.n2915 10.6151
R21147 vdd.n2915 vdd.n2914 10.6151
R21148 vdd.n2914 vdd.n2912 10.6151
R21149 vdd.n2912 vdd.n2911 10.6151
R21150 vdd.n2911 vdd.n2909 10.6151
R21151 vdd.n2909 vdd.n2908 10.6151
R21152 vdd.n2908 vdd.n2906 10.6151
R21153 vdd.n2906 vdd.n2905 10.6151
R21154 vdd.n2905 vdd.n836 10.6151
R21155 vdd.n3264 vdd.n836 10.6151
R21156 vdd.n3265 vdd.n3264 10.6151
R21157 vdd.n3091 vdd.n961 10.6151
R21158 vdd.n3086 vdd.n961 10.6151
R21159 vdd.n3086 vdd.n3085 10.6151
R21160 vdd.n3085 vdd.n3084 10.6151
R21161 vdd.n3084 vdd.n3081 10.6151
R21162 vdd.n3081 vdd.n3080 10.6151
R21163 vdd.n3080 vdd.n3077 10.6151
R21164 vdd.n3077 vdd.n3076 10.6151
R21165 vdd.n3076 vdd.n3073 10.6151
R21166 vdd.n3073 vdd.n3072 10.6151
R21167 vdd.n3072 vdd.n3069 10.6151
R21168 vdd.n3069 vdd.n3068 10.6151
R21169 vdd.n3068 vdd.n3065 10.6151
R21170 vdd.n3065 vdd.n3064 10.6151
R21171 vdd.n3064 vdd.n3061 10.6151
R21172 vdd.n3061 vdd.n3060 10.6151
R21173 vdd.n3060 vdd.n3057 10.6151
R21174 vdd.n3057 vdd.n3056 10.6151
R21175 vdd.n3056 vdd.n3053 10.6151
R21176 vdd.n3053 vdd.n3052 10.6151
R21177 vdd.n3052 vdd.n3049 10.6151
R21178 vdd.n3049 vdd.n3048 10.6151
R21179 vdd.n3048 vdd.n3045 10.6151
R21180 vdd.n3045 vdd.n3044 10.6151
R21181 vdd.n3044 vdd.n3041 10.6151
R21182 vdd.n3041 vdd.n3040 10.6151
R21183 vdd.n3040 vdd.n3037 10.6151
R21184 vdd.n3037 vdd.n3036 10.6151
R21185 vdd.n3036 vdd.n3033 10.6151
R21186 vdd.n3033 vdd.n3032 10.6151
R21187 vdd.n3032 vdd.n3029 10.6151
R21188 vdd.n3027 vdd.n3024 10.6151
R21189 vdd.n3024 vdd.n3023 10.6151
R21190 vdd.n3093 vdd.n3092 10.6151
R21191 vdd.n3093 vdd.n950 10.6151
R21192 vdd.n3103 vdd.n950 10.6151
R21193 vdd.n3104 vdd.n3103 10.6151
R21194 vdd.n3105 vdd.n3104 10.6151
R21195 vdd.n3105 vdd.n938 10.6151
R21196 vdd.n3115 vdd.n938 10.6151
R21197 vdd.n3116 vdd.n3115 10.6151
R21198 vdd.n3117 vdd.n3116 10.6151
R21199 vdd.n3117 vdd.n927 10.6151
R21200 vdd.n3127 vdd.n927 10.6151
R21201 vdd.n3128 vdd.n3127 10.6151
R21202 vdd.n3129 vdd.n3128 10.6151
R21203 vdd.n3129 vdd.n916 10.6151
R21204 vdd.n3139 vdd.n916 10.6151
R21205 vdd.n3140 vdd.n3139 10.6151
R21206 vdd.n3141 vdd.n3140 10.6151
R21207 vdd.n3141 vdd.n903 10.6151
R21208 vdd.n3152 vdd.n903 10.6151
R21209 vdd.n3153 vdd.n3152 10.6151
R21210 vdd.n3154 vdd.n3153 10.6151
R21211 vdd.n3154 vdd.n891 10.6151
R21212 vdd.n3164 vdd.n891 10.6151
R21213 vdd.n3165 vdd.n3164 10.6151
R21214 vdd.n3166 vdd.n3165 10.6151
R21215 vdd.n3166 vdd.n879 10.6151
R21216 vdd.n3176 vdd.n879 10.6151
R21217 vdd.n3177 vdd.n3176 10.6151
R21218 vdd.n3178 vdd.n3177 10.6151
R21219 vdd.n3178 vdd.n866 10.6151
R21220 vdd.n3188 vdd.n866 10.6151
R21221 vdd.n3189 vdd.n3188 10.6151
R21222 vdd.n3190 vdd.n3189 10.6151
R21223 vdd.n3190 vdd.n855 10.6151
R21224 vdd.n3200 vdd.n855 10.6151
R21225 vdd.n3201 vdd.n3200 10.6151
R21226 vdd.n3202 vdd.n3201 10.6151
R21227 vdd.n3202 vdd.n841 10.6151
R21228 vdd.n3257 vdd.n841 10.6151
R21229 vdd.n3258 vdd.n3257 10.6151
R21230 vdd.n3259 vdd.n3258 10.6151
R21231 vdd.n3259 vdd.n810 10.6151
R21232 vdd.n3329 vdd.n810 10.6151
R21233 vdd.n3328 vdd.n3327 10.6151
R21234 vdd.n3327 vdd.n811 10.6151
R21235 vdd.n812 vdd.n811 10.6151
R21236 vdd.n3320 vdd.n812 10.6151
R21237 vdd.n3320 vdd.n3319 10.6151
R21238 vdd.n3319 vdd.n3318 10.6151
R21239 vdd.n3318 vdd.n814 10.6151
R21240 vdd.n3313 vdd.n814 10.6151
R21241 vdd.n3313 vdd.n3312 10.6151
R21242 vdd.n3312 vdd.n3311 10.6151
R21243 vdd.n3311 vdd.n817 10.6151
R21244 vdd.n3306 vdd.n817 10.6151
R21245 vdd.n3306 vdd.n3305 10.6151
R21246 vdd.n3305 vdd.n3304 10.6151
R21247 vdd.n3304 vdd.n820 10.6151
R21248 vdd.n3299 vdd.n820 10.6151
R21249 vdd.n3299 vdd.n731 10.6151
R21250 vdd.n3295 vdd.n731 10.6151
R21251 vdd.n3295 vdd.n3294 10.6151
R21252 vdd.n3294 vdd.n3293 10.6151
R21253 vdd.n3293 vdd.n823 10.6151
R21254 vdd.n3288 vdd.n823 10.6151
R21255 vdd.n3288 vdd.n3287 10.6151
R21256 vdd.n3287 vdd.n3286 10.6151
R21257 vdd.n3286 vdd.n826 10.6151
R21258 vdd.n3281 vdd.n826 10.6151
R21259 vdd.n3281 vdd.n3280 10.6151
R21260 vdd.n3280 vdd.n3279 10.6151
R21261 vdd.n3279 vdd.n829 10.6151
R21262 vdd.n3274 vdd.n829 10.6151
R21263 vdd.n3274 vdd.n3273 10.6151
R21264 vdd.n3271 vdd.n834 10.6151
R21265 vdd.n3266 vdd.n834 10.6151
R21266 vdd.n3247 vdd.n3208 10.6151
R21267 vdd.n3242 vdd.n3208 10.6151
R21268 vdd.n3242 vdd.n3241 10.6151
R21269 vdd.n3241 vdd.n3240 10.6151
R21270 vdd.n3240 vdd.n3210 10.6151
R21271 vdd.n3235 vdd.n3210 10.6151
R21272 vdd.n3235 vdd.n3234 10.6151
R21273 vdd.n3234 vdd.n3233 10.6151
R21274 vdd.n3233 vdd.n3213 10.6151
R21275 vdd.n3228 vdd.n3213 10.6151
R21276 vdd.n3228 vdd.n3227 10.6151
R21277 vdd.n3227 vdd.n3226 10.6151
R21278 vdd.n3226 vdd.n3216 10.6151
R21279 vdd.n3221 vdd.n3216 10.6151
R21280 vdd.n3221 vdd.n3220 10.6151
R21281 vdd.n3220 vdd.n785 10.6151
R21282 vdd.n3364 vdd.n785 10.6151
R21283 vdd.n3364 vdd.n786 10.6151
R21284 vdd.n788 vdd.n786 10.6151
R21285 vdd.n3357 vdd.n788 10.6151
R21286 vdd.n3357 vdd.n3356 10.6151
R21287 vdd.n3356 vdd.n3355 10.6151
R21288 vdd.n3355 vdd.n790 10.6151
R21289 vdd.n3350 vdd.n790 10.6151
R21290 vdd.n3350 vdd.n3349 10.6151
R21291 vdd.n3349 vdd.n3348 10.6151
R21292 vdd.n3348 vdd.n793 10.6151
R21293 vdd.n3343 vdd.n793 10.6151
R21294 vdd.n3343 vdd.n3342 10.6151
R21295 vdd.n3342 vdd.n3341 10.6151
R21296 vdd.n3341 vdd.n796 10.6151
R21297 vdd.n3336 vdd.n3335 10.6151
R21298 vdd.n3335 vdd.n3334 10.6151
R21299 vdd.n2897 vdd.n2896 10.6151
R21300 vdd.n3014 vdd.n2897 10.6151
R21301 vdd.n3014 vdd.n3013 10.6151
R21302 vdd.n3013 vdd.n3012 10.6151
R21303 vdd.n3012 vdd.n3010 10.6151
R21304 vdd.n3010 vdd.n3009 10.6151
R21305 vdd.n3009 vdd.n3007 10.6151
R21306 vdd.n3007 vdd.n3006 10.6151
R21307 vdd.n3006 vdd.n2898 10.6151
R21308 vdd.n2996 vdd.n2898 10.6151
R21309 vdd.n2996 vdd.n2995 10.6151
R21310 vdd.n2995 vdd.n2994 10.6151
R21311 vdd.n2994 vdd.n2992 10.6151
R21312 vdd.n2992 vdd.n2991 10.6151
R21313 vdd.n2991 vdd.n2989 10.6151
R21314 vdd.n2989 vdd.n2988 10.6151
R21315 vdd.n2988 vdd.n2986 10.6151
R21316 vdd.n2986 vdd.n2985 10.6151
R21317 vdd.n2985 vdd.n2983 10.6151
R21318 vdd.n2983 vdd.n2982 10.6151
R21319 vdd.n2982 vdd.n2980 10.6151
R21320 vdd.n2980 vdd.n2979 10.6151
R21321 vdd.n2979 vdd.n2977 10.6151
R21322 vdd.n2977 vdd.n2976 10.6151
R21323 vdd.n2976 vdd.n2974 10.6151
R21324 vdd.n2974 vdd.n2973 10.6151
R21325 vdd.n2973 vdd.n2971 10.6151
R21326 vdd.n2971 vdd.n2970 10.6151
R21327 vdd.n2970 vdd.n2968 10.6151
R21328 vdd.n2968 vdd.n2967 10.6151
R21329 vdd.n2967 vdd.n2965 10.6151
R21330 vdd.n2965 vdd.n2964 10.6151
R21331 vdd.n2964 vdd.n2962 10.6151
R21332 vdd.n2962 vdd.n2961 10.6151
R21333 vdd.n2961 vdd.n2959 10.6151
R21334 vdd.n2959 vdd.n2958 10.6151
R21335 vdd.n2958 vdd.n2956 10.6151
R21336 vdd.n2956 vdd.n2955 10.6151
R21337 vdd.n2955 vdd.n2953 10.6151
R21338 vdd.n2953 vdd.n2952 10.6151
R21339 vdd.n2952 vdd.n2950 10.6151
R21340 vdd.n2950 vdd.n2949 10.6151
R21341 vdd.n2949 vdd.n802 10.6151
R21342 vdd.n2828 vdd.n2827 10.6151
R21343 vdd.n2831 vdd.n2828 10.6151
R21344 vdd.n2832 vdd.n2831 10.6151
R21345 vdd.n2835 vdd.n2832 10.6151
R21346 vdd.n2836 vdd.n2835 10.6151
R21347 vdd.n2839 vdd.n2836 10.6151
R21348 vdd.n2840 vdd.n2839 10.6151
R21349 vdd.n2843 vdd.n2840 10.6151
R21350 vdd.n2844 vdd.n2843 10.6151
R21351 vdd.n2847 vdd.n2844 10.6151
R21352 vdd.n2848 vdd.n2847 10.6151
R21353 vdd.n2851 vdd.n2848 10.6151
R21354 vdd.n2852 vdd.n2851 10.6151
R21355 vdd.n2855 vdd.n2852 10.6151
R21356 vdd.n2856 vdd.n2855 10.6151
R21357 vdd.n2859 vdd.n2856 10.6151
R21358 vdd.n2860 vdd.n2859 10.6151
R21359 vdd.n2863 vdd.n2860 10.6151
R21360 vdd.n2864 vdd.n2863 10.6151
R21361 vdd.n2867 vdd.n2864 10.6151
R21362 vdd.n2868 vdd.n2867 10.6151
R21363 vdd.n2871 vdd.n2868 10.6151
R21364 vdd.n2872 vdd.n2871 10.6151
R21365 vdd.n2875 vdd.n2872 10.6151
R21366 vdd.n2876 vdd.n2875 10.6151
R21367 vdd.n2879 vdd.n2876 10.6151
R21368 vdd.n2880 vdd.n2879 10.6151
R21369 vdd.n2883 vdd.n2880 10.6151
R21370 vdd.n2884 vdd.n2883 10.6151
R21371 vdd.n2887 vdd.n2884 10.6151
R21372 vdd.n2888 vdd.n2887 10.6151
R21373 vdd.n2893 vdd.n2891 10.6151
R21374 vdd.n2894 vdd.n2893 10.6151
R21375 vdd.n3097 vdd.n955 10.6151
R21376 vdd.n3098 vdd.n3097 10.6151
R21377 vdd.n3099 vdd.n3098 10.6151
R21378 vdd.n3099 vdd.n944 10.6151
R21379 vdd.n3109 vdd.n944 10.6151
R21380 vdd.n3110 vdd.n3109 10.6151
R21381 vdd.n3111 vdd.n3110 10.6151
R21382 vdd.n3111 vdd.n933 10.6151
R21383 vdd.n3121 vdd.n933 10.6151
R21384 vdd.n3122 vdd.n3121 10.6151
R21385 vdd.n3123 vdd.n3122 10.6151
R21386 vdd.n3123 vdd.n921 10.6151
R21387 vdd.n3133 vdd.n921 10.6151
R21388 vdd.n3134 vdd.n3133 10.6151
R21389 vdd.n3135 vdd.n3134 10.6151
R21390 vdd.n3135 vdd.n910 10.6151
R21391 vdd.n3145 vdd.n910 10.6151
R21392 vdd.n3146 vdd.n3145 10.6151
R21393 vdd.n3148 vdd.n3146 10.6151
R21394 vdd.n3148 vdd.n3147 10.6151
R21395 vdd.n3159 vdd.n3158 10.6151
R21396 vdd.n3160 vdd.n3159 10.6151
R21397 vdd.n3160 vdd.n885 10.6151
R21398 vdd.n3170 vdd.n885 10.6151
R21399 vdd.n3171 vdd.n3170 10.6151
R21400 vdd.n3172 vdd.n3171 10.6151
R21401 vdd.n3172 vdd.n872 10.6151
R21402 vdd.n3182 vdd.n872 10.6151
R21403 vdd.n3183 vdd.n3182 10.6151
R21404 vdd.n3184 vdd.n3183 10.6151
R21405 vdd.n3184 vdd.n860 10.6151
R21406 vdd.n3194 vdd.n860 10.6151
R21407 vdd.n3195 vdd.n3194 10.6151
R21408 vdd.n3196 vdd.n3195 10.6151
R21409 vdd.n3196 vdd.n849 10.6151
R21410 vdd.n3206 vdd.n849 10.6151
R21411 vdd.n3207 vdd.n3206 10.6151
R21412 vdd.n3253 vdd.n3207 10.6151
R21413 vdd.n3253 vdd.n3252 10.6151
R21414 vdd.n3252 vdd.n3251 10.6151
R21415 vdd.n3251 vdd.n3250 10.6151
R21416 vdd.n3250 vdd.n3248 10.6151
R21417 vdd.n2515 vdd.n1132 10.6151
R21418 vdd.n2516 vdd.n2515 10.6151
R21419 vdd.n2517 vdd.n2516 10.6151
R21420 vdd.n2517 vdd.n1121 10.6151
R21421 vdd.n2527 vdd.n1121 10.6151
R21422 vdd.n2528 vdd.n2527 10.6151
R21423 vdd.n2529 vdd.n2528 10.6151
R21424 vdd.n2529 vdd.n1108 10.6151
R21425 vdd.n2539 vdd.n1108 10.6151
R21426 vdd.n2540 vdd.n2539 10.6151
R21427 vdd.n2541 vdd.n2540 10.6151
R21428 vdd.n2541 vdd.n1097 10.6151
R21429 vdd.n2551 vdd.n1097 10.6151
R21430 vdd.n2552 vdd.n2551 10.6151
R21431 vdd.n2553 vdd.n2552 10.6151
R21432 vdd.n2553 vdd.n1085 10.6151
R21433 vdd.n2563 vdd.n1085 10.6151
R21434 vdd.n2564 vdd.n2563 10.6151
R21435 vdd.n2565 vdd.n2564 10.6151
R21436 vdd.n2565 vdd.n1072 10.6151
R21437 vdd.n2575 vdd.n1072 10.6151
R21438 vdd.n2576 vdd.n2575 10.6151
R21439 vdd.n2578 vdd.n1060 10.6151
R21440 vdd.n2588 vdd.n1060 10.6151
R21441 vdd.n2589 vdd.n2588 10.6151
R21442 vdd.n2590 vdd.n2589 10.6151
R21443 vdd.n2590 vdd.n1048 10.6151
R21444 vdd.n2600 vdd.n1048 10.6151
R21445 vdd.n2601 vdd.n2600 10.6151
R21446 vdd.n2602 vdd.n2601 10.6151
R21447 vdd.n2602 vdd.n1037 10.6151
R21448 vdd.n2612 vdd.n1037 10.6151
R21449 vdd.n2613 vdd.n2612 10.6151
R21450 vdd.n2614 vdd.n2613 10.6151
R21451 vdd.n2614 vdd.n1026 10.6151
R21452 vdd.n2624 vdd.n1026 10.6151
R21453 vdd.n2625 vdd.n2624 10.6151
R21454 vdd.n2628 vdd.n2625 10.6151
R21455 vdd.n2628 vdd.n2627 10.6151
R21456 vdd.n2627 vdd.n2626 10.6151
R21457 vdd.n2626 vdd.n1009 10.6151
R21458 vdd.n2710 vdd.n1009 10.6151
R21459 vdd.n2709 vdd.n2708 10.6151
R21460 vdd.n2708 vdd.n2705 10.6151
R21461 vdd.n2705 vdd.n2704 10.6151
R21462 vdd.n2704 vdd.n2701 10.6151
R21463 vdd.n2701 vdd.n2700 10.6151
R21464 vdd.n2700 vdd.n2697 10.6151
R21465 vdd.n2697 vdd.n2696 10.6151
R21466 vdd.n2696 vdd.n2693 10.6151
R21467 vdd.n2693 vdd.n2692 10.6151
R21468 vdd.n2692 vdd.n2689 10.6151
R21469 vdd.n2689 vdd.n2688 10.6151
R21470 vdd.n2688 vdd.n2685 10.6151
R21471 vdd.n2685 vdd.n2684 10.6151
R21472 vdd.n2684 vdd.n2681 10.6151
R21473 vdd.n2681 vdd.n2680 10.6151
R21474 vdd.n2680 vdd.n2677 10.6151
R21475 vdd.n2677 vdd.n2676 10.6151
R21476 vdd.n2676 vdd.n2673 10.6151
R21477 vdd.n2673 vdd.n2672 10.6151
R21478 vdd.n2672 vdd.n2669 10.6151
R21479 vdd.n2669 vdd.n2668 10.6151
R21480 vdd.n2668 vdd.n2665 10.6151
R21481 vdd.n2665 vdd.n2664 10.6151
R21482 vdd.n2664 vdd.n2661 10.6151
R21483 vdd.n2661 vdd.n2660 10.6151
R21484 vdd.n2660 vdd.n2657 10.6151
R21485 vdd.n2657 vdd.n2656 10.6151
R21486 vdd.n2656 vdd.n2653 10.6151
R21487 vdd.n2653 vdd.n2652 10.6151
R21488 vdd.n2652 vdd.n2649 10.6151
R21489 vdd.n2649 vdd.n2648 10.6151
R21490 vdd.n2645 vdd.n2644 10.6151
R21491 vdd.n2644 vdd.n2642 10.6151
R21492 vdd.n1481 vdd.n1479 10.6151
R21493 vdd.n1479 vdd.n1478 10.6151
R21494 vdd.n1478 vdd.n1476 10.6151
R21495 vdd.n1476 vdd.n1475 10.6151
R21496 vdd.n1475 vdd.n1473 10.6151
R21497 vdd.n1473 vdd.n1472 10.6151
R21498 vdd.n1472 vdd.n1470 10.6151
R21499 vdd.n1470 vdd.n1469 10.6151
R21500 vdd.n1469 vdd.n1467 10.6151
R21501 vdd.n1467 vdd.n1466 10.6151
R21502 vdd.n1466 vdd.n1464 10.6151
R21503 vdd.n1464 vdd.n1463 10.6151
R21504 vdd.n1463 vdd.n1461 10.6151
R21505 vdd.n1461 vdd.n1460 10.6151
R21506 vdd.n1460 vdd.n1458 10.6151
R21507 vdd.n1458 vdd.n1457 10.6151
R21508 vdd.n1457 vdd.n1455 10.6151
R21509 vdd.n1455 vdd.n1454 10.6151
R21510 vdd.n1454 vdd.n1452 10.6151
R21511 vdd.n1452 vdd.n1451 10.6151
R21512 vdd.n1451 vdd.n1449 10.6151
R21513 vdd.n1449 vdd.n1448 10.6151
R21514 vdd.n1448 vdd.n1446 10.6151
R21515 vdd.n1446 vdd.n1445 10.6151
R21516 vdd.n1445 vdd.n1443 10.6151
R21517 vdd.n1443 vdd.n1442 10.6151
R21518 vdd.n1442 vdd.n1440 10.6151
R21519 vdd.n1440 vdd.n1439 10.6151
R21520 vdd.n1439 vdd.n1318 10.6151
R21521 vdd.n1410 vdd.n1318 10.6151
R21522 vdd.n1411 vdd.n1410 10.6151
R21523 vdd.n1413 vdd.n1411 10.6151
R21524 vdd.n1414 vdd.n1413 10.6151
R21525 vdd.n1423 vdd.n1414 10.6151
R21526 vdd.n1423 vdd.n1422 10.6151
R21527 vdd.n1422 vdd.n1421 10.6151
R21528 vdd.n1421 vdd.n1419 10.6151
R21529 vdd.n1419 vdd.n1418 10.6151
R21530 vdd.n1418 vdd.n1416 10.6151
R21531 vdd.n1416 vdd.n1415 10.6151
R21532 vdd.n1415 vdd.n1013 10.6151
R21533 vdd.n2640 vdd.n1013 10.6151
R21534 vdd.n2641 vdd.n2640 10.6151
R21535 vdd.n1282 vdd.n1281 10.6151
R21536 vdd.n1285 vdd.n1282 10.6151
R21537 vdd.n1286 vdd.n1285 10.6151
R21538 vdd.n1289 vdd.n1286 10.6151
R21539 vdd.n1290 vdd.n1289 10.6151
R21540 vdd.n1293 vdd.n1290 10.6151
R21541 vdd.n1294 vdd.n1293 10.6151
R21542 vdd.n1297 vdd.n1294 10.6151
R21543 vdd.n1298 vdd.n1297 10.6151
R21544 vdd.n1301 vdd.n1298 10.6151
R21545 vdd.n1302 vdd.n1301 10.6151
R21546 vdd.n1305 vdd.n1302 10.6151
R21547 vdd.n1306 vdd.n1305 10.6151
R21548 vdd.n1309 vdd.n1306 10.6151
R21549 vdd.n1310 vdd.n1309 10.6151
R21550 vdd.n1313 vdd.n1310 10.6151
R21551 vdd.n1515 vdd.n1313 10.6151
R21552 vdd.n1515 vdd.n1514 10.6151
R21553 vdd.n1514 vdd.n1512 10.6151
R21554 vdd.n1512 vdd.n1509 10.6151
R21555 vdd.n1509 vdd.n1508 10.6151
R21556 vdd.n1508 vdd.n1505 10.6151
R21557 vdd.n1505 vdd.n1504 10.6151
R21558 vdd.n1504 vdd.n1501 10.6151
R21559 vdd.n1501 vdd.n1500 10.6151
R21560 vdd.n1500 vdd.n1497 10.6151
R21561 vdd.n1497 vdd.n1496 10.6151
R21562 vdd.n1496 vdd.n1493 10.6151
R21563 vdd.n1493 vdd.n1492 10.6151
R21564 vdd.n1492 vdd.n1489 10.6151
R21565 vdd.n1489 vdd.n1488 10.6151
R21566 vdd.n1485 vdd.n1484 10.6151
R21567 vdd.n1484 vdd.n1482 10.6151
R21568 vdd.n2306 vdd.t39 10.5435
R21569 vdd.n656 vdd.t16 10.5435
R21570 vdd.n316 vdd.n298 10.4732
R21571 vdd.n257 vdd.n239 10.4732
R21572 vdd.n214 vdd.n196 10.4732
R21573 vdd.n155 vdd.n137 10.4732
R21574 vdd.n113 vdd.n95 10.4732
R21575 vdd.n54 vdd.n36 10.4732
R21576 vdd.n2190 vdd.n2172 10.4732
R21577 vdd.n2249 vdd.n2231 10.4732
R21578 vdd.n2088 vdd.n2070 10.4732
R21579 vdd.n2147 vdd.n2129 10.4732
R21580 vdd.n1987 vdd.n1969 10.4732
R21581 vdd.n2046 vdd.n2028 10.4732
R21582 vdd.t60 vdd.n2280 10.3167
R21583 vdd.n3572 vdd.t6 10.3167
R21584 vdd.n1957 vdd.t52 10.09
R21585 vdd.n3666 vdd.t18 10.09
R21586 vdd.n2475 vdd.n2474 9.98956
R21587 vdd.n3488 vdd.n731 9.98956
R21588 vdd.n3365 vdd.n3364 9.98956
R21589 vdd.n2367 vdd.n1515 9.98956
R21590 vdd.t44 vdd.n1610 9.86327
R21591 vdd.n3657 vdd.t139 9.86327
R21592 vdd.n2712 vdd.t286 9.7499
R21593 vdd.t269 vdd.n957 9.7499
R21594 vdd.n315 vdd.n300 9.69747
R21595 vdd.n256 vdd.n241 9.69747
R21596 vdd.n213 vdd.n198 9.69747
R21597 vdd.n154 vdd.n139 9.69747
R21598 vdd.n112 vdd.n97 9.69747
R21599 vdd.n53 vdd.n38 9.69747
R21600 vdd.n2189 vdd.n2174 9.69747
R21601 vdd.n2248 vdd.n2233 9.69747
R21602 vdd.n2087 vdd.n2072 9.69747
R21603 vdd.n2146 vdd.n2131 9.69747
R21604 vdd.n1986 vdd.n1971 9.69747
R21605 vdd.n2045 vdd.n2030 9.69747
R21606 vdd.n1916 vdd.t32 9.63654
R21607 vdd.n3603 vdd.t66 9.63654
R21608 vdd.n331 vdd.n330 9.45567
R21609 vdd.n272 vdd.n271 9.45567
R21610 vdd.n229 vdd.n228 9.45567
R21611 vdd.n170 vdd.n169 9.45567
R21612 vdd.n128 vdd.n127 9.45567
R21613 vdd.n69 vdd.n68 9.45567
R21614 vdd.n2205 vdd.n2204 9.45567
R21615 vdd.n2264 vdd.n2263 9.45567
R21616 vdd.n2103 vdd.n2102 9.45567
R21617 vdd.n2162 vdd.n2161 9.45567
R21618 vdd.n2002 vdd.n2001 9.45567
R21619 vdd.n2061 vdd.n2060 9.45567
R21620 vdd.n1890 vdd.t87 9.40981
R21621 vdd.n3635 vdd.t14 9.40981
R21622 vdd.n2437 vdd.n1207 9.3005
R21623 vdd.n2436 vdd.n2435 9.3005
R21624 vdd.n1213 vdd.n1212 9.3005
R21625 vdd.n2430 vdd.n1217 9.3005
R21626 vdd.n2429 vdd.n1218 9.3005
R21627 vdd.n2428 vdd.n1219 9.3005
R21628 vdd.n1223 vdd.n1220 9.3005
R21629 vdd.n2423 vdd.n1224 9.3005
R21630 vdd.n2422 vdd.n1225 9.3005
R21631 vdd.n2421 vdd.n1226 9.3005
R21632 vdd.n1230 vdd.n1227 9.3005
R21633 vdd.n2416 vdd.n1231 9.3005
R21634 vdd.n2415 vdd.n1232 9.3005
R21635 vdd.n2414 vdd.n1233 9.3005
R21636 vdd.n1237 vdd.n1234 9.3005
R21637 vdd.n2409 vdd.n1238 9.3005
R21638 vdd.n2408 vdd.n1239 9.3005
R21639 vdd.n2407 vdd.n1240 9.3005
R21640 vdd.n1244 vdd.n1241 9.3005
R21641 vdd.n2402 vdd.n1245 9.3005
R21642 vdd.n2401 vdd.n1246 9.3005
R21643 vdd.n2400 vdd.n2399 9.3005
R21644 vdd.n2398 vdd.n1247 9.3005
R21645 vdd.n2397 vdd.n2396 9.3005
R21646 vdd.n1253 vdd.n1252 9.3005
R21647 vdd.n2391 vdd.n1257 9.3005
R21648 vdd.n2390 vdd.n1258 9.3005
R21649 vdd.n2389 vdd.n1259 9.3005
R21650 vdd.n1263 vdd.n1260 9.3005
R21651 vdd.n2384 vdd.n1264 9.3005
R21652 vdd.n2383 vdd.n1265 9.3005
R21653 vdd.n2382 vdd.n1266 9.3005
R21654 vdd.n1270 vdd.n1267 9.3005
R21655 vdd.n2377 vdd.n1271 9.3005
R21656 vdd.n2376 vdd.n1272 9.3005
R21657 vdd.n2375 vdd.n1273 9.3005
R21658 vdd.n1277 vdd.n1274 9.3005
R21659 vdd.n2370 vdd.n1278 9.3005
R21660 vdd.n2439 vdd.n2438 9.3005
R21661 vdd.n2461 vdd.n1178 9.3005
R21662 vdd.n2460 vdd.n1186 9.3005
R21663 vdd.n1190 vdd.n1187 9.3005
R21664 vdd.n2455 vdd.n1191 9.3005
R21665 vdd.n2454 vdd.n1192 9.3005
R21666 vdd.n2453 vdd.n1193 9.3005
R21667 vdd.n1197 vdd.n1194 9.3005
R21668 vdd.n2448 vdd.n1198 9.3005
R21669 vdd.n2447 vdd.n1199 9.3005
R21670 vdd.n2446 vdd.n1200 9.3005
R21671 vdd.n1204 vdd.n1201 9.3005
R21672 vdd.n2441 vdd.n1205 9.3005
R21673 vdd.n2440 vdd.n1206 9.3005
R21674 vdd.n2473 vdd.n2472 9.3005
R21675 vdd.n1182 vdd.n1181 9.3005
R21676 vdd.n2270 vdd.n2269 9.3005
R21677 vdd.n1579 vdd.n1578 9.3005
R21678 vdd.n2284 vdd.n2283 9.3005
R21679 vdd.n2285 vdd.n1577 9.3005
R21680 vdd.n2287 vdd.n2286 9.3005
R21681 vdd.n1568 vdd.n1567 9.3005
R21682 vdd.n2301 vdd.n2300 9.3005
R21683 vdd.n2302 vdd.n1566 9.3005
R21684 vdd.n2304 vdd.n2303 9.3005
R21685 vdd.n1557 vdd.n1556 9.3005
R21686 vdd.n2317 vdd.n2316 9.3005
R21687 vdd.n2318 vdd.n1555 9.3005
R21688 vdd.n2320 vdd.n2319 9.3005
R21689 vdd.n1545 vdd.n1544 9.3005
R21690 vdd.n2334 vdd.n2333 9.3005
R21691 vdd.n2335 vdd.n1543 9.3005
R21692 vdd.n2337 vdd.n2336 9.3005
R21693 vdd.n1533 vdd.n1532 9.3005
R21694 vdd.n2353 vdd.n2352 9.3005
R21695 vdd.n2354 vdd.n1531 9.3005
R21696 vdd.n2356 vdd.n2355 9.3005
R21697 vdd.n307 vdd.n306 9.3005
R21698 vdd.n302 vdd.n301 9.3005
R21699 vdd.n313 vdd.n312 9.3005
R21700 vdd.n315 vdd.n314 9.3005
R21701 vdd.n298 vdd.n297 9.3005
R21702 vdd.n321 vdd.n320 9.3005
R21703 vdd.n323 vdd.n322 9.3005
R21704 vdd.n295 vdd.n292 9.3005
R21705 vdd.n330 vdd.n329 9.3005
R21706 vdd.n248 vdd.n247 9.3005
R21707 vdd.n243 vdd.n242 9.3005
R21708 vdd.n254 vdd.n253 9.3005
R21709 vdd.n256 vdd.n255 9.3005
R21710 vdd.n239 vdd.n238 9.3005
R21711 vdd.n262 vdd.n261 9.3005
R21712 vdd.n264 vdd.n263 9.3005
R21713 vdd.n236 vdd.n233 9.3005
R21714 vdd.n271 vdd.n270 9.3005
R21715 vdd.n205 vdd.n204 9.3005
R21716 vdd.n200 vdd.n199 9.3005
R21717 vdd.n211 vdd.n210 9.3005
R21718 vdd.n213 vdd.n212 9.3005
R21719 vdd.n196 vdd.n195 9.3005
R21720 vdd.n219 vdd.n218 9.3005
R21721 vdd.n221 vdd.n220 9.3005
R21722 vdd.n193 vdd.n190 9.3005
R21723 vdd.n228 vdd.n227 9.3005
R21724 vdd.n146 vdd.n145 9.3005
R21725 vdd.n141 vdd.n140 9.3005
R21726 vdd.n152 vdd.n151 9.3005
R21727 vdd.n154 vdd.n153 9.3005
R21728 vdd.n137 vdd.n136 9.3005
R21729 vdd.n160 vdd.n159 9.3005
R21730 vdd.n162 vdd.n161 9.3005
R21731 vdd.n134 vdd.n131 9.3005
R21732 vdd.n169 vdd.n168 9.3005
R21733 vdd.n104 vdd.n103 9.3005
R21734 vdd.n99 vdd.n98 9.3005
R21735 vdd.n110 vdd.n109 9.3005
R21736 vdd.n112 vdd.n111 9.3005
R21737 vdd.n95 vdd.n94 9.3005
R21738 vdd.n118 vdd.n117 9.3005
R21739 vdd.n120 vdd.n119 9.3005
R21740 vdd.n92 vdd.n89 9.3005
R21741 vdd.n127 vdd.n126 9.3005
R21742 vdd.n45 vdd.n44 9.3005
R21743 vdd.n40 vdd.n39 9.3005
R21744 vdd.n51 vdd.n50 9.3005
R21745 vdd.n53 vdd.n52 9.3005
R21746 vdd.n36 vdd.n35 9.3005
R21747 vdd.n59 vdd.n58 9.3005
R21748 vdd.n61 vdd.n60 9.3005
R21749 vdd.n33 vdd.n30 9.3005
R21750 vdd.n68 vdd.n67 9.3005
R21751 vdd.n3410 vdd.n3409 9.3005
R21752 vdd.n3413 vdd.n766 9.3005
R21753 vdd.n3414 vdd.n765 9.3005
R21754 vdd.n3417 vdd.n764 9.3005
R21755 vdd.n3418 vdd.n763 9.3005
R21756 vdd.n3421 vdd.n762 9.3005
R21757 vdd.n3422 vdd.n761 9.3005
R21758 vdd.n3425 vdd.n760 9.3005
R21759 vdd.n3426 vdd.n759 9.3005
R21760 vdd.n3429 vdd.n758 9.3005
R21761 vdd.n3430 vdd.n757 9.3005
R21762 vdd.n3433 vdd.n756 9.3005
R21763 vdd.n3434 vdd.n755 9.3005
R21764 vdd.n3437 vdd.n754 9.3005
R21765 vdd.n3438 vdd.n753 9.3005
R21766 vdd.n3441 vdd.n752 9.3005
R21767 vdd.n3442 vdd.n751 9.3005
R21768 vdd.n3445 vdd.n750 9.3005
R21769 vdd.n3446 vdd.n749 9.3005
R21770 vdd.n3449 vdd.n748 9.3005
R21771 vdd.n3453 vdd.n3452 9.3005
R21772 vdd.n3454 vdd.n747 9.3005
R21773 vdd.n3458 vdd.n3455 9.3005
R21774 vdd.n3461 vdd.n746 9.3005
R21775 vdd.n3462 vdd.n745 9.3005
R21776 vdd.n3465 vdd.n744 9.3005
R21777 vdd.n3466 vdd.n743 9.3005
R21778 vdd.n3469 vdd.n742 9.3005
R21779 vdd.n3470 vdd.n741 9.3005
R21780 vdd.n3473 vdd.n740 9.3005
R21781 vdd.n3474 vdd.n739 9.3005
R21782 vdd.n3477 vdd.n738 9.3005
R21783 vdd.n3478 vdd.n737 9.3005
R21784 vdd.n3481 vdd.n736 9.3005
R21785 vdd.n3482 vdd.n735 9.3005
R21786 vdd.n3485 vdd.n730 9.3005
R21787 vdd.n3491 vdd.n727 9.3005
R21788 vdd.n3492 vdd.n726 9.3005
R21789 vdd.n3506 vdd.n3505 9.3005
R21790 vdd.n3507 vdd.n681 9.3005
R21791 vdd.n3509 vdd.n3508 9.3005
R21792 vdd.n671 vdd.n670 9.3005
R21793 vdd.n3523 vdd.n3522 9.3005
R21794 vdd.n3524 vdd.n669 9.3005
R21795 vdd.n3526 vdd.n3525 9.3005
R21796 vdd.n660 vdd.n659 9.3005
R21797 vdd.n3539 vdd.n3538 9.3005
R21798 vdd.n3540 vdd.n658 9.3005
R21799 vdd.n3542 vdd.n3541 9.3005
R21800 vdd.n648 vdd.n647 9.3005
R21801 vdd.n3556 vdd.n3555 9.3005
R21802 vdd.n3557 vdd.n646 9.3005
R21803 vdd.n3559 vdd.n3558 9.3005
R21804 vdd.n637 vdd.n636 9.3005
R21805 vdd.n3575 vdd.n3574 9.3005
R21806 vdd.n3576 vdd.n635 9.3005
R21807 vdd.n3578 vdd.n3577 9.3005
R21808 vdd.n336 vdd.n334 9.3005
R21809 vdd.n683 vdd.n682 9.3005
R21810 vdd.n3670 vdd.n3669 9.3005
R21811 vdd.n337 vdd.n335 9.3005
R21812 vdd.n3663 vdd.n346 9.3005
R21813 vdd.n3662 vdd.n347 9.3005
R21814 vdd.n3661 vdd.n348 9.3005
R21815 vdd.n355 vdd.n349 9.3005
R21816 vdd.n3655 vdd.n356 9.3005
R21817 vdd.n3654 vdd.n357 9.3005
R21818 vdd.n3653 vdd.n358 9.3005
R21819 vdd.n366 vdd.n359 9.3005
R21820 vdd.n3647 vdd.n367 9.3005
R21821 vdd.n3646 vdd.n368 9.3005
R21822 vdd.n3645 vdd.n369 9.3005
R21823 vdd.n377 vdd.n370 9.3005
R21824 vdd.n3639 vdd.n378 9.3005
R21825 vdd.n3638 vdd.n379 9.3005
R21826 vdd.n3637 vdd.n380 9.3005
R21827 vdd.n388 vdd.n381 9.3005
R21828 vdd.n3631 vdd.n389 9.3005
R21829 vdd.n3630 vdd.n390 9.3005
R21830 vdd.n3629 vdd.n391 9.3005
R21831 vdd.n466 vdd.n463 9.3005
R21832 vdd.n470 vdd.n469 9.3005
R21833 vdd.n471 vdd.n462 9.3005
R21834 vdd.n475 vdd.n472 9.3005
R21835 vdd.n476 vdd.n461 9.3005
R21836 vdd.n480 vdd.n479 9.3005
R21837 vdd.n481 vdd.n460 9.3005
R21838 vdd.n485 vdd.n482 9.3005
R21839 vdd.n486 vdd.n459 9.3005
R21840 vdd.n490 vdd.n489 9.3005
R21841 vdd.n491 vdd.n458 9.3005
R21842 vdd.n495 vdd.n492 9.3005
R21843 vdd.n496 vdd.n457 9.3005
R21844 vdd.n500 vdd.n499 9.3005
R21845 vdd.n501 vdd.n456 9.3005
R21846 vdd.n505 vdd.n502 9.3005
R21847 vdd.n506 vdd.n455 9.3005
R21848 vdd.n510 vdd.n509 9.3005
R21849 vdd.n511 vdd.n454 9.3005
R21850 vdd.n515 vdd.n512 9.3005
R21851 vdd.n516 vdd.n451 9.3005
R21852 vdd.n520 vdd.n519 9.3005
R21853 vdd.n521 vdd.n450 9.3005
R21854 vdd.n525 vdd.n522 9.3005
R21855 vdd.n526 vdd.n449 9.3005
R21856 vdd.n530 vdd.n529 9.3005
R21857 vdd.n531 vdd.n448 9.3005
R21858 vdd.n535 vdd.n532 9.3005
R21859 vdd.n536 vdd.n447 9.3005
R21860 vdd.n540 vdd.n539 9.3005
R21861 vdd.n541 vdd.n446 9.3005
R21862 vdd.n545 vdd.n542 9.3005
R21863 vdd.n546 vdd.n445 9.3005
R21864 vdd.n550 vdd.n549 9.3005
R21865 vdd.n551 vdd.n444 9.3005
R21866 vdd.n555 vdd.n552 9.3005
R21867 vdd.n556 vdd.n443 9.3005
R21868 vdd.n560 vdd.n559 9.3005
R21869 vdd.n561 vdd.n442 9.3005
R21870 vdd.n565 vdd.n562 9.3005
R21871 vdd.n566 vdd.n439 9.3005
R21872 vdd.n570 vdd.n569 9.3005
R21873 vdd.n571 vdd.n438 9.3005
R21874 vdd.n575 vdd.n572 9.3005
R21875 vdd.n576 vdd.n437 9.3005
R21876 vdd.n580 vdd.n579 9.3005
R21877 vdd.n581 vdd.n436 9.3005
R21878 vdd.n585 vdd.n582 9.3005
R21879 vdd.n586 vdd.n435 9.3005
R21880 vdd.n590 vdd.n589 9.3005
R21881 vdd.n591 vdd.n434 9.3005
R21882 vdd.n595 vdd.n592 9.3005
R21883 vdd.n596 vdd.n433 9.3005
R21884 vdd.n600 vdd.n599 9.3005
R21885 vdd.n601 vdd.n432 9.3005
R21886 vdd.n605 vdd.n602 9.3005
R21887 vdd.n606 vdd.n431 9.3005
R21888 vdd.n610 vdd.n609 9.3005
R21889 vdd.n611 vdd.n430 9.3005
R21890 vdd.n615 vdd.n612 9.3005
R21891 vdd.n617 vdd.n429 9.3005
R21892 vdd.n619 vdd.n618 9.3005
R21893 vdd.n3623 vdd.n3622 9.3005
R21894 vdd.n465 vdd.n464 9.3005
R21895 vdd.n3501 vdd.n3500 9.3005
R21896 vdd.n676 vdd.n675 9.3005
R21897 vdd.n3514 vdd.n3513 9.3005
R21898 vdd.n3515 vdd.n674 9.3005
R21899 vdd.n3517 vdd.n3516 9.3005
R21900 vdd.n666 vdd.n665 9.3005
R21901 vdd.n3531 vdd.n3530 9.3005
R21902 vdd.n3532 vdd.n664 9.3005
R21903 vdd.n3534 vdd.n3533 9.3005
R21904 vdd.n653 vdd.n652 9.3005
R21905 vdd.n3547 vdd.n3546 9.3005
R21906 vdd.n3548 vdd.n651 9.3005
R21907 vdd.n3550 vdd.n3549 9.3005
R21908 vdd.n642 vdd.n641 9.3005
R21909 vdd.n3564 vdd.n3563 9.3005
R21910 vdd.n3565 vdd.n640 9.3005
R21911 vdd.n3570 vdd.n3566 9.3005
R21912 vdd.n3569 vdd.n3568 9.3005
R21913 vdd.n3567 vdd.n631 9.3005
R21914 vdd.n3583 vdd.n630 9.3005
R21915 vdd.n3585 vdd.n3584 9.3005
R21916 vdd.n3586 vdd.n629 9.3005
R21917 vdd.n3588 vdd.n3587 9.3005
R21918 vdd.n3590 vdd.n628 9.3005
R21919 vdd.n3592 vdd.n3591 9.3005
R21920 vdd.n3593 vdd.n627 9.3005
R21921 vdd.n3595 vdd.n3594 9.3005
R21922 vdd.n3597 vdd.n626 9.3005
R21923 vdd.n3599 vdd.n3598 9.3005
R21924 vdd.n3600 vdd.n625 9.3005
R21925 vdd.n3602 vdd.n3601 9.3005
R21926 vdd.n3605 vdd.n624 9.3005
R21927 vdd.n3607 vdd.n3606 9.3005
R21928 vdd.n3608 vdd.n623 9.3005
R21929 vdd.n3610 vdd.n3609 9.3005
R21930 vdd.n3612 vdd.n622 9.3005
R21931 vdd.n3614 vdd.n3613 9.3005
R21932 vdd.n3615 vdd.n621 9.3005
R21933 vdd.n3617 vdd.n3616 9.3005
R21934 vdd.n3619 vdd.n620 9.3005
R21935 vdd.n3621 vdd.n3620 9.3005
R21936 vdd.n3499 vdd.n686 9.3005
R21937 vdd.n3498 vdd.n3497 9.3005
R21938 vdd.n3367 vdd.n687 9.3005
R21939 vdd.n3376 vdd.n783 9.3005
R21940 vdd.n3379 vdd.n782 9.3005
R21941 vdd.n3380 vdd.n781 9.3005
R21942 vdd.n3383 vdd.n780 9.3005
R21943 vdd.n3384 vdd.n779 9.3005
R21944 vdd.n3387 vdd.n778 9.3005
R21945 vdd.n3388 vdd.n777 9.3005
R21946 vdd.n3391 vdd.n776 9.3005
R21947 vdd.n3392 vdd.n775 9.3005
R21948 vdd.n3395 vdd.n774 9.3005
R21949 vdd.n3396 vdd.n773 9.3005
R21950 vdd.n3399 vdd.n772 9.3005
R21951 vdd.n3400 vdd.n771 9.3005
R21952 vdd.n3403 vdd.n770 9.3005
R21953 vdd.n3407 vdd.n3406 9.3005
R21954 vdd.n3408 vdd.n767 9.3005
R21955 vdd.n2366 vdd.n2365 9.3005
R21956 vdd.n2361 vdd.n1517 9.3005
R21957 vdd.n1885 vdd.n1884 9.3005
R21958 vdd.n1886 vdd.n1640 9.3005
R21959 vdd.n1888 vdd.n1887 9.3005
R21960 vdd.n1630 vdd.n1629 9.3005
R21961 vdd.n1902 vdd.n1901 9.3005
R21962 vdd.n1903 vdd.n1628 9.3005
R21963 vdd.n1905 vdd.n1904 9.3005
R21964 vdd.n1620 vdd.n1619 9.3005
R21965 vdd.n1919 vdd.n1918 9.3005
R21966 vdd.n1920 vdd.n1618 9.3005
R21967 vdd.n1922 vdd.n1921 9.3005
R21968 vdd.n1607 vdd.n1606 9.3005
R21969 vdd.n1935 vdd.n1934 9.3005
R21970 vdd.n1936 vdd.n1605 9.3005
R21971 vdd.n1938 vdd.n1937 9.3005
R21972 vdd.n1596 vdd.n1595 9.3005
R21973 vdd.n1952 vdd.n1951 9.3005
R21974 vdd.n1953 vdd.n1594 9.3005
R21975 vdd.n1955 vdd.n1954 9.3005
R21976 vdd.n1585 vdd.n1584 9.3005
R21977 vdd.n2275 vdd.n2274 9.3005
R21978 vdd.n2276 vdd.n1583 9.3005
R21979 vdd.n2278 vdd.n2277 9.3005
R21980 vdd.n1573 vdd.n1572 9.3005
R21981 vdd.n2292 vdd.n2291 9.3005
R21982 vdd.n2293 vdd.n1571 9.3005
R21983 vdd.n2295 vdd.n2294 9.3005
R21984 vdd.n1563 vdd.n1562 9.3005
R21985 vdd.n2309 vdd.n2308 9.3005
R21986 vdd.n2310 vdd.n1561 9.3005
R21987 vdd.n2312 vdd.n2311 9.3005
R21988 vdd.n1550 vdd.n1549 9.3005
R21989 vdd.n2325 vdd.n2324 9.3005
R21990 vdd.n2326 vdd.n1548 9.3005
R21991 vdd.n2328 vdd.n2327 9.3005
R21992 vdd.n1540 vdd.n1539 9.3005
R21993 vdd.n2342 vdd.n2341 9.3005
R21994 vdd.n2343 vdd.n1537 9.3005
R21995 vdd.n2347 vdd.n2346 9.3005
R21996 vdd.n2345 vdd.n1538 9.3005
R21997 vdd.n2344 vdd.n1528 9.3005
R21998 vdd.n1642 vdd.n1641 9.3005
R21999 vdd.n1778 vdd.n1777 9.3005
R22000 vdd.n1779 vdd.n1768 9.3005
R22001 vdd.n1781 vdd.n1780 9.3005
R22002 vdd.n1782 vdd.n1767 9.3005
R22003 vdd.n1784 vdd.n1783 9.3005
R22004 vdd.n1785 vdd.n1762 9.3005
R22005 vdd.n1787 vdd.n1786 9.3005
R22006 vdd.n1788 vdd.n1761 9.3005
R22007 vdd.n1790 vdd.n1789 9.3005
R22008 vdd.n1791 vdd.n1756 9.3005
R22009 vdd.n1793 vdd.n1792 9.3005
R22010 vdd.n1794 vdd.n1755 9.3005
R22011 vdd.n1796 vdd.n1795 9.3005
R22012 vdd.n1797 vdd.n1750 9.3005
R22013 vdd.n1799 vdd.n1798 9.3005
R22014 vdd.n1800 vdd.n1749 9.3005
R22015 vdd.n1802 vdd.n1801 9.3005
R22016 vdd.n1803 vdd.n1744 9.3005
R22017 vdd.n1805 vdd.n1804 9.3005
R22018 vdd.n1806 vdd.n1743 9.3005
R22019 vdd.n1808 vdd.n1807 9.3005
R22020 vdd.n1812 vdd.n1739 9.3005
R22021 vdd.n1814 vdd.n1813 9.3005
R22022 vdd.n1815 vdd.n1738 9.3005
R22023 vdd.n1817 vdd.n1816 9.3005
R22024 vdd.n1818 vdd.n1733 9.3005
R22025 vdd.n1820 vdd.n1819 9.3005
R22026 vdd.n1821 vdd.n1732 9.3005
R22027 vdd.n1823 vdd.n1822 9.3005
R22028 vdd.n1824 vdd.n1727 9.3005
R22029 vdd.n1826 vdd.n1825 9.3005
R22030 vdd.n1827 vdd.n1726 9.3005
R22031 vdd.n1829 vdd.n1828 9.3005
R22032 vdd.n1830 vdd.n1721 9.3005
R22033 vdd.n1832 vdd.n1831 9.3005
R22034 vdd.n1833 vdd.n1720 9.3005
R22035 vdd.n1835 vdd.n1834 9.3005
R22036 vdd.n1836 vdd.n1715 9.3005
R22037 vdd.n1838 vdd.n1837 9.3005
R22038 vdd.n1839 vdd.n1714 9.3005
R22039 vdd.n1841 vdd.n1840 9.3005
R22040 vdd.n1842 vdd.n1709 9.3005
R22041 vdd.n1844 vdd.n1843 9.3005
R22042 vdd.n1845 vdd.n1708 9.3005
R22043 vdd.n1847 vdd.n1846 9.3005
R22044 vdd.n1848 vdd.n1701 9.3005
R22045 vdd.n1850 vdd.n1849 9.3005
R22046 vdd.n1851 vdd.n1700 9.3005
R22047 vdd.n1853 vdd.n1852 9.3005
R22048 vdd.n1854 vdd.n1695 9.3005
R22049 vdd.n1856 vdd.n1855 9.3005
R22050 vdd.n1857 vdd.n1694 9.3005
R22051 vdd.n1859 vdd.n1858 9.3005
R22052 vdd.n1860 vdd.n1689 9.3005
R22053 vdd.n1862 vdd.n1861 9.3005
R22054 vdd.n1863 vdd.n1688 9.3005
R22055 vdd.n1865 vdd.n1864 9.3005
R22056 vdd.n1866 vdd.n1683 9.3005
R22057 vdd.n1868 vdd.n1867 9.3005
R22058 vdd.n1869 vdd.n1682 9.3005
R22059 vdd.n1871 vdd.n1870 9.3005
R22060 vdd.n1647 vdd.n1646 9.3005
R22061 vdd.n1877 vdd.n1876 9.3005
R22062 vdd.n1776 vdd.n1775 9.3005
R22063 vdd.n1880 vdd.n1879 9.3005
R22064 vdd.n1636 vdd.n1635 9.3005
R22065 vdd.n1894 vdd.n1893 9.3005
R22066 vdd.n1895 vdd.n1634 9.3005
R22067 vdd.n1897 vdd.n1896 9.3005
R22068 vdd.n1625 vdd.n1624 9.3005
R22069 vdd.n1911 vdd.n1910 9.3005
R22070 vdd.n1912 vdd.n1623 9.3005
R22071 vdd.n1914 vdd.n1913 9.3005
R22072 vdd.n1614 vdd.n1613 9.3005
R22073 vdd.n1927 vdd.n1926 9.3005
R22074 vdd.n1928 vdd.n1612 9.3005
R22075 vdd.n1930 vdd.n1929 9.3005
R22076 vdd.n1602 vdd.n1601 9.3005
R22077 vdd.n1944 vdd.n1943 9.3005
R22078 vdd.n1945 vdd.n1600 9.3005
R22079 vdd.n1947 vdd.n1946 9.3005
R22080 vdd.n1591 vdd.n1590 9.3005
R22081 vdd.n1960 vdd.n1959 9.3005
R22082 vdd.n1961 vdd.n1589 9.3005
R22083 vdd.n1878 vdd.n1645 9.3005
R22084 vdd.n2181 vdd.n2180 9.3005
R22085 vdd.n2176 vdd.n2175 9.3005
R22086 vdd.n2187 vdd.n2186 9.3005
R22087 vdd.n2189 vdd.n2188 9.3005
R22088 vdd.n2172 vdd.n2171 9.3005
R22089 vdd.n2195 vdd.n2194 9.3005
R22090 vdd.n2197 vdd.n2196 9.3005
R22091 vdd.n2169 vdd.n2166 9.3005
R22092 vdd.n2204 vdd.n2203 9.3005
R22093 vdd.n2240 vdd.n2239 9.3005
R22094 vdd.n2235 vdd.n2234 9.3005
R22095 vdd.n2246 vdd.n2245 9.3005
R22096 vdd.n2248 vdd.n2247 9.3005
R22097 vdd.n2231 vdd.n2230 9.3005
R22098 vdd.n2254 vdd.n2253 9.3005
R22099 vdd.n2256 vdd.n2255 9.3005
R22100 vdd.n2228 vdd.n2225 9.3005
R22101 vdd.n2263 vdd.n2262 9.3005
R22102 vdd.n2079 vdd.n2078 9.3005
R22103 vdd.n2074 vdd.n2073 9.3005
R22104 vdd.n2085 vdd.n2084 9.3005
R22105 vdd.n2087 vdd.n2086 9.3005
R22106 vdd.n2070 vdd.n2069 9.3005
R22107 vdd.n2093 vdd.n2092 9.3005
R22108 vdd.n2095 vdd.n2094 9.3005
R22109 vdd.n2067 vdd.n2064 9.3005
R22110 vdd.n2102 vdd.n2101 9.3005
R22111 vdd.n2138 vdd.n2137 9.3005
R22112 vdd.n2133 vdd.n2132 9.3005
R22113 vdd.n2144 vdd.n2143 9.3005
R22114 vdd.n2146 vdd.n2145 9.3005
R22115 vdd.n2129 vdd.n2128 9.3005
R22116 vdd.n2152 vdd.n2151 9.3005
R22117 vdd.n2154 vdd.n2153 9.3005
R22118 vdd.n2126 vdd.n2123 9.3005
R22119 vdd.n2161 vdd.n2160 9.3005
R22120 vdd.n1978 vdd.n1977 9.3005
R22121 vdd.n1973 vdd.n1972 9.3005
R22122 vdd.n1984 vdd.n1983 9.3005
R22123 vdd.n1986 vdd.n1985 9.3005
R22124 vdd.n1969 vdd.n1968 9.3005
R22125 vdd.n1992 vdd.n1991 9.3005
R22126 vdd.n1994 vdd.n1993 9.3005
R22127 vdd.n1966 vdd.n1963 9.3005
R22128 vdd.n2001 vdd.n2000 9.3005
R22129 vdd.n2037 vdd.n2036 9.3005
R22130 vdd.n2032 vdd.n2031 9.3005
R22131 vdd.n2043 vdd.n2042 9.3005
R22132 vdd.n2045 vdd.n2044 9.3005
R22133 vdd.n2028 vdd.n2027 9.3005
R22134 vdd.n2051 vdd.n2050 9.3005
R22135 vdd.n2053 vdd.n2052 9.3005
R22136 vdd.n2025 vdd.n2022 9.3005
R22137 vdd.n2060 vdd.n2059 9.3005
R22138 vdd.n1916 vdd.t128 9.18308
R22139 vdd.n3603 vdd.t2 9.18308
R22140 vdd.n1610 vdd.t76 8.95635
R22141 vdd.n2358 vdd.t169 8.95635
R22142 vdd.n723 vdd.t186 8.95635
R22143 vdd.t74 vdd.n3657 8.95635
R22144 vdd.n312 vdd.n311 8.92171
R22145 vdd.n253 vdd.n252 8.92171
R22146 vdd.n210 vdd.n209 8.92171
R22147 vdd.n151 vdd.n150 8.92171
R22148 vdd.n109 vdd.n108 8.92171
R22149 vdd.n50 vdd.n49 8.92171
R22150 vdd.n2186 vdd.n2185 8.92171
R22151 vdd.n2245 vdd.n2244 8.92171
R22152 vdd.n2084 vdd.n2083 8.92171
R22153 vdd.n2143 vdd.n2142 8.92171
R22154 vdd.n1983 vdd.n1982 8.92171
R22155 vdd.n2042 vdd.n2041 8.92171
R22156 vdd.n231 vdd.n129 8.81535
R22157 vdd.n2164 vdd.n2062 8.81535
R22158 vdd.n1957 vdd.t0 8.72962
R22159 vdd.t116 vdd.n3666 8.72962
R22160 vdd.n2280 vdd.t8 8.50289
R22161 vdd.n3572 vdd.t64 8.50289
R22162 vdd.n28 vdd.n14 8.42249
R22163 vdd.n2306 vdd.t37 8.27616
R22164 vdd.t112 vdd.n656 8.27616
R22165 vdd.n3672 vdd.n3671 8.16225
R22166 vdd.n2268 vdd.n2267 8.16225
R22167 vdd.n308 vdd.n302 8.14595
R22168 vdd.n249 vdd.n243 8.14595
R22169 vdd.n206 vdd.n200 8.14595
R22170 vdd.n147 vdd.n141 8.14595
R22171 vdd.n105 vdd.n99 8.14595
R22172 vdd.n46 vdd.n40 8.14595
R22173 vdd.n2182 vdd.n2176 8.14595
R22174 vdd.n2241 vdd.n2235 8.14595
R22175 vdd.n2080 vdd.n2074 8.14595
R22176 vdd.n2139 vdd.n2133 8.14595
R22177 vdd.n1979 vdd.n1973 8.14595
R22178 vdd.n2038 vdd.n2032 8.14595
R22179 vdd.n1553 vdd.t92 8.04943
R22180 vdd.n3528 vdd.t50 8.04943
R22181 vdd.n2513 vdd.n1134 7.70933
R22182 vdd.n2513 vdd.n1137 7.70933
R22183 vdd.n2519 vdd.n1123 7.70933
R22184 vdd.n2525 vdd.n1123 7.70933
R22185 vdd.n2525 vdd.n1116 7.70933
R22186 vdd.n2531 vdd.n1116 7.70933
R22187 vdd.n2531 vdd.n1119 7.70933
R22188 vdd.n2537 vdd.n1112 7.70933
R22189 vdd.n2543 vdd.n1106 7.70933
R22190 vdd.n2549 vdd.n1093 7.70933
R22191 vdd.n2555 vdd.n1093 7.70933
R22192 vdd.n2561 vdd.n1087 7.70933
R22193 vdd.n2567 vdd.n1080 7.70933
R22194 vdd.n2567 vdd.n1083 7.70933
R22195 vdd.n2573 vdd.n1076 7.70933
R22196 vdd.n2580 vdd.n1062 7.70933
R22197 vdd.n2586 vdd.n1062 7.70933
R22198 vdd.n2592 vdd.n1056 7.70933
R22199 vdd.n2598 vdd.n1052 7.70933
R22200 vdd.n2604 vdd.n1046 7.70933
R22201 vdd.n2622 vdd.n1028 7.70933
R22202 vdd.n2622 vdd.n1021 7.70933
R22203 vdd.n2630 vdd.n1021 7.70933
R22204 vdd.n2712 vdd.n1005 7.70933
R22205 vdd.n3095 vdd.n957 7.70933
R22206 vdd.n3107 vdd.n946 7.70933
R22207 vdd.n3107 vdd.n940 7.70933
R22208 vdd.n3113 vdd.n940 7.70933
R22209 vdd.n3125 vdd.n931 7.70933
R22210 vdd.n3131 vdd.n925 7.70933
R22211 vdd.n3143 vdd.n912 7.70933
R22212 vdd.n3150 vdd.n905 7.70933
R22213 vdd.n3150 vdd.n908 7.70933
R22214 vdd.n3156 vdd.n901 7.70933
R22215 vdd.n3162 vdd.n887 7.70933
R22216 vdd.n3168 vdd.n887 7.70933
R22217 vdd.n3174 vdd.n881 7.70933
R22218 vdd.n3180 vdd.n874 7.70933
R22219 vdd.n3180 vdd.n877 7.70933
R22220 vdd.n3186 vdd.n870 7.70933
R22221 vdd.n3192 vdd.n864 7.70933
R22222 vdd.n3198 vdd.n851 7.70933
R22223 vdd.n3204 vdd.n851 7.70933
R22224 vdd.n3204 vdd.n843 7.70933
R22225 vdd.n3255 vdd.n843 7.70933
R22226 vdd.n3255 vdd.n846 7.70933
R22227 vdd.n3261 vdd.n805 7.70933
R22228 vdd.n3331 vdd.n805 7.70933
R22229 vdd.n307 vdd.n304 7.3702
R22230 vdd.n248 vdd.n245 7.3702
R22231 vdd.n205 vdd.n202 7.3702
R22232 vdd.n146 vdd.n143 7.3702
R22233 vdd.n104 vdd.n101 7.3702
R22234 vdd.n45 vdd.n42 7.3702
R22235 vdd.n2181 vdd.n2178 7.3702
R22236 vdd.n2240 vdd.n2237 7.3702
R22237 vdd.n2079 vdd.n2076 7.3702
R22238 vdd.n2138 vdd.n2135 7.3702
R22239 vdd.n1978 vdd.n1975 7.3702
R22240 vdd.n2037 vdd.n2034 7.3702
R22241 vdd.n1106 vdd.t289 7.36923
R22242 vdd.n3186 vdd.t266 7.36923
R22243 vdd.n2339 vdd.t42 7.1425
R22244 vdd.n2537 vdd.t241 7.1425
R22245 vdd.n1425 vdd.t237 7.1425
R22246 vdd.n3119 vdd.t240 7.1425
R22247 vdd.n864 vdd.t250 7.1425
R22248 vdd.n679 vdd.t81 7.1425
R22249 vdd.n1813 vdd.n1812 6.98232
R22250 vdd.n2401 vdd.n2400 6.98232
R22251 vdd.n566 vdd.n565 6.98232
R22252 vdd.n3413 vdd.n3410 6.98232
R22253 vdd.t10 vdd.n1552 6.91577
R22254 vdd.n3536 vdd.t25 6.91577
R22255 vdd.n1425 vdd.t238 6.80241
R22256 vdd.n3119 vdd.t284 6.80241
R22257 vdd.n2298 vdd.t4 6.68904
R22258 vdd.n3552 vdd.t79 6.68904
R22259 vdd.t90 vdd.n1581 6.46231
R22260 vdd.n2561 vdd.t248 6.46231
R22261 vdd.t253 vdd.n1056 6.46231
R22262 vdd.n3143 vdd.t258 6.46231
R22263 vdd.t274 vdd.n881 6.46231
R22264 vdd.n3580 vdd.t56 6.46231
R22265 vdd.n3672 vdd.n333 6.38151
R22266 vdd.n2267 vdd.n2266 6.38151
R22267 vdd.n2637 vdd.t281 6.34895
R22268 vdd.n3016 vdd.t271 6.34895
R22269 vdd.n3158 vdd.n897 6.2444
R22270 vdd.n2577 vdd.n2576 6.2444
R22271 vdd.n1949 vdd.t110 6.23558
R22272 vdd.t48 vdd.n344 6.23558
R22273 vdd.t94 vdd.n1609 6.00885
R22274 vdd.n3651 vdd.t20 6.00885
R22275 vdd.n2598 vdd.t279 5.89549
R22276 vdd.n925 vdd.t254 5.89549
R22277 vdd.n308 vdd.n307 5.81868
R22278 vdd.n249 vdd.n248 5.81868
R22279 vdd.n206 vdd.n205 5.81868
R22280 vdd.n147 vdd.n146 5.81868
R22281 vdd.n105 vdd.n104 5.81868
R22282 vdd.n46 vdd.n45 5.81868
R22283 vdd.n2182 vdd.n2181 5.81868
R22284 vdd.n2241 vdd.n2240 5.81868
R22285 vdd.n2080 vdd.n2079 5.81868
R22286 vdd.n2139 vdd.n2138 5.81868
R22287 vdd.n1979 vdd.n1978 5.81868
R22288 vdd.n2038 vdd.n2037 5.81868
R22289 vdd.n1908 vdd.t84 5.78212
R22290 vdd.n3642 vdd.t12 5.78212
R22291 vdd.n2720 vdd.n2719 5.77611
R22292 vdd.n1349 vdd.n1348 5.77611
R22293 vdd.n3028 vdd.n3027 5.77611
R22294 vdd.n3272 vdd.n3271 5.77611
R22295 vdd.n3336 vdd.n801 5.77611
R22296 vdd.n2891 vdd.n2825 5.77611
R22297 vdd.n2645 vdd.n1012 5.77611
R22298 vdd.n1485 vdd.n1317 5.77611
R22299 vdd.n1775 vdd.n1774 5.62474
R22300 vdd.n2364 vdd.n2361 5.62474
R22301 vdd.n3623 vdd.n428 5.62474
R22302 vdd.n3497 vdd.n690 5.62474
R22303 vdd.n1632 vdd.t84 5.55539
R22304 vdd.n2573 vdd.t268 5.55539
R22305 vdd.n901 vdd.t244 5.55539
R22306 vdd.t12 vdd.n3641 5.55539
R22307 vdd.n1924 vdd.t94 5.32866
R22308 vdd.t20 vdd.n3650 5.32866
R22309 vdd.n1940 vdd.t110 5.10193
R22310 vdd.n3659 vdd.t48 5.10193
R22311 vdd.n311 vdd.n302 5.04292
R22312 vdd.n252 vdd.n243 5.04292
R22313 vdd.n209 vdd.n200 5.04292
R22314 vdd.n150 vdd.n141 5.04292
R22315 vdd.n108 vdd.n99 5.04292
R22316 vdd.n49 vdd.n40 5.04292
R22317 vdd.n2185 vdd.n2176 5.04292
R22318 vdd.n2244 vdd.n2235 5.04292
R22319 vdd.n2083 vdd.n2074 5.04292
R22320 vdd.n2142 vdd.n2133 5.04292
R22321 vdd.n1982 vdd.n1973 5.04292
R22322 vdd.n2041 vdd.n2032 5.04292
R22323 vdd.n2272 vdd.t90 4.8752
R22324 vdd.t247 vdd.t260 4.8752
R22325 vdd.t290 vdd.t236 4.8752
R22326 vdd.t56 vdd.n340 4.8752
R22327 vdd.n2721 vdd.n2720 4.83952
R22328 vdd.n1348 vdd.n1347 4.83952
R22329 vdd.n3029 vdd.n3028 4.83952
R22330 vdd.n3273 vdd.n3272 4.83952
R22331 vdd.n801 vdd.n796 4.83952
R22332 vdd.n2888 vdd.n2825 4.83952
R22333 vdd.n2648 vdd.n1012 4.83952
R22334 vdd.n1488 vdd.n1317 4.83952
R22335 vdd.n1399 vdd.t256 4.76184
R22336 vdd.n3101 vdd.t242 4.76184
R22337 vdd.n2369 vdd.n2368 4.74817
R22338 vdd.n1521 vdd.n1516 4.74817
R22339 vdd.n1183 vdd.n1180 4.74817
R22340 vdd.n2462 vdd.n1179 4.74817
R22341 vdd.n2467 vdd.n1180 4.74817
R22342 vdd.n2466 vdd.n1179 4.74817
R22343 vdd.n3490 vdd.n3489 4.74817
R22344 vdd.n3487 vdd.n3486 4.74817
R22345 vdd.n3487 vdd.n732 4.74817
R22346 vdd.n3489 vdd.n729 4.74817
R22347 vdd.n3372 vdd.n784 4.74817
R22348 vdd.n3368 vdd.n3366 4.74817
R22349 vdd.n3371 vdd.n3366 4.74817
R22350 vdd.n3375 vdd.n784 4.74817
R22351 vdd.n2368 vdd.n1279 4.74817
R22352 vdd.n1518 vdd.n1516 4.74817
R22353 vdd.n333 vdd.n332 4.7074
R22354 vdd.n231 vdd.n230 4.7074
R22355 vdd.n2266 vdd.n2265 4.7074
R22356 vdd.n2164 vdd.n2163 4.7074
R22357 vdd.n1575 vdd.t4 4.64847
R22358 vdd.t249 vdd.n1087 4.64847
R22359 vdd.n2592 vdd.t288 4.64847
R22360 vdd.t277 vdd.n912 4.64847
R22361 vdd.n3174 vdd.t273 4.64847
R22362 vdd.n3561 vdd.t79 4.64847
R22363 vdd.n1076 vdd.t217 4.53511
R22364 vdd.n3156 vdd.t190 4.53511
R22365 vdd.n2314 vdd.t10 4.42174
R22366 vdd.n2519 vdd.t165 4.42174
R22367 vdd.n1399 vdd.t206 4.42174
R22368 vdd.n3101 vdd.t213 4.42174
R22369 vdd.n846 vdd.t161 4.42174
R22370 vdd.t25 vdd.n655 4.42174
R22371 vdd.n3147 vdd.n897 4.37123
R22372 vdd.n2578 vdd.n2577 4.37123
R22373 vdd.n2616 vdd.t275 4.30838
R22374 vdd.n3004 vdd.t262 4.30838
R22375 vdd.n312 vdd.n300 4.26717
R22376 vdd.n253 vdd.n241 4.26717
R22377 vdd.n210 vdd.n198 4.26717
R22378 vdd.n151 vdd.n139 4.26717
R22379 vdd.n109 vdd.n97 4.26717
R22380 vdd.n50 vdd.n38 4.26717
R22381 vdd.n2186 vdd.n2174 4.26717
R22382 vdd.n2245 vdd.n2233 4.26717
R22383 vdd.n2084 vdd.n2072 4.26717
R22384 vdd.n2143 vdd.n2131 4.26717
R22385 vdd.n1983 vdd.n1971 4.26717
R22386 vdd.n2042 vdd.n2030 4.26717
R22387 vdd.n2330 vdd.t42 4.19501
R22388 vdd.n3520 vdd.t81 4.19501
R22389 vdd.n333 vdd.n231 4.10845
R22390 vdd.n2266 vdd.n2164 4.10845
R22391 vdd.n289 vdd.t148 4.06363
R22392 vdd.n289 vdd.t31 4.06363
R22393 vdd.n287 vdd.t41 4.06363
R22394 vdd.n287 vdd.t69 4.06363
R22395 vdd.n285 vdd.t109 4.06363
R22396 vdd.n285 vdd.t153 4.06363
R22397 vdd.n283 vdd.t19 4.06363
R22398 vdd.n283 vdd.t71 4.06363
R22399 vdd.n281 vdd.t73 4.06363
R22400 vdd.n281 vdd.t126 4.06363
R22401 vdd.n279 vdd.t130 4.06363
R22402 vdd.n279 vdd.t7 4.06363
R22403 vdd.n277 vdd.t35 4.06363
R22404 vdd.n277 vdd.t101 4.06363
R22405 vdd.n275 vdd.t131 4.06363
R22406 vdd.n275 vdd.t149 4.06363
R22407 vdd.n273 vdd.t154 4.06363
R22408 vdd.n273 vdd.t46 4.06363
R22409 vdd.n187 vdd.t132 4.06363
R22410 vdd.n187 vdd.t13 4.06363
R22411 vdd.n185 vdd.t21 4.06363
R22412 vdd.n185 vdd.t47 4.06363
R22413 vdd.n183 vdd.t99 4.06363
R22414 vdd.n183 vdd.t140 4.06363
R22415 vdd.n181 vdd.t158 4.06363
R22416 vdd.n181 vdd.t49 4.06363
R22417 vdd.n179 vdd.t57 4.06363
R22418 vdd.n179 vdd.t117 4.06363
R22419 vdd.n177 vdd.t118 4.06363
R22420 vdd.n177 vdd.t150 4.06363
R22421 vdd.n175 vdd.t17 4.06363
R22422 vdd.n175 vdd.t80 4.06363
R22423 vdd.n173 vdd.t121 4.06363
R22424 vdd.n173 vdd.t133 4.06363
R22425 vdd.n171 vdd.t142 4.06363
R22426 vdd.n171 vdd.t23 4.06363
R22427 vdd.n86 vdd.t67 4.06363
R22428 vdd.n86 vdd.t145 4.06363
R22429 vdd.n84 vdd.t100 4.06363
R22430 vdd.n84 vdd.t3 4.06363
R22431 vdd.n82 vdd.t75 4.06363
R22432 vdd.n82 vdd.t155 4.06363
R22433 vdd.n80 vdd.t54 4.06363
R22434 vdd.n80 vdd.t136 4.06363
R22435 vdd.n78 vdd.t89 4.06363
R22436 vdd.n78 vdd.t119 4.06363
R22437 vdd.n76 vdd.t65 4.06363
R22438 vdd.n76 vdd.t144 4.06363
R22439 vdd.n74 vdd.t34 4.06363
R22440 vdd.n74 vdd.t127 4.06363
R22441 vdd.n72 vdd.t26 4.06363
R22442 vdd.n72 vdd.t113 4.06363
R22443 vdd.n70 vdd.t51 4.06363
R22444 vdd.n70 vdd.t134 4.06363
R22445 vdd.n2206 vdd.t108 4.06363
R22446 vdd.n2206 vdd.t106 4.06363
R22447 vdd.n2208 vdd.t59 4.06363
R22448 vdd.n2208 vdd.t30 4.06363
R22449 vdd.n2210 vdd.t28 4.06363
R22450 vdd.n2210 vdd.t104 4.06363
R22451 vdd.n2212 vdd.t78 4.06363
R22452 vdd.n2212 vdd.t29 4.06363
R22453 vdd.n2214 vdd.t24 4.06363
R22454 vdd.n2214 vdd.t125 4.06363
R22455 vdd.n2216 vdd.t123 4.06363
R22456 vdd.n2216 vdd.t72 4.06363
R22457 vdd.n2218 vdd.t63 4.06363
R22458 vdd.n2218 vdd.t157 4.06363
R22459 vdd.n2220 vdd.t151 4.06363
R22460 vdd.n2220 vdd.t107 4.06363
R22461 vdd.n2222 vdd.t103 4.06363
R22462 vdd.n2222 vdd.t58 4.06363
R22463 vdd.n2104 vdd.t97 4.06363
R22464 vdd.n2104 vdd.t93 4.06363
R22465 vdd.n2106 vdd.t38 4.06363
R22466 vdd.n2106 vdd.t11 4.06363
R22467 vdd.n2108 vdd.t5 4.06363
R22468 vdd.n2108 vdd.t86 4.06363
R22469 vdd.n2110 vdd.t61 4.06363
R22470 vdd.n2110 vdd.t9 4.06363
R22471 vdd.n2112 vdd.t1 4.06363
R22472 vdd.n2112 vdd.t115 4.06363
R22473 vdd.n2114 vdd.t111 4.06363
R22474 vdd.n2114 vdd.t55 4.06363
R22475 vdd.n2116 vdd.t45 4.06363
R22476 vdd.n2116 vdd.t143 4.06363
R22477 vdd.n2118 vdd.t138 4.06363
R22478 vdd.n2118 vdd.t95 4.06363
R22479 vdd.n2120 vdd.t85 4.06363
R22480 vdd.n2120 vdd.t33 4.06363
R22481 vdd.n2003 vdd.t135 4.06363
R22482 vdd.n2003 vdd.t159 4.06363
R22483 vdd.n2005 vdd.t114 4.06363
R22484 vdd.n2005 vdd.t27 4.06363
R22485 vdd.n2007 vdd.t98 4.06363
R22486 vdd.n2007 vdd.t40 4.06363
R22487 vdd.n2009 vdd.t146 4.06363
R22488 vdd.n2009 vdd.t68 4.06363
R22489 vdd.n2011 vdd.t120 4.06363
R22490 vdd.n2011 vdd.t91 4.06363
R22491 vdd.n2013 vdd.t137 4.06363
R22492 vdd.n2013 vdd.t53 4.06363
R22493 vdd.n2015 vdd.t156 4.06363
R22494 vdd.n2015 vdd.t77 4.06363
R22495 vdd.n2017 vdd.t129 4.06363
R22496 vdd.n2017 vdd.t102 4.06363
R22497 vdd.n2019 vdd.t147 4.06363
R22498 vdd.n2019 vdd.t70 4.06363
R22499 vdd.n1112 vdd.t283 3.96828
R22500 vdd.n2610 vdd.t259 3.96828
R22501 vdd.n2998 vdd.t278 3.96828
R22502 vdd.n3192 vdd.t267 3.96828
R22503 vdd.n26 vdd.t307 3.9605
R22504 vdd.n26 vdd.t292 3.9605
R22505 vdd.n23 vdd.t296 3.9605
R22506 vdd.n23 vdd.t302 3.9605
R22507 vdd.n21 vdd.t303 3.9605
R22508 vdd.n21 vdd.t306 3.9605
R22509 vdd.n20 vdd.t304 3.9605
R22510 vdd.n20 vdd.t295 3.9605
R22511 vdd.n15 vdd.t300 3.9605
R22512 vdd.n15 vdd.t297 3.9605
R22513 vdd.n16 vdd.t301 3.9605
R22514 vdd.n16 vdd.t294 3.9605
R22515 vdd.n18 vdd.t299 3.9605
R22516 vdd.n18 vdd.t305 3.9605
R22517 vdd.n25 vdd.t293 3.9605
R22518 vdd.n25 vdd.t298 3.9605
R22519 vdd.n2543 vdd.t283 3.74155
R22520 vdd.n1046 vdd.t259 3.74155
R22521 vdd.n3125 vdd.t278 3.74155
R22522 vdd.n870 vdd.t267 3.74155
R22523 vdd.n7 vdd.t291 3.61217
R22524 vdd.n7 vdd.t255 3.61217
R22525 vdd.n8 vdd.t263 3.61217
R22526 vdd.n8 vdd.t285 3.61217
R22527 vdd.n10 vdd.t272 3.61217
R22528 vdd.n10 vdd.t243 3.61217
R22529 vdd.n12 vdd.t252 3.61217
R22530 vdd.n12 vdd.t270 3.61217
R22531 vdd.n5 vdd.t287 3.61217
R22532 vdd.n5 vdd.t265 3.61217
R22533 vdd.n3 vdd.t257 3.61217
R22534 vdd.n3 vdd.t282 3.61217
R22535 vdd.n1 vdd.t239 3.61217
R22536 vdd.n1 vdd.t276 3.61217
R22537 vdd.n0 vdd.t280 3.61217
R22538 vdd.n0 vdd.t261 3.61217
R22539 vdd.n316 vdd.n315 3.49141
R22540 vdd.n257 vdd.n256 3.49141
R22541 vdd.n214 vdd.n213 3.49141
R22542 vdd.n155 vdd.n154 3.49141
R22543 vdd.n113 vdd.n112 3.49141
R22544 vdd.n54 vdd.n53 3.49141
R22545 vdd.n2190 vdd.n2189 3.49141
R22546 vdd.n2249 vdd.n2248 3.49141
R22547 vdd.n2088 vdd.n2087 3.49141
R22548 vdd.n2147 vdd.n2146 3.49141
R22549 vdd.n1987 vdd.n1986 3.49141
R22550 vdd.n2046 vdd.n2045 3.49141
R22551 vdd.t275 vdd.n1028 3.40145
R22552 vdd.n2784 vdd.t286 3.40145
R22553 vdd.n3088 vdd.t269 3.40145
R22554 vdd.n3113 vdd.t262 3.40145
R22555 vdd.n2331 vdd.t92 3.28809
R22556 vdd.n1137 vdd.t165 3.28809
R22557 vdd.n2637 vdd.t206 3.28809
R22558 vdd.n3016 vdd.t213 3.28809
R22559 vdd.n3261 vdd.t161 3.28809
R22560 vdd.n3519 vdd.t50 3.28809
R22561 vdd.t37 vdd.n1559 3.06136
R22562 vdd.n2555 vdd.t249 3.06136
R22563 vdd.n1437 vdd.t288 3.06136
R22564 vdd.n3137 vdd.t277 3.06136
R22565 vdd.t273 vdd.n874 3.06136
R22566 vdd.n3544 vdd.t112 3.06136
R22567 vdd.n2630 vdd.t256 2.94799
R22568 vdd.t242 vdd.n946 2.94799
R22569 vdd.n2289 vdd.t8 2.83463
R22570 vdd.n644 vdd.t64 2.83463
R22571 vdd.n319 vdd.n298 2.71565
R22572 vdd.n260 vdd.n239 2.71565
R22573 vdd.n217 vdd.n196 2.71565
R22574 vdd.n158 vdd.n137 2.71565
R22575 vdd.n116 vdd.n95 2.71565
R22576 vdd.n57 vdd.n36 2.71565
R22577 vdd.n2193 vdd.n2172 2.71565
R22578 vdd.n2252 vdd.n2231 2.71565
R22579 vdd.n2091 vdd.n2070 2.71565
R22580 vdd.n2150 vdd.n2129 2.71565
R22581 vdd.n1990 vdd.n1969 2.71565
R22582 vdd.n2049 vdd.n2028 2.71565
R22583 vdd.t0 vdd.n1587 2.6079
R22584 vdd.n3667 vdd.t116 2.6079
R22585 vdd.n2604 vdd.t260 2.49453
R22586 vdd.n931 vdd.t290 2.49453
R22587 vdd.n306 vdd.n305 2.4129
R22588 vdd.n247 vdd.n246 2.4129
R22589 vdd.n204 vdd.n203 2.4129
R22590 vdd.n145 vdd.n144 2.4129
R22591 vdd.n103 vdd.n102 2.4129
R22592 vdd.n44 vdd.n43 2.4129
R22593 vdd.n2180 vdd.n2179 2.4129
R22594 vdd.n2239 vdd.n2238 2.4129
R22595 vdd.n2078 vdd.n2077 2.4129
R22596 vdd.n2137 vdd.n2136 2.4129
R22597 vdd.n1977 vdd.n1976 2.4129
R22598 vdd.n2036 vdd.n2035 2.4129
R22599 vdd.n1941 vdd.t76 2.38117
R22600 vdd.n2349 vdd.t169 2.38117
R22601 vdd.n3503 vdd.t186 2.38117
R22602 vdd.n3658 vdd.t74 2.38117
R22603 vdd.n2474 vdd.n1180 2.27742
R22604 vdd.n2474 vdd.n1179 2.27742
R22605 vdd.n3488 vdd.n3487 2.27742
R22606 vdd.n3489 vdd.n3488 2.27742
R22607 vdd.n3366 vdd.n3365 2.27742
R22608 vdd.n3365 vdd.n784 2.27742
R22609 vdd.n2368 vdd.n2367 2.27742
R22610 vdd.n2367 vdd.n1516 2.27742
R22611 vdd.t128 vdd.n1616 2.15444
R22612 vdd.n1083 vdd.t268 2.15444
R22613 vdd.n2580 vdd.t246 2.15444
R22614 vdd.n908 vdd.t245 2.15444
R22615 vdd.n3162 vdd.t244 2.15444
R22616 vdd.n3649 vdd.t2 2.15444
R22617 vdd.n320 vdd.n296 1.93989
R22618 vdd.n261 vdd.n237 1.93989
R22619 vdd.n218 vdd.n194 1.93989
R22620 vdd.n159 vdd.n135 1.93989
R22621 vdd.n117 vdd.n93 1.93989
R22622 vdd.n58 vdd.n34 1.93989
R22623 vdd.n2194 vdd.n2170 1.93989
R22624 vdd.n2253 vdd.n2229 1.93989
R22625 vdd.n2092 vdd.n2068 1.93989
R22626 vdd.n2151 vdd.n2127 1.93989
R22627 vdd.n1991 vdd.n1967 1.93989
R22628 vdd.n2050 vdd.n2026 1.93989
R22629 vdd.n1899 vdd.t87 1.92771
R22630 vdd.t14 vdd.n375 1.92771
R22631 vdd.n1437 vdd.t279 1.81434
R22632 vdd.n3137 vdd.t254 1.81434
R22633 vdd.n1907 vdd.t32 1.70098
R22634 vdd.n3643 vdd.t66 1.70098
R22635 vdd.n1932 vdd.t44 1.47425
R22636 vdd.n361 vdd.t139 1.47425
R22637 vdd.t281 vdd.n1005 1.36088
R22638 vdd.n3095 vdd.t271 1.36088
R22639 vdd.n1598 vdd.t52 1.24752
R22640 vdd.t248 vdd.n1080 1.24752
R22641 vdd.n2586 vdd.t253 1.24752
R22642 vdd.t258 vdd.n905 1.24752
R22643 vdd.n3168 vdd.t274 1.24752
R22644 vdd.t18 vdd.n3665 1.24752
R22645 vdd.n2267 vdd.n28 1.21639
R22646 vdd vdd.n3672 1.20856
R22647 vdd.n331 vdd.n291 1.16414
R22648 vdd.n324 vdd.n323 1.16414
R22649 vdd.n272 vdd.n232 1.16414
R22650 vdd.n265 vdd.n264 1.16414
R22651 vdd.n229 vdd.n189 1.16414
R22652 vdd.n222 vdd.n221 1.16414
R22653 vdd.n170 vdd.n130 1.16414
R22654 vdd.n163 vdd.n162 1.16414
R22655 vdd.n128 vdd.n88 1.16414
R22656 vdd.n121 vdd.n120 1.16414
R22657 vdd.n69 vdd.n29 1.16414
R22658 vdd.n62 vdd.n61 1.16414
R22659 vdd.n2205 vdd.n2165 1.16414
R22660 vdd.n2198 vdd.n2197 1.16414
R22661 vdd.n2264 vdd.n2224 1.16414
R22662 vdd.n2257 vdd.n2256 1.16414
R22663 vdd.n2103 vdd.n2063 1.16414
R22664 vdd.n2096 vdd.n2095 1.16414
R22665 vdd.n2162 vdd.n2122 1.16414
R22666 vdd.n2155 vdd.n2154 1.16414
R22667 vdd.n2002 vdd.n1962 1.16414
R22668 vdd.n1995 vdd.n1994 1.16414
R22669 vdd.n2061 vdd.n2021 1.16414
R22670 vdd.n2054 vdd.n2053 1.16414
R22671 vdd.n2281 vdd.t60 1.02079
R22672 vdd.t217 vdd.t246 1.02079
R22673 vdd.t245 vdd.t190 1.02079
R22674 vdd.t6 vdd.n633 1.02079
R22675 vdd.n1778 vdd.n1774 0.970197
R22676 vdd.n2365 vdd.n2364 0.970197
R22677 vdd.n618 vdd.n428 0.970197
R22678 vdd.n3367 vdd.n690 0.970197
R22679 vdd.n2610 vdd.t238 0.907421
R22680 vdd.n2998 vdd.t284 0.907421
R22681 vdd.n2297 vdd.t39 0.794056
R22682 vdd.n3553 vdd.t16 0.794056
R22683 vdd.n2322 vdd.t96 0.567326
R22684 vdd.n1119 vdd.t241 0.567326
R22685 vdd.n2616 vdd.t237 0.567326
R22686 vdd.n3004 vdd.t240 0.567326
R22687 vdd.n3198 vdd.t250 0.567326
R22688 vdd.t22 vdd.n662 0.567326
R22689 vdd.n2355 vdd.n1181 0.530988
R22690 vdd.n726 vdd.n682 0.530988
R22691 vdd.n464 vdd.n391 0.530988
R22692 vdd.n3622 vdd.n3621 0.530988
R22693 vdd.n3499 vdd.n3498 0.530988
R22694 vdd.n2344 vdd.n1517 0.530988
R22695 vdd.n1776 vdd.n1641 0.530988
R22696 vdd.n1878 vdd.n1877 0.530988
R22697 vdd.n4 vdd.n2 0.459552
R22698 vdd.n11 vdd.n9 0.459552
R22699 vdd.n329 vdd.n328 0.388379
R22700 vdd.n295 vdd.n293 0.388379
R22701 vdd.n270 vdd.n269 0.388379
R22702 vdd.n236 vdd.n234 0.388379
R22703 vdd.n227 vdd.n226 0.388379
R22704 vdd.n193 vdd.n191 0.388379
R22705 vdd.n168 vdd.n167 0.388379
R22706 vdd.n134 vdd.n132 0.388379
R22707 vdd.n126 vdd.n125 0.388379
R22708 vdd.n92 vdd.n90 0.388379
R22709 vdd.n67 vdd.n66 0.388379
R22710 vdd.n33 vdd.n31 0.388379
R22711 vdd.n2203 vdd.n2202 0.388379
R22712 vdd.n2169 vdd.n2167 0.388379
R22713 vdd.n2262 vdd.n2261 0.388379
R22714 vdd.n2228 vdd.n2226 0.388379
R22715 vdd.n2101 vdd.n2100 0.388379
R22716 vdd.n2067 vdd.n2065 0.388379
R22717 vdd.n2160 vdd.n2159 0.388379
R22718 vdd.n2126 vdd.n2124 0.388379
R22719 vdd.n2000 vdd.n1999 0.388379
R22720 vdd.n1966 vdd.n1964 0.388379
R22721 vdd.n2059 vdd.n2058 0.388379
R22722 vdd.n2025 vdd.n2023 0.388379
R22723 vdd.n19 vdd.n17 0.387128
R22724 vdd.n24 vdd.n22 0.387128
R22725 vdd.n6 vdd.n4 0.358259
R22726 vdd.n13 vdd.n11 0.358259
R22727 vdd.n276 vdd.n274 0.358259
R22728 vdd.n278 vdd.n276 0.358259
R22729 vdd.n280 vdd.n278 0.358259
R22730 vdd.n282 vdd.n280 0.358259
R22731 vdd.n284 vdd.n282 0.358259
R22732 vdd.n286 vdd.n284 0.358259
R22733 vdd.n288 vdd.n286 0.358259
R22734 vdd.n290 vdd.n288 0.358259
R22735 vdd.n332 vdd.n290 0.358259
R22736 vdd.n174 vdd.n172 0.358259
R22737 vdd.n176 vdd.n174 0.358259
R22738 vdd.n178 vdd.n176 0.358259
R22739 vdd.n180 vdd.n178 0.358259
R22740 vdd.n182 vdd.n180 0.358259
R22741 vdd.n184 vdd.n182 0.358259
R22742 vdd.n186 vdd.n184 0.358259
R22743 vdd.n188 vdd.n186 0.358259
R22744 vdd.n230 vdd.n188 0.358259
R22745 vdd.n73 vdd.n71 0.358259
R22746 vdd.n75 vdd.n73 0.358259
R22747 vdd.n77 vdd.n75 0.358259
R22748 vdd.n79 vdd.n77 0.358259
R22749 vdd.n81 vdd.n79 0.358259
R22750 vdd.n83 vdd.n81 0.358259
R22751 vdd.n85 vdd.n83 0.358259
R22752 vdd.n87 vdd.n85 0.358259
R22753 vdd.n129 vdd.n87 0.358259
R22754 vdd.n2265 vdd.n2223 0.358259
R22755 vdd.n2223 vdd.n2221 0.358259
R22756 vdd.n2221 vdd.n2219 0.358259
R22757 vdd.n2219 vdd.n2217 0.358259
R22758 vdd.n2217 vdd.n2215 0.358259
R22759 vdd.n2215 vdd.n2213 0.358259
R22760 vdd.n2213 vdd.n2211 0.358259
R22761 vdd.n2211 vdd.n2209 0.358259
R22762 vdd.n2209 vdd.n2207 0.358259
R22763 vdd.n2163 vdd.n2121 0.358259
R22764 vdd.n2121 vdd.n2119 0.358259
R22765 vdd.n2119 vdd.n2117 0.358259
R22766 vdd.n2117 vdd.n2115 0.358259
R22767 vdd.n2115 vdd.n2113 0.358259
R22768 vdd.n2113 vdd.n2111 0.358259
R22769 vdd.n2111 vdd.n2109 0.358259
R22770 vdd.n2109 vdd.n2107 0.358259
R22771 vdd.n2107 vdd.n2105 0.358259
R22772 vdd.n2062 vdd.n2020 0.358259
R22773 vdd.n2020 vdd.n2018 0.358259
R22774 vdd.n2018 vdd.n2016 0.358259
R22775 vdd.n2016 vdd.n2014 0.358259
R22776 vdd.n2014 vdd.n2012 0.358259
R22777 vdd.n2012 vdd.n2010 0.358259
R22778 vdd.n2010 vdd.n2008 0.358259
R22779 vdd.n2008 vdd.n2006 0.358259
R22780 vdd.n2006 vdd.n2004 0.358259
R22781 vdd.n2549 vdd.t289 0.340595
R22782 vdd.n1052 vdd.t247 0.340595
R22783 vdd.n3131 vdd.t236 0.340595
R22784 vdd.n877 vdd.t266 0.340595
R22785 vdd.n14 vdd.n6 0.334552
R22786 vdd.n14 vdd.n13 0.334552
R22787 vdd.n27 vdd.n19 0.21707
R22788 vdd.n27 vdd.n24 0.21707
R22789 vdd.n330 vdd.n292 0.155672
R22790 vdd.n322 vdd.n292 0.155672
R22791 vdd.n322 vdd.n321 0.155672
R22792 vdd.n321 vdd.n297 0.155672
R22793 vdd.n314 vdd.n297 0.155672
R22794 vdd.n314 vdd.n313 0.155672
R22795 vdd.n313 vdd.n301 0.155672
R22796 vdd.n306 vdd.n301 0.155672
R22797 vdd.n271 vdd.n233 0.155672
R22798 vdd.n263 vdd.n233 0.155672
R22799 vdd.n263 vdd.n262 0.155672
R22800 vdd.n262 vdd.n238 0.155672
R22801 vdd.n255 vdd.n238 0.155672
R22802 vdd.n255 vdd.n254 0.155672
R22803 vdd.n254 vdd.n242 0.155672
R22804 vdd.n247 vdd.n242 0.155672
R22805 vdd.n228 vdd.n190 0.155672
R22806 vdd.n220 vdd.n190 0.155672
R22807 vdd.n220 vdd.n219 0.155672
R22808 vdd.n219 vdd.n195 0.155672
R22809 vdd.n212 vdd.n195 0.155672
R22810 vdd.n212 vdd.n211 0.155672
R22811 vdd.n211 vdd.n199 0.155672
R22812 vdd.n204 vdd.n199 0.155672
R22813 vdd.n169 vdd.n131 0.155672
R22814 vdd.n161 vdd.n131 0.155672
R22815 vdd.n161 vdd.n160 0.155672
R22816 vdd.n160 vdd.n136 0.155672
R22817 vdd.n153 vdd.n136 0.155672
R22818 vdd.n153 vdd.n152 0.155672
R22819 vdd.n152 vdd.n140 0.155672
R22820 vdd.n145 vdd.n140 0.155672
R22821 vdd.n127 vdd.n89 0.155672
R22822 vdd.n119 vdd.n89 0.155672
R22823 vdd.n119 vdd.n118 0.155672
R22824 vdd.n118 vdd.n94 0.155672
R22825 vdd.n111 vdd.n94 0.155672
R22826 vdd.n111 vdd.n110 0.155672
R22827 vdd.n110 vdd.n98 0.155672
R22828 vdd.n103 vdd.n98 0.155672
R22829 vdd.n68 vdd.n30 0.155672
R22830 vdd.n60 vdd.n30 0.155672
R22831 vdd.n60 vdd.n59 0.155672
R22832 vdd.n59 vdd.n35 0.155672
R22833 vdd.n52 vdd.n35 0.155672
R22834 vdd.n52 vdd.n51 0.155672
R22835 vdd.n51 vdd.n39 0.155672
R22836 vdd.n44 vdd.n39 0.155672
R22837 vdd.n2204 vdd.n2166 0.155672
R22838 vdd.n2196 vdd.n2166 0.155672
R22839 vdd.n2196 vdd.n2195 0.155672
R22840 vdd.n2195 vdd.n2171 0.155672
R22841 vdd.n2188 vdd.n2171 0.155672
R22842 vdd.n2188 vdd.n2187 0.155672
R22843 vdd.n2187 vdd.n2175 0.155672
R22844 vdd.n2180 vdd.n2175 0.155672
R22845 vdd.n2263 vdd.n2225 0.155672
R22846 vdd.n2255 vdd.n2225 0.155672
R22847 vdd.n2255 vdd.n2254 0.155672
R22848 vdd.n2254 vdd.n2230 0.155672
R22849 vdd.n2247 vdd.n2230 0.155672
R22850 vdd.n2247 vdd.n2246 0.155672
R22851 vdd.n2246 vdd.n2234 0.155672
R22852 vdd.n2239 vdd.n2234 0.155672
R22853 vdd.n2102 vdd.n2064 0.155672
R22854 vdd.n2094 vdd.n2064 0.155672
R22855 vdd.n2094 vdd.n2093 0.155672
R22856 vdd.n2093 vdd.n2069 0.155672
R22857 vdd.n2086 vdd.n2069 0.155672
R22858 vdd.n2086 vdd.n2085 0.155672
R22859 vdd.n2085 vdd.n2073 0.155672
R22860 vdd.n2078 vdd.n2073 0.155672
R22861 vdd.n2161 vdd.n2123 0.155672
R22862 vdd.n2153 vdd.n2123 0.155672
R22863 vdd.n2153 vdd.n2152 0.155672
R22864 vdd.n2152 vdd.n2128 0.155672
R22865 vdd.n2145 vdd.n2128 0.155672
R22866 vdd.n2145 vdd.n2144 0.155672
R22867 vdd.n2144 vdd.n2132 0.155672
R22868 vdd.n2137 vdd.n2132 0.155672
R22869 vdd.n2001 vdd.n1963 0.155672
R22870 vdd.n1993 vdd.n1963 0.155672
R22871 vdd.n1993 vdd.n1992 0.155672
R22872 vdd.n1992 vdd.n1968 0.155672
R22873 vdd.n1985 vdd.n1968 0.155672
R22874 vdd.n1985 vdd.n1984 0.155672
R22875 vdd.n1984 vdd.n1972 0.155672
R22876 vdd.n1977 vdd.n1972 0.155672
R22877 vdd.n2060 vdd.n2022 0.155672
R22878 vdd.n2052 vdd.n2022 0.155672
R22879 vdd.n2052 vdd.n2051 0.155672
R22880 vdd.n2051 vdd.n2027 0.155672
R22881 vdd.n2044 vdd.n2027 0.155672
R22882 vdd.n2044 vdd.n2043 0.155672
R22883 vdd.n2043 vdd.n2031 0.155672
R22884 vdd.n2036 vdd.n2031 0.155672
R22885 vdd.n1186 vdd.n1178 0.152939
R22886 vdd.n1190 vdd.n1186 0.152939
R22887 vdd.n1191 vdd.n1190 0.152939
R22888 vdd.n1192 vdd.n1191 0.152939
R22889 vdd.n1193 vdd.n1192 0.152939
R22890 vdd.n1197 vdd.n1193 0.152939
R22891 vdd.n1198 vdd.n1197 0.152939
R22892 vdd.n1199 vdd.n1198 0.152939
R22893 vdd.n1200 vdd.n1199 0.152939
R22894 vdd.n1204 vdd.n1200 0.152939
R22895 vdd.n1205 vdd.n1204 0.152939
R22896 vdd.n1206 vdd.n1205 0.152939
R22897 vdd.n2438 vdd.n1206 0.152939
R22898 vdd.n2438 vdd.n2437 0.152939
R22899 vdd.n2437 vdd.n2436 0.152939
R22900 vdd.n2436 vdd.n1212 0.152939
R22901 vdd.n1217 vdd.n1212 0.152939
R22902 vdd.n1218 vdd.n1217 0.152939
R22903 vdd.n1219 vdd.n1218 0.152939
R22904 vdd.n1223 vdd.n1219 0.152939
R22905 vdd.n1224 vdd.n1223 0.152939
R22906 vdd.n1225 vdd.n1224 0.152939
R22907 vdd.n1226 vdd.n1225 0.152939
R22908 vdd.n1230 vdd.n1226 0.152939
R22909 vdd.n1231 vdd.n1230 0.152939
R22910 vdd.n1232 vdd.n1231 0.152939
R22911 vdd.n1233 vdd.n1232 0.152939
R22912 vdd.n1237 vdd.n1233 0.152939
R22913 vdd.n1238 vdd.n1237 0.152939
R22914 vdd.n1239 vdd.n1238 0.152939
R22915 vdd.n1240 vdd.n1239 0.152939
R22916 vdd.n1244 vdd.n1240 0.152939
R22917 vdd.n1245 vdd.n1244 0.152939
R22918 vdd.n1246 vdd.n1245 0.152939
R22919 vdd.n2399 vdd.n1246 0.152939
R22920 vdd.n2399 vdd.n2398 0.152939
R22921 vdd.n2398 vdd.n2397 0.152939
R22922 vdd.n2397 vdd.n1252 0.152939
R22923 vdd.n1257 vdd.n1252 0.152939
R22924 vdd.n1258 vdd.n1257 0.152939
R22925 vdd.n1259 vdd.n1258 0.152939
R22926 vdd.n1263 vdd.n1259 0.152939
R22927 vdd.n1264 vdd.n1263 0.152939
R22928 vdd.n1265 vdd.n1264 0.152939
R22929 vdd.n1266 vdd.n1265 0.152939
R22930 vdd.n1270 vdd.n1266 0.152939
R22931 vdd.n1271 vdd.n1270 0.152939
R22932 vdd.n1272 vdd.n1271 0.152939
R22933 vdd.n1273 vdd.n1272 0.152939
R22934 vdd.n1277 vdd.n1273 0.152939
R22935 vdd.n1278 vdd.n1277 0.152939
R22936 vdd.n2473 vdd.n1181 0.152939
R22937 vdd.n2269 vdd.n1578 0.152939
R22938 vdd.n2284 vdd.n1578 0.152939
R22939 vdd.n2285 vdd.n2284 0.152939
R22940 vdd.n2286 vdd.n2285 0.152939
R22941 vdd.n2286 vdd.n1567 0.152939
R22942 vdd.n2301 vdd.n1567 0.152939
R22943 vdd.n2302 vdd.n2301 0.152939
R22944 vdd.n2303 vdd.n2302 0.152939
R22945 vdd.n2303 vdd.n1556 0.152939
R22946 vdd.n2317 vdd.n1556 0.152939
R22947 vdd.n2318 vdd.n2317 0.152939
R22948 vdd.n2319 vdd.n2318 0.152939
R22949 vdd.n2319 vdd.n1544 0.152939
R22950 vdd.n2334 vdd.n1544 0.152939
R22951 vdd.n2335 vdd.n2334 0.152939
R22952 vdd.n2336 vdd.n2335 0.152939
R22953 vdd.n2336 vdd.n1532 0.152939
R22954 vdd.n2353 vdd.n1532 0.152939
R22955 vdd.n2354 vdd.n2353 0.152939
R22956 vdd.n2355 vdd.n2354 0.152939
R22957 vdd.n735 vdd.n730 0.152939
R22958 vdd.n736 vdd.n735 0.152939
R22959 vdd.n737 vdd.n736 0.152939
R22960 vdd.n738 vdd.n737 0.152939
R22961 vdd.n739 vdd.n738 0.152939
R22962 vdd.n740 vdd.n739 0.152939
R22963 vdd.n741 vdd.n740 0.152939
R22964 vdd.n742 vdd.n741 0.152939
R22965 vdd.n743 vdd.n742 0.152939
R22966 vdd.n744 vdd.n743 0.152939
R22967 vdd.n745 vdd.n744 0.152939
R22968 vdd.n746 vdd.n745 0.152939
R22969 vdd.n3455 vdd.n746 0.152939
R22970 vdd.n3455 vdd.n3454 0.152939
R22971 vdd.n3454 vdd.n3453 0.152939
R22972 vdd.n3453 vdd.n748 0.152939
R22973 vdd.n749 vdd.n748 0.152939
R22974 vdd.n750 vdd.n749 0.152939
R22975 vdd.n751 vdd.n750 0.152939
R22976 vdd.n752 vdd.n751 0.152939
R22977 vdd.n753 vdd.n752 0.152939
R22978 vdd.n754 vdd.n753 0.152939
R22979 vdd.n755 vdd.n754 0.152939
R22980 vdd.n756 vdd.n755 0.152939
R22981 vdd.n757 vdd.n756 0.152939
R22982 vdd.n758 vdd.n757 0.152939
R22983 vdd.n759 vdd.n758 0.152939
R22984 vdd.n760 vdd.n759 0.152939
R22985 vdd.n761 vdd.n760 0.152939
R22986 vdd.n762 vdd.n761 0.152939
R22987 vdd.n763 vdd.n762 0.152939
R22988 vdd.n764 vdd.n763 0.152939
R22989 vdd.n765 vdd.n764 0.152939
R22990 vdd.n766 vdd.n765 0.152939
R22991 vdd.n3409 vdd.n766 0.152939
R22992 vdd.n3409 vdd.n3408 0.152939
R22993 vdd.n3408 vdd.n3407 0.152939
R22994 vdd.n3407 vdd.n770 0.152939
R22995 vdd.n771 vdd.n770 0.152939
R22996 vdd.n772 vdd.n771 0.152939
R22997 vdd.n773 vdd.n772 0.152939
R22998 vdd.n774 vdd.n773 0.152939
R22999 vdd.n775 vdd.n774 0.152939
R23000 vdd.n776 vdd.n775 0.152939
R23001 vdd.n777 vdd.n776 0.152939
R23002 vdd.n778 vdd.n777 0.152939
R23003 vdd.n779 vdd.n778 0.152939
R23004 vdd.n780 vdd.n779 0.152939
R23005 vdd.n781 vdd.n780 0.152939
R23006 vdd.n782 vdd.n781 0.152939
R23007 vdd.n783 vdd.n782 0.152939
R23008 vdd.n727 vdd.n726 0.152939
R23009 vdd.n3506 vdd.n682 0.152939
R23010 vdd.n3507 vdd.n3506 0.152939
R23011 vdd.n3508 vdd.n3507 0.152939
R23012 vdd.n3508 vdd.n670 0.152939
R23013 vdd.n3523 vdd.n670 0.152939
R23014 vdd.n3524 vdd.n3523 0.152939
R23015 vdd.n3525 vdd.n3524 0.152939
R23016 vdd.n3525 vdd.n659 0.152939
R23017 vdd.n3539 vdd.n659 0.152939
R23018 vdd.n3540 vdd.n3539 0.152939
R23019 vdd.n3541 vdd.n3540 0.152939
R23020 vdd.n3541 vdd.n647 0.152939
R23021 vdd.n3556 vdd.n647 0.152939
R23022 vdd.n3557 vdd.n3556 0.152939
R23023 vdd.n3558 vdd.n3557 0.152939
R23024 vdd.n3558 vdd.n636 0.152939
R23025 vdd.n3575 vdd.n636 0.152939
R23026 vdd.n3576 vdd.n3575 0.152939
R23027 vdd.n3577 vdd.n3576 0.152939
R23028 vdd.n3577 vdd.n334 0.152939
R23029 vdd.n3670 vdd.n335 0.152939
R23030 vdd.n346 vdd.n335 0.152939
R23031 vdd.n347 vdd.n346 0.152939
R23032 vdd.n348 vdd.n347 0.152939
R23033 vdd.n355 vdd.n348 0.152939
R23034 vdd.n356 vdd.n355 0.152939
R23035 vdd.n357 vdd.n356 0.152939
R23036 vdd.n358 vdd.n357 0.152939
R23037 vdd.n366 vdd.n358 0.152939
R23038 vdd.n367 vdd.n366 0.152939
R23039 vdd.n368 vdd.n367 0.152939
R23040 vdd.n369 vdd.n368 0.152939
R23041 vdd.n377 vdd.n369 0.152939
R23042 vdd.n378 vdd.n377 0.152939
R23043 vdd.n379 vdd.n378 0.152939
R23044 vdd.n380 vdd.n379 0.152939
R23045 vdd.n388 vdd.n380 0.152939
R23046 vdd.n389 vdd.n388 0.152939
R23047 vdd.n390 vdd.n389 0.152939
R23048 vdd.n391 vdd.n390 0.152939
R23049 vdd.n464 vdd.n463 0.152939
R23050 vdd.n470 vdd.n463 0.152939
R23051 vdd.n471 vdd.n470 0.152939
R23052 vdd.n472 vdd.n471 0.152939
R23053 vdd.n472 vdd.n461 0.152939
R23054 vdd.n480 vdd.n461 0.152939
R23055 vdd.n481 vdd.n480 0.152939
R23056 vdd.n482 vdd.n481 0.152939
R23057 vdd.n482 vdd.n459 0.152939
R23058 vdd.n490 vdd.n459 0.152939
R23059 vdd.n491 vdd.n490 0.152939
R23060 vdd.n492 vdd.n491 0.152939
R23061 vdd.n492 vdd.n457 0.152939
R23062 vdd.n500 vdd.n457 0.152939
R23063 vdd.n501 vdd.n500 0.152939
R23064 vdd.n502 vdd.n501 0.152939
R23065 vdd.n502 vdd.n455 0.152939
R23066 vdd.n510 vdd.n455 0.152939
R23067 vdd.n511 vdd.n510 0.152939
R23068 vdd.n512 vdd.n511 0.152939
R23069 vdd.n512 vdd.n451 0.152939
R23070 vdd.n520 vdd.n451 0.152939
R23071 vdd.n521 vdd.n520 0.152939
R23072 vdd.n522 vdd.n521 0.152939
R23073 vdd.n522 vdd.n449 0.152939
R23074 vdd.n530 vdd.n449 0.152939
R23075 vdd.n531 vdd.n530 0.152939
R23076 vdd.n532 vdd.n531 0.152939
R23077 vdd.n532 vdd.n447 0.152939
R23078 vdd.n540 vdd.n447 0.152939
R23079 vdd.n541 vdd.n540 0.152939
R23080 vdd.n542 vdd.n541 0.152939
R23081 vdd.n542 vdd.n445 0.152939
R23082 vdd.n550 vdd.n445 0.152939
R23083 vdd.n551 vdd.n550 0.152939
R23084 vdd.n552 vdd.n551 0.152939
R23085 vdd.n552 vdd.n443 0.152939
R23086 vdd.n560 vdd.n443 0.152939
R23087 vdd.n561 vdd.n560 0.152939
R23088 vdd.n562 vdd.n561 0.152939
R23089 vdd.n562 vdd.n439 0.152939
R23090 vdd.n570 vdd.n439 0.152939
R23091 vdd.n571 vdd.n570 0.152939
R23092 vdd.n572 vdd.n571 0.152939
R23093 vdd.n572 vdd.n437 0.152939
R23094 vdd.n580 vdd.n437 0.152939
R23095 vdd.n581 vdd.n580 0.152939
R23096 vdd.n582 vdd.n581 0.152939
R23097 vdd.n582 vdd.n435 0.152939
R23098 vdd.n590 vdd.n435 0.152939
R23099 vdd.n591 vdd.n590 0.152939
R23100 vdd.n592 vdd.n591 0.152939
R23101 vdd.n592 vdd.n433 0.152939
R23102 vdd.n600 vdd.n433 0.152939
R23103 vdd.n601 vdd.n600 0.152939
R23104 vdd.n602 vdd.n601 0.152939
R23105 vdd.n602 vdd.n431 0.152939
R23106 vdd.n610 vdd.n431 0.152939
R23107 vdd.n611 vdd.n610 0.152939
R23108 vdd.n612 vdd.n611 0.152939
R23109 vdd.n612 vdd.n429 0.152939
R23110 vdd.n619 vdd.n429 0.152939
R23111 vdd.n3622 vdd.n619 0.152939
R23112 vdd.n3500 vdd.n3499 0.152939
R23113 vdd.n3500 vdd.n675 0.152939
R23114 vdd.n3514 vdd.n675 0.152939
R23115 vdd.n3515 vdd.n3514 0.152939
R23116 vdd.n3516 vdd.n3515 0.152939
R23117 vdd.n3516 vdd.n665 0.152939
R23118 vdd.n3531 vdd.n665 0.152939
R23119 vdd.n3532 vdd.n3531 0.152939
R23120 vdd.n3533 vdd.n3532 0.152939
R23121 vdd.n3533 vdd.n652 0.152939
R23122 vdd.n3547 vdd.n652 0.152939
R23123 vdd.n3548 vdd.n3547 0.152939
R23124 vdd.n3549 vdd.n3548 0.152939
R23125 vdd.n3549 vdd.n641 0.152939
R23126 vdd.n3564 vdd.n641 0.152939
R23127 vdd.n3565 vdd.n3564 0.152939
R23128 vdd.n3566 vdd.n3565 0.152939
R23129 vdd.n3568 vdd.n3566 0.152939
R23130 vdd.n3568 vdd.n3567 0.152939
R23131 vdd.n3567 vdd.n630 0.152939
R23132 vdd.n3585 vdd.n630 0.152939
R23133 vdd.n3586 vdd.n3585 0.152939
R23134 vdd.n3587 vdd.n3586 0.152939
R23135 vdd.n3587 vdd.n628 0.152939
R23136 vdd.n3592 vdd.n628 0.152939
R23137 vdd.n3593 vdd.n3592 0.152939
R23138 vdd.n3594 vdd.n3593 0.152939
R23139 vdd.n3594 vdd.n626 0.152939
R23140 vdd.n3599 vdd.n626 0.152939
R23141 vdd.n3600 vdd.n3599 0.152939
R23142 vdd.n3601 vdd.n3600 0.152939
R23143 vdd.n3601 vdd.n624 0.152939
R23144 vdd.n3607 vdd.n624 0.152939
R23145 vdd.n3608 vdd.n3607 0.152939
R23146 vdd.n3609 vdd.n3608 0.152939
R23147 vdd.n3609 vdd.n622 0.152939
R23148 vdd.n3614 vdd.n622 0.152939
R23149 vdd.n3615 vdd.n3614 0.152939
R23150 vdd.n3616 vdd.n3615 0.152939
R23151 vdd.n3616 vdd.n620 0.152939
R23152 vdd.n3621 vdd.n620 0.152939
R23153 vdd.n3498 vdd.n687 0.152939
R23154 vdd.n2366 vdd.n1517 0.152939
R23155 vdd.n1885 vdd.n1641 0.152939
R23156 vdd.n1886 vdd.n1885 0.152939
R23157 vdd.n1887 vdd.n1886 0.152939
R23158 vdd.n1887 vdd.n1629 0.152939
R23159 vdd.n1902 vdd.n1629 0.152939
R23160 vdd.n1903 vdd.n1902 0.152939
R23161 vdd.n1904 vdd.n1903 0.152939
R23162 vdd.n1904 vdd.n1619 0.152939
R23163 vdd.n1919 vdd.n1619 0.152939
R23164 vdd.n1920 vdd.n1919 0.152939
R23165 vdd.n1921 vdd.n1920 0.152939
R23166 vdd.n1921 vdd.n1606 0.152939
R23167 vdd.n1935 vdd.n1606 0.152939
R23168 vdd.n1936 vdd.n1935 0.152939
R23169 vdd.n1937 vdd.n1936 0.152939
R23170 vdd.n1937 vdd.n1595 0.152939
R23171 vdd.n1952 vdd.n1595 0.152939
R23172 vdd.n1953 vdd.n1952 0.152939
R23173 vdd.n1954 vdd.n1953 0.152939
R23174 vdd.n1954 vdd.n1584 0.152939
R23175 vdd.n2275 vdd.n1584 0.152939
R23176 vdd.n2276 vdd.n2275 0.152939
R23177 vdd.n2277 vdd.n2276 0.152939
R23178 vdd.n2277 vdd.n1572 0.152939
R23179 vdd.n2292 vdd.n1572 0.152939
R23180 vdd.n2293 vdd.n2292 0.152939
R23181 vdd.n2294 vdd.n2293 0.152939
R23182 vdd.n2294 vdd.n1562 0.152939
R23183 vdd.n2309 vdd.n1562 0.152939
R23184 vdd.n2310 vdd.n2309 0.152939
R23185 vdd.n2311 vdd.n2310 0.152939
R23186 vdd.n2311 vdd.n1549 0.152939
R23187 vdd.n2325 vdd.n1549 0.152939
R23188 vdd.n2326 vdd.n2325 0.152939
R23189 vdd.n2327 vdd.n2326 0.152939
R23190 vdd.n2327 vdd.n1539 0.152939
R23191 vdd.n2342 vdd.n1539 0.152939
R23192 vdd.n2343 vdd.n2342 0.152939
R23193 vdd.n2346 vdd.n2343 0.152939
R23194 vdd.n2346 vdd.n2345 0.152939
R23195 vdd.n2345 vdd.n2344 0.152939
R23196 vdd.n1877 vdd.n1646 0.152939
R23197 vdd.n1870 vdd.n1646 0.152939
R23198 vdd.n1870 vdd.n1869 0.152939
R23199 vdd.n1869 vdd.n1868 0.152939
R23200 vdd.n1868 vdd.n1683 0.152939
R23201 vdd.n1864 vdd.n1683 0.152939
R23202 vdd.n1864 vdd.n1863 0.152939
R23203 vdd.n1863 vdd.n1862 0.152939
R23204 vdd.n1862 vdd.n1689 0.152939
R23205 vdd.n1858 vdd.n1689 0.152939
R23206 vdd.n1858 vdd.n1857 0.152939
R23207 vdd.n1857 vdd.n1856 0.152939
R23208 vdd.n1856 vdd.n1695 0.152939
R23209 vdd.n1852 vdd.n1695 0.152939
R23210 vdd.n1852 vdd.n1851 0.152939
R23211 vdd.n1851 vdd.n1850 0.152939
R23212 vdd.n1850 vdd.n1701 0.152939
R23213 vdd.n1846 vdd.n1701 0.152939
R23214 vdd.n1846 vdd.n1845 0.152939
R23215 vdd.n1845 vdd.n1844 0.152939
R23216 vdd.n1844 vdd.n1709 0.152939
R23217 vdd.n1840 vdd.n1709 0.152939
R23218 vdd.n1840 vdd.n1839 0.152939
R23219 vdd.n1839 vdd.n1838 0.152939
R23220 vdd.n1838 vdd.n1715 0.152939
R23221 vdd.n1834 vdd.n1715 0.152939
R23222 vdd.n1834 vdd.n1833 0.152939
R23223 vdd.n1833 vdd.n1832 0.152939
R23224 vdd.n1832 vdd.n1721 0.152939
R23225 vdd.n1828 vdd.n1721 0.152939
R23226 vdd.n1828 vdd.n1827 0.152939
R23227 vdd.n1827 vdd.n1826 0.152939
R23228 vdd.n1826 vdd.n1727 0.152939
R23229 vdd.n1822 vdd.n1727 0.152939
R23230 vdd.n1822 vdd.n1821 0.152939
R23231 vdd.n1821 vdd.n1820 0.152939
R23232 vdd.n1820 vdd.n1733 0.152939
R23233 vdd.n1816 vdd.n1733 0.152939
R23234 vdd.n1816 vdd.n1815 0.152939
R23235 vdd.n1815 vdd.n1814 0.152939
R23236 vdd.n1814 vdd.n1739 0.152939
R23237 vdd.n1807 vdd.n1739 0.152939
R23238 vdd.n1807 vdd.n1806 0.152939
R23239 vdd.n1806 vdd.n1805 0.152939
R23240 vdd.n1805 vdd.n1744 0.152939
R23241 vdd.n1801 vdd.n1744 0.152939
R23242 vdd.n1801 vdd.n1800 0.152939
R23243 vdd.n1800 vdd.n1799 0.152939
R23244 vdd.n1799 vdd.n1750 0.152939
R23245 vdd.n1795 vdd.n1750 0.152939
R23246 vdd.n1795 vdd.n1794 0.152939
R23247 vdd.n1794 vdd.n1793 0.152939
R23248 vdd.n1793 vdd.n1756 0.152939
R23249 vdd.n1789 vdd.n1756 0.152939
R23250 vdd.n1789 vdd.n1788 0.152939
R23251 vdd.n1788 vdd.n1787 0.152939
R23252 vdd.n1787 vdd.n1762 0.152939
R23253 vdd.n1783 vdd.n1762 0.152939
R23254 vdd.n1783 vdd.n1782 0.152939
R23255 vdd.n1782 vdd.n1781 0.152939
R23256 vdd.n1781 vdd.n1768 0.152939
R23257 vdd.n1777 vdd.n1768 0.152939
R23258 vdd.n1777 vdd.n1776 0.152939
R23259 vdd.n1879 vdd.n1878 0.152939
R23260 vdd.n1879 vdd.n1635 0.152939
R23261 vdd.n1894 vdd.n1635 0.152939
R23262 vdd.n1895 vdd.n1894 0.152939
R23263 vdd.n1896 vdd.n1895 0.152939
R23264 vdd.n1896 vdd.n1624 0.152939
R23265 vdd.n1911 vdd.n1624 0.152939
R23266 vdd.n1912 vdd.n1911 0.152939
R23267 vdd.n1913 vdd.n1912 0.152939
R23268 vdd.n1913 vdd.n1613 0.152939
R23269 vdd.n1927 vdd.n1613 0.152939
R23270 vdd.n1928 vdd.n1927 0.152939
R23271 vdd.n1929 vdd.n1928 0.152939
R23272 vdd.n1929 vdd.n1601 0.152939
R23273 vdd.n1944 vdd.n1601 0.152939
R23274 vdd.n1945 vdd.n1944 0.152939
R23275 vdd.n1946 vdd.n1945 0.152939
R23276 vdd.n1946 vdd.n1590 0.152939
R23277 vdd.n1960 vdd.n1590 0.152939
R23278 vdd.n1961 vdd.n1960 0.152939
R23279 vdd.n1882 vdd.t224 0.113865
R23280 vdd.t173 vdd.n386 0.113865
R23281 vdd.n2474 vdd.n2473 0.110256
R23282 vdd.n3488 vdd.n727 0.110256
R23283 vdd.n3365 vdd.n687 0.110256
R23284 vdd.n2367 vdd.n2366 0.110256
R23285 vdd.n2269 vdd.n2268 0.0695946
R23286 vdd.n3671 vdd.n334 0.0695946
R23287 vdd.n3671 vdd.n3670 0.0695946
R23288 vdd.n2268 vdd.n1961 0.0695946
R23289 vdd.n2474 vdd.n1178 0.0431829
R23290 vdd.n2367 vdd.n1278 0.0431829
R23291 vdd.n3488 vdd.n730 0.0431829
R23292 vdd.n3365 vdd.n783 0.0431829
R23293 vdd vdd.n28 0.00833333
R23294 a_n2804_13878.n2 a_n2804_13878.n0 98.9633
R23295 a_n2804_13878.n5 a_n2804_13878.n3 98.7517
R23296 a_n2804_13878.n25 a_n2804_13878.n24 98.6055
R23297 a_n2804_13878.n27 a_n2804_13878.n26 98.6055
R23298 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R23299 a_n2804_13878.n13 a_n2804_13878.n12 98.6055
R23300 a_n2804_13878.n11 a_n2804_13878.n10 98.6055
R23301 a_n2804_13878.n9 a_n2804_13878.n8 98.6055
R23302 a_n2804_13878.n7 a_n2804_13878.n6 98.6055
R23303 a_n2804_13878.n5 a_n2804_13878.n4 98.6055
R23304 a_n2804_13878.n29 a_n2804_13878.n28 98.6054
R23305 a_n2804_13878.n23 a_n2804_13878.n22 98.6054
R23306 a_n2804_13878.n15 a_n2804_13878.t1 74.6477
R23307 a_n2804_13878.n20 a_n2804_13878.t2 74.2899
R23308 a_n2804_13878.n17 a_n2804_13878.t3 74.2899
R23309 a_n2804_13878.n16 a_n2804_13878.t0 74.2899
R23310 a_n2804_13878.n19 a_n2804_13878.n18 70.6783
R23311 a_n2804_13878.n15 a_n2804_13878.n14 70.6783
R23312 a_n2804_13878.n21 a_n2804_13878.n13 15.7159
R23313 a_n2804_13878.n23 a_n2804_13878.n21 12.6495
R23314 a_n2804_13878.n21 a_n2804_13878.n20 8.38735
R23315 a_n2804_13878.n22 a_n2804_13878.t15 3.61217
R23316 a_n2804_13878.n22 a_n2804_13878.t24 3.61217
R23317 a_n2804_13878.n24 a_n2804_13878.t28 3.61217
R23318 a_n2804_13878.n24 a_n2804_13878.t14 3.61217
R23319 a_n2804_13878.n26 a_n2804_13878.t18 3.61217
R23320 a_n2804_13878.n26 a_n2804_13878.t19 3.61217
R23321 a_n2804_13878.n1 a_n2804_13878.t8 3.61217
R23322 a_n2804_13878.n1 a_n2804_13878.t20 3.61217
R23323 a_n2804_13878.n0 a_n2804_13878.t25 3.61217
R23324 a_n2804_13878.n0 a_n2804_13878.t31 3.61217
R23325 a_n2804_13878.n18 a_n2804_13878.t6 3.61217
R23326 a_n2804_13878.n18 a_n2804_13878.t7 3.61217
R23327 a_n2804_13878.n14 a_n2804_13878.t4 3.61217
R23328 a_n2804_13878.n14 a_n2804_13878.t5 3.61217
R23329 a_n2804_13878.n12 a_n2804_13878.t21 3.61217
R23330 a_n2804_13878.n12 a_n2804_13878.t9 3.61217
R23331 a_n2804_13878.n10 a_n2804_13878.t26 3.61217
R23332 a_n2804_13878.n10 a_n2804_13878.t11 3.61217
R23333 a_n2804_13878.n8 a_n2804_13878.t10 3.61217
R23334 a_n2804_13878.n8 a_n2804_13878.t13 3.61217
R23335 a_n2804_13878.n6 a_n2804_13878.t23 3.61217
R23336 a_n2804_13878.n6 a_n2804_13878.t16 3.61217
R23337 a_n2804_13878.n4 a_n2804_13878.t27 3.61217
R23338 a_n2804_13878.n4 a_n2804_13878.t17 3.61217
R23339 a_n2804_13878.n3 a_n2804_13878.t12 3.61217
R23340 a_n2804_13878.n3 a_n2804_13878.t22 3.61217
R23341 a_n2804_13878.n29 a_n2804_13878.t29 3.61217
R23342 a_n2804_13878.t30 a_n2804_13878.n29 3.61217
R23343 a_n2804_13878.n16 a_n2804_13878.n15 0.358259
R23344 a_n2804_13878.n19 a_n2804_13878.n17 0.358259
R23345 a_n2804_13878.n20 a_n2804_13878.n19 0.358259
R23346 a_n2804_13878.n28 a_n2804_13878.n2 0.358259
R23347 a_n2804_13878.n28 a_n2804_13878.n27 0.358259
R23348 a_n2804_13878.n27 a_n2804_13878.n25 0.358259
R23349 a_n2804_13878.n25 a_n2804_13878.n23 0.358259
R23350 a_n2804_13878.n7 a_n2804_13878.n5 0.146627
R23351 a_n2804_13878.n9 a_n2804_13878.n7 0.146627
R23352 a_n2804_13878.n11 a_n2804_13878.n9 0.146627
R23353 a_n2804_13878.n13 a_n2804_13878.n11 0.146627
R23354 a_n2804_13878.n17 a_n2804_13878.n16 0.101793
R23355 a_n2982_8322.n12 a_n2982_8322.t27 74.6477
R23356 a_n2982_8322.n1 a_n2982_8322.t6 74.6477
R23357 a_n2982_8322.n28 a_n2982_8322.t21 74.6474
R23358 a_n2982_8322.n20 a_n2982_8322.t1 74.2899
R23359 a_n2982_8322.n13 a_n2982_8322.t25 74.2899
R23360 a_n2982_8322.n14 a_n2982_8322.t28 74.2899
R23361 a_n2982_8322.n17 a_n2982_8322.t29 74.2899
R23362 a_n2982_8322.n10 a_n2982_8322.t0 74.2899
R23363 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R23364 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R23365 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R23366 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R23367 a_n2982_8322.n12 a_n2982_8322.n11 70.6783
R23368 a_n2982_8322.n16 a_n2982_8322.n15 70.6783
R23369 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R23370 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R23371 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R23372 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R23373 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R23374 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R23375 a_n2982_8322.n18 a_n2982_8322.n10 24.9022
R23376 a_n2982_8322.n19 a_n2982_8322.t32 9.69161
R23377 a_n2982_8322.n18 a_n2982_8322.n17 8.38735
R23378 a_n2982_8322.n20 a_n2982_8322.n19 6.90998
R23379 a_n2982_8322.n19 a_n2982_8322.n18 5.3452
R23380 a_n2982_8322.n27 a_n2982_8322.t14 3.61217
R23381 a_n2982_8322.n27 a_n2982_8322.t10 3.61217
R23382 a_n2982_8322.n25 a_n2982_8322.t20 3.61217
R23383 a_n2982_8322.n25 a_n2982_8322.t8 3.61217
R23384 a_n2982_8322.n23 a_n2982_8322.t5 3.61217
R23385 a_n2982_8322.n23 a_n2982_8322.t4 3.61217
R23386 a_n2982_8322.n21 a_n2982_8322.t18 3.61217
R23387 a_n2982_8322.n21 a_n2982_8322.t17 3.61217
R23388 a_n2982_8322.n11 a_n2982_8322.t31 3.61217
R23389 a_n2982_8322.n11 a_n2982_8322.t30 3.61217
R23390 a_n2982_8322.n15 a_n2982_8322.t26 3.61217
R23391 a_n2982_8322.n15 a_n2982_8322.t24 3.61217
R23392 a_n2982_8322.n0 a_n2982_8322.t19 3.61217
R23393 a_n2982_8322.n0 a_n2982_8322.t15 3.61217
R23394 a_n2982_8322.n2 a_n2982_8322.t22 3.61217
R23395 a_n2982_8322.n2 a_n2982_8322.t12 3.61217
R23396 a_n2982_8322.n4 a_n2982_8322.t3 3.61217
R23397 a_n2982_8322.n4 a_n2982_8322.t2 3.61217
R23398 a_n2982_8322.n6 a_n2982_8322.t16 3.61217
R23399 a_n2982_8322.n6 a_n2982_8322.t9 3.61217
R23400 a_n2982_8322.n8 a_n2982_8322.t13 3.61217
R23401 a_n2982_8322.n8 a_n2982_8322.t11 3.61217
R23402 a_n2982_8322.n30 a_n2982_8322.t7 3.61217
R23403 a_n2982_8322.t23 a_n2982_8322.n30 3.61217
R23404 a_n2982_8322.n17 a_n2982_8322.n16 0.358259
R23405 a_n2982_8322.n16 a_n2982_8322.n14 0.358259
R23406 a_n2982_8322.n13 a_n2982_8322.n12 0.358259
R23407 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R23408 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R23409 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R23410 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R23411 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R23412 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R23413 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R23414 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R23415 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R23416 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R23417 a_n2982_8322.n14 a_n2982_8322.n13 0.101793
R23418 a_n2982_8322.t37 a_n2982_8322.t33 0.0788333
R23419 a_n2982_8322.t36 a_n2982_8322.t34 0.0788333
R23420 a_n2982_8322.t32 a_n2982_8322.t35 0.0788333
R23421 a_n2982_8322.t36 a_n2982_8322.t37 0.0318333
R23422 a_n2982_8322.t32 a_n2982_8322.t34 0.0318333
R23423 a_n2982_8322.t33 a_n2982_8322.t34 0.0318333
R23424 a_n2982_8322.t35 a_n2982_8322.t36 0.0318333
R23425 output.n41 output.n15 289.615
R23426 output.n72 output.n46 289.615
R23427 output.n104 output.n78 289.615
R23428 output.n136 output.n110 289.615
R23429 output.n77 output.n45 197.26
R23430 output.n77 output.n76 196.298
R23431 output.n109 output.n108 196.298
R23432 output.n141 output.n140 196.298
R23433 output.n42 output.n41 185
R23434 output.n40 output.n39 185
R23435 output.n19 output.n18 185
R23436 output.n34 output.n33 185
R23437 output.n32 output.n31 185
R23438 output.n23 output.n22 185
R23439 output.n26 output.n25 185
R23440 output.n73 output.n72 185
R23441 output.n71 output.n70 185
R23442 output.n50 output.n49 185
R23443 output.n65 output.n64 185
R23444 output.n63 output.n62 185
R23445 output.n54 output.n53 185
R23446 output.n57 output.n56 185
R23447 output.n105 output.n104 185
R23448 output.n103 output.n102 185
R23449 output.n82 output.n81 185
R23450 output.n97 output.n96 185
R23451 output.n95 output.n94 185
R23452 output.n86 output.n85 185
R23453 output.n89 output.n88 185
R23454 output.n137 output.n136 185
R23455 output.n135 output.n134 185
R23456 output.n114 output.n113 185
R23457 output.n129 output.n128 185
R23458 output.n127 output.n126 185
R23459 output.n118 output.n117 185
R23460 output.n121 output.n120 185
R23461 output.t1 output.n24 147.661
R23462 output.t0 output.n55 147.661
R23463 output.t2 output.n87 147.661
R23464 output.t19 output.n119 147.661
R23465 output.n41 output.n40 104.615
R23466 output.n40 output.n18 104.615
R23467 output.n33 output.n18 104.615
R23468 output.n33 output.n32 104.615
R23469 output.n32 output.n22 104.615
R23470 output.n25 output.n22 104.615
R23471 output.n72 output.n71 104.615
R23472 output.n71 output.n49 104.615
R23473 output.n64 output.n49 104.615
R23474 output.n64 output.n63 104.615
R23475 output.n63 output.n53 104.615
R23476 output.n56 output.n53 104.615
R23477 output.n104 output.n103 104.615
R23478 output.n103 output.n81 104.615
R23479 output.n96 output.n81 104.615
R23480 output.n96 output.n95 104.615
R23481 output.n95 output.n85 104.615
R23482 output.n88 output.n85 104.615
R23483 output.n136 output.n135 104.615
R23484 output.n135 output.n113 104.615
R23485 output.n128 output.n113 104.615
R23486 output.n128 output.n127 104.615
R23487 output.n127 output.n117 104.615
R23488 output.n120 output.n117 104.615
R23489 output.n1 output.t16 77.056
R23490 output.n14 output.t18 76.6694
R23491 output.n1 output.n0 72.7095
R23492 output.n3 output.n2 72.7095
R23493 output.n5 output.n4 72.7095
R23494 output.n7 output.n6 72.7095
R23495 output.n9 output.n8 72.7095
R23496 output.n11 output.n10 72.7095
R23497 output.n13 output.n12 72.7095
R23498 output.n25 output.t1 52.3082
R23499 output.n56 output.t0 52.3082
R23500 output.n88 output.t2 52.3082
R23501 output.n120 output.t19 52.3082
R23502 output.n26 output.n24 15.6674
R23503 output.n57 output.n55 15.6674
R23504 output.n89 output.n87 15.6674
R23505 output.n121 output.n119 15.6674
R23506 output.n27 output.n23 12.8005
R23507 output.n58 output.n54 12.8005
R23508 output.n90 output.n86 12.8005
R23509 output.n122 output.n118 12.8005
R23510 output.n31 output.n30 12.0247
R23511 output.n62 output.n61 12.0247
R23512 output.n94 output.n93 12.0247
R23513 output.n126 output.n125 12.0247
R23514 output.n34 output.n21 11.249
R23515 output.n65 output.n52 11.249
R23516 output.n97 output.n84 11.249
R23517 output.n129 output.n116 11.249
R23518 output.n35 output.n19 10.4732
R23519 output.n66 output.n50 10.4732
R23520 output.n98 output.n82 10.4732
R23521 output.n130 output.n114 10.4732
R23522 output.n39 output.n38 9.69747
R23523 output.n70 output.n69 9.69747
R23524 output.n102 output.n101 9.69747
R23525 output.n134 output.n133 9.69747
R23526 output.n45 output.n44 9.45567
R23527 output.n76 output.n75 9.45567
R23528 output.n108 output.n107 9.45567
R23529 output.n140 output.n139 9.45567
R23530 output.n44 output.n43 9.3005
R23531 output.n17 output.n16 9.3005
R23532 output.n38 output.n37 9.3005
R23533 output.n36 output.n35 9.3005
R23534 output.n21 output.n20 9.3005
R23535 output.n30 output.n29 9.3005
R23536 output.n28 output.n27 9.3005
R23537 output.n75 output.n74 9.3005
R23538 output.n48 output.n47 9.3005
R23539 output.n69 output.n68 9.3005
R23540 output.n67 output.n66 9.3005
R23541 output.n52 output.n51 9.3005
R23542 output.n61 output.n60 9.3005
R23543 output.n59 output.n58 9.3005
R23544 output.n107 output.n106 9.3005
R23545 output.n80 output.n79 9.3005
R23546 output.n101 output.n100 9.3005
R23547 output.n99 output.n98 9.3005
R23548 output.n84 output.n83 9.3005
R23549 output.n93 output.n92 9.3005
R23550 output.n91 output.n90 9.3005
R23551 output.n139 output.n138 9.3005
R23552 output.n112 output.n111 9.3005
R23553 output.n133 output.n132 9.3005
R23554 output.n131 output.n130 9.3005
R23555 output.n116 output.n115 9.3005
R23556 output.n125 output.n124 9.3005
R23557 output.n123 output.n122 9.3005
R23558 output.n42 output.n17 8.92171
R23559 output.n73 output.n48 8.92171
R23560 output.n105 output.n80 8.92171
R23561 output.n137 output.n112 8.92171
R23562 output output.n141 8.15037
R23563 output.n43 output.n15 8.14595
R23564 output.n74 output.n46 8.14595
R23565 output.n106 output.n78 8.14595
R23566 output.n138 output.n110 8.14595
R23567 output.n45 output.n15 5.81868
R23568 output.n76 output.n46 5.81868
R23569 output.n108 output.n78 5.81868
R23570 output.n140 output.n110 5.81868
R23571 output.n43 output.n42 5.04292
R23572 output.n74 output.n73 5.04292
R23573 output.n106 output.n105 5.04292
R23574 output.n138 output.n137 5.04292
R23575 output.n28 output.n24 4.38594
R23576 output.n59 output.n55 4.38594
R23577 output.n91 output.n87 4.38594
R23578 output.n123 output.n119 4.38594
R23579 output.n39 output.n17 4.26717
R23580 output.n70 output.n48 4.26717
R23581 output.n102 output.n80 4.26717
R23582 output.n134 output.n112 4.26717
R23583 output.n0 output.t12 3.9605
R23584 output.n0 output.t10 3.9605
R23585 output.n2 output.t4 3.9605
R23586 output.n2 output.t6 3.9605
R23587 output.n4 output.t7 3.9605
R23588 output.n4 output.t14 3.9605
R23589 output.n6 output.t17 3.9605
R23590 output.n6 output.t5 3.9605
R23591 output.n8 output.t8 3.9605
R23592 output.n8 output.t13 3.9605
R23593 output.n10 output.t15 3.9605
R23594 output.n10 output.t3 3.9605
R23595 output.n12 output.t11 3.9605
R23596 output.n12 output.t9 3.9605
R23597 output.n38 output.n19 3.49141
R23598 output.n69 output.n50 3.49141
R23599 output.n101 output.n82 3.49141
R23600 output.n133 output.n114 3.49141
R23601 output.n35 output.n34 2.71565
R23602 output.n66 output.n65 2.71565
R23603 output.n98 output.n97 2.71565
R23604 output.n130 output.n129 2.71565
R23605 output.n31 output.n21 1.93989
R23606 output.n62 output.n52 1.93989
R23607 output.n94 output.n84 1.93989
R23608 output.n126 output.n116 1.93989
R23609 output.n30 output.n23 1.16414
R23610 output.n61 output.n54 1.16414
R23611 output.n93 output.n86 1.16414
R23612 output.n125 output.n118 1.16414
R23613 output.n141 output.n109 0.962709
R23614 output.n109 output.n77 0.962709
R23615 output.n27 output.n26 0.388379
R23616 output.n58 output.n57 0.388379
R23617 output.n90 output.n89 0.388379
R23618 output.n122 output.n121 0.388379
R23619 output.n14 output.n13 0.387128
R23620 output.n13 output.n11 0.387128
R23621 output.n11 output.n9 0.387128
R23622 output.n9 output.n7 0.387128
R23623 output.n7 output.n5 0.387128
R23624 output.n5 output.n3 0.387128
R23625 output.n3 output.n1 0.387128
R23626 output.n44 output.n16 0.155672
R23627 output.n37 output.n16 0.155672
R23628 output.n37 output.n36 0.155672
R23629 output.n36 output.n20 0.155672
R23630 output.n29 output.n20 0.155672
R23631 output.n29 output.n28 0.155672
R23632 output.n75 output.n47 0.155672
R23633 output.n68 output.n47 0.155672
R23634 output.n68 output.n67 0.155672
R23635 output.n67 output.n51 0.155672
R23636 output.n60 output.n51 0.155672
R23637 output.n60 output.n59 0.155672
R23638 output.n107 output.n79 0.155672
R23639 output.n100 output.n79 0.155672
R23640 output.n100 output.n99 0.155672
R23641 output.n99 output.n83 0.155672
R23642 output.n92 output.n83 0.155672
R23643 output.n92 output.n91 0.155672
R23644 output.n139 output.n111 0.155672
R23645 output.n132 output.n111 0.155672
R23646 output.n132 output.n131 0.155672
R23647 output.n131 output.n115 0.155672
R23648 output.n124 output.n115 0.155672
R23649 output.n124 output.n123 0.155672
R23650 output output.n14 0.126227
R23651 minus.n33 minus.t20 321.495
R23652 minus.n7 minus.t6 321.495
R23653 minus.n50 minus.t18 297.12
R23654 minus.n48 minus.t15 297.12
R23655 minus.n28 minus.t16 297.12
R23656 minus.n42 minus.t11 297.12
R23657 minus.n30 minus.t12 297.12
R23658 minus.n36 minus.t7 297.12
R23659 minus.n32 minus.t19 297.12
R23660 minus.n6 minus.t5 297.12
R23661 minus.n10 minus.t9 297.12
R23662 minus.n12 minus.t8 297.12
R23663 minus.n16 minus.t10 297.12
R23664 minus.n18 minus.t14 297.12
R23665 minus.n22 minus.t13 297.12
R23666 minus.n24 minus.t17 297.12
R23667 minus.n56 minus.t4 243.255
R23668 minus.n55 minus.n53 224.169
R23669 minus.n55 minus.n54 223.454
R23670 minus.n35 minus.n34 161.3
R23671 minus.n36 minus.n31 161.3
R23672 minus.n38 minus.n37 161.3
R23673 minus.n39 minus.n30 161.3
R23674 minus.n41 minus.n40 161.3
R23675 minus.n42 minus.n29 161.3
R23676 minus.n44 minus.n43 161.3
R23677 minus.n45 minus.n28 161.3
R23678 minus.n47 minus.n46 161.3
R23679 minus.n48 minus.n27 161.3
R23680 minus.n49 minus.n26 161.3
R23681 minus.n51 minus.n50 161.3
R23682 minus.n25 minus.n24 161.3
R23683 minus.n23 minus.n0 161.3
R23684 minus.n22 minus.n21 161.3
R23685 minus.n20 minus.n1 161.3
R23686 minus.n19 minus.n18 161.3
R23687 minus.n17 minus.n2 161.3
R23688 minus.n16 minus.n15 161.3
R23689 minus.n14 minus.n3 161.3
R23690 minus.n13 minus.n12 161.3
R23691 minus.n11 minus.n4 161.3
R23692 minus.n10 minus.n9 161.3
R23693 minus.n8 minus.n5 161.3
R23694 minus.n8 minus.n7 44.9377
R23695 minus.n34 minus.n33 44.9377
R23696 minus.n50 minus.n49 37.246
R23697 minus.n24 minus.n23 37.246
R23698 minus.n48 minus.n47 32.8641
R23699 minus.n35 minus.n32 32.8641
R23700 minus.n6 minus.n5 32.8641
R23701 minus.n22 minus.n1 32.8641
R23702 minus.n52 minus.n51 30.2486
R23703 minus.n43 minus.n28 28.4823
R23704 minus.n37 minus.n36 28.4823
R23705 minus.n11 minus.n10 28.4823
R23706 minus.n18 minus.n17 28.4823
R23707 minus.n42 minus.n41 24.1005
R23708 minus.n41 minus.n30 24.1005
R23709 minus.n12 minus.n3 24.1005
R23710 minus.n16 minus.n3 24.1005
R23711 minus.n54 minus.t3 19.8005
R23712 minus.n54 minus.t2 19.8005
R23713 minus.n53 minus.t1 19.8005
R23714 minus.n53 minus.t0 19.8005
R23715 minus.n43 minus.n42 19.7187
R23716 minus.n37 minus.n30 19.7187
R23717 minus.n12 minus.n11 19.7187
R23718 minus.n17 minus.n16 19.7187
R23719 minus.n33 minus.n32 17.0522
R23720 minus.n7 minus.n6 17.0522
R23721 minus.n47 minus.n28 15.3369
R23722 minus.n36 minus.n35 15.3369
R23723 minus.n10 minus.n5 15.3369
R23724 minus.n18 minus.n1 15.3369
R23725 minus.n52 minus.n25 12.0706
R23726 minus minus.n57 11.7484
R23727 minus.n49 minus.n48 10.955
R23728 minus.n23 minus.n22 10.955
R23729 minus.n57 minus.n56 4.80222
R23730 minus.n57 minus.n52 0.972091
R23731 minus.n56 minus.n55 0.716017
R23732 minus.n51 minus.n26 0.189894
R23733 minus.n27 minus.n26 0.189894
R23734 minus.n46 minus.n27 0.189894
R23735 minus.n46 minus.n45 0.189894
R23736 minus.n45 minus.n44 0.189894
R23737 minus.n44 minus.n29 0.189894
R23738 minus.n40 minus.n29 0.189894
R23739 minus.n40 minus.n39 0.189894
R23740 minus.n39 minus.n38 0.189894
R23741 minus.n38 minus.n31 0.189894
R23742 minus.n34 minus.n31 0.189894
R23743 minus.n9 minus.n8 0.189894
R23744 minus.n9 minus.n4 0.189894
R23745 minus.n13 minus.n4 0.189894
R23746 minus.n14 minus.n13 0.189894
R23747 minus.n15 minus.n14 0.189894
R23748 minus.n15 minus.n2 0.189894
R23749 minus.n19 minus.n2 0.189894
R23750 minus.n20 minus.n19 0.189894
R23751 minus.n21 minus.n20 0.189894
R23752 minus.n21 minus.n0 0.189894
R23753 minus.n25 minus.n0 0.189894
R23754 diffpairibias.n0 diffpairibias.t18 436.822
R23755 diffpairibias.n21 diffpairibias.t19 435.479
R23756 diffpairibias.n20 diffpairibias.t16 435.479
R23757 diffpairibias.n19 diffpairibias.t17 435.479
R23758 diffpairibias.n18 diffpairibias.t21 435.479
R23759 diffpairibias.n0 diffpairibias.t22 435.479
R23760 diffpairibias.n1 diffpairibias.t20 435.479
R23761 diffpairibias.n2 diffpairibias.t23 435.479
R23762 diffpairibias.n10 diffpairibias.t0 377.536
R23763 diffpairibias.n10 diffpairibias.t8 376.193
R23764 diffpairibias.n11 diffpairibias.t10 376.193
R23765 diffpairibias.n12 diffpairibias.t6 376.193
R23766 diffpairibias.n13 diffpairibias.t2 376.193
R23767 diffpairibias.n14 diffpairibias.t12 376.193
R23768 diffpairibias.n15 diffpairibias.t4 376.193
R23769 diffpairibias.n16 diffpairibias.t14 376.193
R23770 diffpairibias.n3 diffpairibias.t1 113.368
R23771 diffpairibias.n3 diffpairibias.t9 112.698
R23772 diffpairibias.n4 diffpairibias.t11 112.698
R23773 diffpairibias.n5 diffpairibias.t7 112.698
R23774 diffpairibias.n6 diffpairibias.t3 112.698
R23775 diffpairibias.n7 diffpairibias.t13 112.698
R23776 diffpairibias.n8 diffpairibias.t5 112.698
R23777 diffpairibias.n9 diffpairibias.t15 112.698
R23778 diffpairibias.n17 diffpairibias.n16 4.77242
R23779 diffpairibias.n17 diffpairibias.n9 4.30807
R23780 diffpairibias.n18 diffpairibias.n17 4.13945
R23781 diffpairibias.n16 diffpairibias.n15 1.34352
R23782 diffpairibias.n15 diffpairibias.n14 1.34352
R23783 diffpairibias.n14 diffpairibias.n13 1.34352
R23784 diffpairibias.n13 diffpairibias.n12 1.34352
R23785 diffpairibias.n12 diffpairibias.n11 1.34352
R23786 diffpairibias.n11 diffpairibias.n10 1.34352
R23787 diffpairibias.n2 diffpairibias.n1 1.34352
R23788 diffpairibias.n1 diffpairibias.n0 1.34352
R23789 diffpairibias.n19 diffpairibias.n18 1.34352
R23790 diffpairibias.n20 diffpairibias.n19 1.34352
R23791 diffpairibias.n21 diffpairibias.n20 1.34352
R23792 diffpairibias.n22 diffpairibias.n21 0.862419
R23793 diffpairibias diffpairibias.n22 0.684875
R23794 diffpairibias.n9 diffpairibias.n8 0.672012
R23795 diffpairibias.n8 diffpairibias.n7 0.672012
R23796 diffpairibias.n7 diffpairibias.n6 0.672012
R23797 diffpairibias.n6 diffpairibias.n5 0.672012
R23798 diffpairibias.n5 diffpairibias.n4 0.672012
R23799 diffpairibias.n4 diffpairibias.n3 0.672012
R23800 diffpairibias.n22 diffpairibias.n2 0.190907
R23801 outputibias.n27 outputibias.n1 289.615
R23802 outputibias.n58 outputibias.n32 289.615
R23803 outputibias.n90 outputibias.n64 289.615
R23804 outputibias.n122 outputibias.n96 289.615
R23805 outputibias.n28 outputibias.n27 185
R23806 outputibias.n26 outputibias.n25 185
R23807 outputibias.n5 outputibias.n4 185
R23808 outputibias.n20 outputibias.n19 185
R23809 outputibias.n18 outputibias.n17 185
R23810 outputibias.n9 outputibias.n8 185
R23811 outputibias.n12 outputibias.n11 185
R23812 outputibias.n59 outputibias.n58 185
R23813 outputibias.n57 outputibias.n56 185
R23814 outputibias.n36 outputibias.n35 185
R23815 outputibias.n51 outputibias.n50 185
R23816 outputibias.n49 outputibias.n48 185
R23817 outputibias.n40 outputibias.n39 185
R23818 outputibias.n43 outputibias.n42 185
R23819 outputibias.n91 outputibias.n90 185
R23820 outputibias.n89 outputibias.n88 185
R23821 outputibias.n68 outputibias.n67 185
R23822 outputibias.n83 outputibias.n82 185
R23823 outputibias.n81 outputibias.n80 185
R23824 outputibias.n72 outputibias.n71 185
R23825 outputibias.n75 outputibias.n74 185
R23826 outputibias.n123 outputibias.n122 185
R23827 outputibias.n121 outputibias.n120 185
R23828 outputibias.n100 outputibias.n99 185
R23829 outputibias.n115 outputibias.n114 185
R23830 outputibias.n113 outputibias.n112 185
R23831 outputibias.n104 outputibias.n103 185
R23832 outputibias.n107 outputibias.n106 185
R23833 outputibias.n0 outputibias.t10 178.945
R23834 outputibias.n133 outputibias.t8 177.018
R23835 outputibias.n132 outputibias.t11 177.018
R23836 outputibias.n0 outputibias.t9 177.018
R23837 outputibias.t7 outputibias.n10 147.661
R23838 outputibias.t3 outputibias.n41 147.661
R23839 outputibias.t1 outputibias.n73 147.661
R23840 outputibias.t5 outputibias.n105 147.661
R23841 outputibias.n128 outputibias.t6 132.363
R23842 outputibias.n128 outputibias.t2 130.436
R23843 outputibias.n129 outputibias.t0 130.436
R23844 outputibias.n130 outputibias.t4 130.436
R23845 outputibias.n27 outputibias.n26 104.615
R23846 outputibias.n26 outputibias.n4 104.615
R23847 outputibias.n19 outputibias.n4 104.615
R23848 outputibias.n19 outputibias.n18 104.615
R23849 outputibias.n18 outputibias.n8 104.615
R23850 outputibias.n11 outputibias.n8 104.615
R23851 outputibias.n58 outputibias.n57 104.615
R23852 outputibias.n57 outputibias.n35 104.615
R23853 outputibias.n50 outputibias.n35 104.615
R23854 outputibias.n50 outputibias.n49 104.615
R23855 outputibias.n49 outputibias.n39 104.615
R23856 outputibias.n42 outputibias.n39 104.615
R23857 outputibias.n90 outputibias.n89 104.615
R23858 outputibias.n89 outputibias.n67 104.615
R23859 outputibias.n82 outputibias.n67 104.615
R23860 outputibias.n82 outputibias.n81 104.615
R23861 outputibias.n81 outputibias.n71 104.615
R23862 outputibias.n74 outputibias.n71 104.615
R23863 outputibias.n122 outputibias.n121 104.615
R23864 outputibias.n121 outputibias.n99 104.615
R23865 outputibias.n114 outputibias.n99 104.615
R23866 outputibias.n114 outputibias.n113 104.615
R23867 outputibias.n113 outputibias.n103 104.615
R23868 outputibias.n106 outputibias.n103 104.615
R23869 outputibias.n63 outputibias.n31 95.6354
R23870 outputibias.n63 outputibias.n62 94.6732
R23871 outputibias.n95 outputibias.n94 94.6732
R23872 outputibias.n127 outputibias.n126 94.6732
R23873 outputibias.n11 outputibias.t7 52.3082
R23874 outputibias.n42 outputibias.t3 52.3082
R23875 outputibias.n74 outputibias.t1 52.3082
R23876 outputibias.n106 outputibias.t5 52.3082
R23877 outputibias.n12 outputibias.n10 15.6674
R23878 outputibias.n43 outputibias.n41 15.6674
R23879 outputibias.n75 outputibias.n73 15.6674
R23880 outputibias.n107 outputibias.n105 15.6674
R23881 outputibias.n13 outputibias.n9 12.8005
R23882 outputibias.n44 outputibias.n40 12.8005
R23883 outputibias.n76 outputibias.n72 12.8005
R23884 outputibias.n108 outputibias.n104 12.8005
R23885 outputibias.n17 outputibias.n16 12.0247
R23886 outputibias.n48 outputibias.n47 12.0247
R23887 outputibias.n80 outputibias.n79 12.0247
R23888 outputibias.n112 outputibias.n111 12.0247
R23889 outputibias.n20 outputibias.n7 11.249
R23890 outputibias.n51 outputibias.n38 11.249
R23891 outputibias.n83 outputibias.n70 11.249
R23892 outputibias.n115 outputibias.n102 11.249
R23893 outputibias.n21 outputibias.n5 10.4732
R23894 outputibias.n52 outputibias.n36 10.4732
R23895 outputibias.n84 outputibias.n68 10.4732
R23896 outputibias.n116 outputibias.n100 10.4732
R23897 outputibias.n25 outputibias.n24 9.69747
R23898 outputibias.n56 outputibias.n55 9.69747
R23899 outputibias.n88 outputibias.n87 9.69747
R23900 outputibias.n120 outputibias.n119 9.69747
R23901 outputibias.n31 outputibias.n30 9.45567
R23902 outputibias.n62 outputibias.n61 9.45567
R23903 outputibias.n94 outputibias.n93 9.45567
R23904 outputibias.n126 outputibias.n125 9.45567
R23905 outputibias.n30 outputibias.n29 9.3005
R23906 outputibias.n3 outputibias.n2 9.3005
R23907 outputibias.n24 outputibias.n23 9.3005
R23908 outputibias.n22 outputibias.n21 9.3005
R23909 outputibias.n7 outputibias.n6 9.3005
R23910 outputibias.n16 outputibias.n15 9.3005
R23911 outputibias.n14 outputibias.n13 9.3005
R23912 outputibias.n61 outputibias.n60 9.3005
R23913 outputibias.n34 outputibias.n33 9.3005
R23914 outputibias.n55 outputibias.n54 9.3005
R23915 outputibias.n53 outputibias.n52 9.3005
R23916 outputibias.n38 outputibias.n37 9.3005
R23917 outputibias.n47 outputibias.n46 9.3005
R23918 outputibias.n45 outputibias.n44 9.3005
R23919 outputibias.n93 outputibias.n92 9.3005
R23920 outputibias.n66 outputibias.n65 9.3005
R23921 outputibias.n87 outputibias.n86 9.3005
R23922 outputibias.n85 outputibias.n84 9.3005
R23923 outputibias.n70 outputibias.n69 9.3005
R23924 outputibias.n79 outputibias.n78 9.3005
R23925 outputibias.n77 outputibias.n76 9.3005
R23926 outputibias.n125 outputibias.n124 9.3005
R23927 outputibias.n98 outputibias.n97 9.3005
R23928 outputibias.n119 outputibias.n118 9.3005
R23929 outputibias.n117 outputibias.n116 9.3005
R23930 outputibias.n102 outputibias.n101 9.3005
R23931 outputibias.n111 outputibias.n110 9.3005
R23932 outputibias.n109 outputibias.n108 9.3005
R23933 outputibias.n28 outputibias.n3 8.92171
R23934 outputibias.n59 outputibias.n34 8.92171
R23935 outputibias.n91 outputibias.n66 8.92171
R23936 outputibias.n123 outputibias.n98 8.92171
R23937 outputibias.n29 outputibias.n1 8.14595
R23938 outputibias.n60 outputibias.n32 8.14595
R23939 outputibias.n92 outputibias.n64 8.14595
R23940 outputibias.n124 outputibias.n96 8.14595
R23941 outputibias.n31 outputibias.n1 5.81868
R23942 outputibias.n62 outputibias.n32 5.81868
R23943 outputibias.n94 outputibias.n64 5.81868
R23944 outputibias.n126 outputibias.n96 5.81868
R23945 outputibias.n131 outputibias.n130 5.20947
R23946 outputibias.n29 outputibias.n28 5.04292
R23947 outputibias.n60 outputibias.n59 5.04292
R23948 outputibias.n92 outputibias.n91 5.04292
R23949 outputibias.n124 outputibias.n123 5.04292
R23950 outputibias.n131 outputibias.n127 4.42209
R23951 outputibias.n14 outputibias.n10 4.38594
R23952 outputibias.n45 outputibias.n41 4.38594
R23953 outputibias.n77 outputibias.n73 4.38594
R23954 outputibias.n109 outputibias.n105 4.38594
R23955 outputibias.n132 outputibias.n131 4.28454
R23956 outputibias.n25 outputibias.n3 4.26717
R23957 outputibias.n56 outputibias.n34 4.26717
R23958 outputibias.n88 outputibias.n66 4.26717
R23959 outputibias.n120 outputibias.n98 4.26717
R23960 outputibias.n24 outputibias.n5 3.49141
R23961 outputibias.n55 outputibias.n36 3.49141
R23962 outputibias.n87 outputibias.n68 3.49141
R23963 outputibias.n119 outputibias.n100 3.49141
R23964 outputibias.n21 outputibias.n20 2.71565
R23965 outputibias.n52 outputibias.n51 2.71565
R23966 outputibias.n84 outputibias.n83 2.71565
R23967 outputibias.n116 outputibias.n115 2.71565
R23968 outputibias.n17 outputibias.n7 1.93989
R23969 outputibias.n48 outputibias.n38 1.93989
R23970 outputibias.n80 outputibias.n70 1.93989
R23971 outputibias.n112 outputibias.n102 1.93989
R23972 outputibias.n130 outputibias.n129 1.9266
R23973 outputibias.n129 outputibias.n128 1.9266
R23974 outputibias.n133 outputibias.n132 1.92658
R23975 outputibias.n134 outputibias.n133 1.29913
R23976 outputibias.n16 outputibias.n9 1.16414
R23977 outputibias.n47 outputibias.n40 1.16414
R23978 outputibias.n79 outputibias.n72 1.16414
R23979 outputibias.n111 outputibias.n104 1.16414
R23980 outputibias.n127 outputibias.n95 0.962709
R23981 outputibias.n95 outputibias.n63 0.962709
R23982 outputibias.n13 outputibias.n12 0.388379
R23983 outputibias.n44 outputibias.n43 0.388379
R23984 outputibias.n76 outputibias.n75 0.388379
R23985 outputibias.n108 outputibias.n107 0.388379
R23986 outputibias.n134 outputibias.n0 0.337251
R23987 outputibias outputibias.n134 0.302375
R23988 outputibias.n30 outputibias.n2 0.155672
R23989 outputibias.n23 outputibias.n2 0.155672
R23990 outputibias.n23 outputibias.n22 0.155672
R23991 outputibias.n22 outputibias.n6 0.155672
R23992 outputibias.n15 outputibias.n6 0.155672
R23993 outputibias.n15 outputibias.n14 0.155672
R23994 outputibias.n61 outputibias.n33 0.155672
R23995 outputibias.n54 outputibias.n33 0.155672
R23996 outputibias.n54 outputibias.n53 0.155672
R23997 outputibias.n53 outputibias.n37 0.155672
R23998 outputibias.n46 outputibias.n37 0.155672
R23999 outputibias.n46 outputibias.n45 0.155672
R24000 outputibias.n93 outputibias.n65 0.155672
R24001 outputibias.n86 outputibias.n65 0.155672
R24002 outputibias.n86 outputibias.n85 0.155672
R24003 outputibias.n85 outputibias.n69 0.155672
R24004 outputibias.n78 outputibias.n69 0.155672
R24005 outputibias.n78 outputibias.n77 0.155672
R24006 outputibias.n125 outputibias.n97 0.155672
R24007 outputibias.n118 outputibias.n97 0.155672
R24008 outputibias.n118 outputibias.n117 0.155672
R24009 outputibias.n117 outputibias.n101 0.155672
R24010 outputibias.n110 outputibias.n101 0.155672
R24011 outputibias.n110 outputibias.n109 0.155672
C0 CSoutput outputibias 0.032386f
C1 vdd CSoutput 0.14236p
C2 minus diffpairibias 3.1e-19
C3 commonsourceibias output 0.006829f
C4 vdd plus 0.098689f
C5 CSoutput minus 2.93147f
C6 plus diffpairibias 3.12e-19
C7 commonsourceibias outputibias 0.003902f
C8 CSoutput plus 0.847799f
C9 vdd commonsourceibias 0.004262f
C10 commonsourceibias diffpairibias 0.06482f
C11 minus plus 8.948191f
C12 CSoutput commonsourceibias 42.168602f
C13 minus commonsourceibias 0.318966f
C14 plus commonsourceibias 0.273048f
C15 output outputibias 2.34152f
C16 vdd output 7.23429f
C17 CSoutput output 6.13881f
C18 diffpairibias gnd 48.980038f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.144975p
C22 plus gnd 31.0858f
C23 minus gnd 26.46894f
C24 CSoutput gnd 0.107423p
C25 vdd gnd 0.542244p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t10 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t3 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t1 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t0 gnd 0.108319f
C162 outputibias.t2 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t8 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 minus.n0 gnd 0.030586f
C221 minus.n1 gnd 0.006941f
C222 minus.n2 gnd 0.030586f
C223 minus.n3 gnd 0.006941f
C224 minus.n4 gnd 0.030586f
C225 minus.n5 gnd 0.006941f
C226 minus.t6 gnd 0.447195f
C227 minus.t5 gnd 0.432615f
C228 minus.n6 gnd 0.196371f
C229 minus.n7 gnd 0.180147f
C230 minus.n8 gnd 0.129434f
C231 minus.n9 gnd 0.030586f
C232 minus.t9 gnd 0.432615f
C233 minus.n10 gnd 0.192181f
C234 minus.n11 gnd 0.006941f
C235 minus.t8 gnd 0.432615f
C236 minus.n12 gnd 0.192181f
C237 minus.n13 gnd 0.030586f
C238 minus.n14 gnd 0.030586f
C239 minus.n15 gnd 0.030586f
C240 minus.t10 gnd 0.432615f
C241 minus.n16 gnd 0.192181f
C242 minus.n17 gnd 0.006941f
C243 minus.t14 gnd 0.432615f
C244 minus.n18 gnd 0.192181f
C245 minus.n19 gnd 0.030586f
C246 minus.n20 gnd 0.030586f
C247 minus.n21 gnd 0.030586f
C248 minus.t13 gnd 0.432615f
C249 minus.n22 gnd 0.192181f
C250 minus.n23 gnd 0.006941f
C251 minus.t17 gnd 0.432615f
C252 minus.n24 gnd 0.191333f
C253 minus.n25 gnd 0.352582f
C254 minus.n26 gnd 0.030586f
C255 minus.t18 gnd 0.432615f
C256 minus.t15 gnd 0.432615f
C257 minus.n27 gnd 0.030586f
C258 minus.t16 gnd 0.432615f
C259 minus.n28 gnd 0.192181f
C260 minus.n29 gnd 0.030586f
C261 minus.t11 gnd 0.432615f
C262 minus.t12 gnd 0.432615f
C263 minus.n30 gnd 0.192181f
C264 minus.n31 gnd 0.030586f
C265 minus.t7 gnd 0.432615f
C266 minus.t19 gnd 0.432615f
C267 minus.n32 gnd 0.196371f
C268 minus.t20 gnd 0.447195f
C269 minus.n33 gnd 0.180147f
C270 minus.n34 gnd 0.129434f
C271 minus.n35 gnd 0.006941f
C272 minus.n36 gnd 0.192181f
C273 minus.n37 gnd 0.006941f
C274 minus.n38 gnd 0.030586f
C275 minus.n39 gnd 0.030586f
C276 minus.n40 gnd 0.030586f
C277 minus.n41 gnd 0.006941f
C278 minus.n42 gnd 0.192181f
C279 minus.n43 gnd 0.006941f
C280 minus.n44 gnd 0.030586f
C281 minus.n45 gnd 0.030586f
C282 minus.n46 gnd 0.030586f
C283 minus.n47 gnd 0.006941f
C284 minus.n48 gnd 0.192181f
C285 minus.n49 gnd 0.006941f
C286 minus.n50 gnd 0.191333f
C287 minus.n51 gnd 0.887772f
C288 minus.n52 gnd 1.34998f
C289 minus.t1 gnd 0.009429f
C290 minus.t0 gnd 0.009429f
C291 minus.n53 gnd 0.031004f
C292 minus.t3 gnd 0.009429f
C293 minus.t2 gnd 0.009429f
C294 minus.n54 gnd 0.030579f
C295 minus.n55 gnd 0.260982f
C296 minus.t4 gnd 0.05248f
C297 minus.n56 gnd 0.142415f
C298 minus.n57 gnd 2.06205f
C299 output.t16 gnd 0.464308f
C300 output.t12 gnd 0.044422f
C301 output.t10 gnd 0.044422f
C302 output.n0 gnd 0.364624f
C303 output.n1 gnd 0.614102f
C304 output.t4 gnd 0.044422f
C305 output.t6 gnd 0.044422f
C306 output.n2 gnd 0.364624f
C307 output.n3 gnd 0.350265f
C308 output.t7 gnd 0.044422f
C309 output.t14 gnd 0.044422f
C310 output.n4 gnd 0.364624f
C311 output.n5 gnd 0.350265f
C312 output.t17 gnd 0.044422f
C313 output.t5 gnd 0.044422f
C314 output.n6 gnd 0.364624f
C315 output.n7 gnd 0.350265f
C316 output.t8 gnd 0.044422f
C317 output.t13 gnd 0.044422f
C318 output.n8 gnd 0.364624f
C319 output.n9 gnd 0.350265f
C320 output.t15 gnd 0.044422f
C321 output.t3 gnd 0.044422f
C322 output.n10 gnd 0.364624f
C323 output.n11 gnd 0.350265f
C324 output.t11 gnd 0.044422f
C325 output.t9 gnd 0.044422f
C326 output.n12 gnd 0.364624f
C327 output.n13 gnd 0.350265f
C328 output.t18 gnd 0.462979f
C329 output.n14 gnd 0.28994f
C330 output.n15 gnd 0.015803f
C331 output.n16 gnd 0.011243f
C332 output.n17 gnd 0.006041f
C333 output.n18 gnd 0.01428f
C334 output.n19 gnd 0.006397f
C335 output.n20 gnd 0.011243f
C336 output.n21 gnd 0.006041f
C337 output.n22 gnd 0.01428f
C338 output.n23 gnd 0.006397f
C339 output.n24 gnd 0.048111f
C340 output.t1 gnd 0.023274f
C341 output.n25 gnd 0.01071f
C342 output.n26 gnd 0.008435f
C343 output.n27 gnd 0.006041f
C344 output.n28 gnd 0.267512f
C345 output.n29 gnd 0.011243f
C346 output.n30 gnd 0.006041f
C347 output.n31 gnd 0.006397f
C348 output.n32 gnd 0.01428f
C349 output.n33 gnd 0.01428f
C350 output.n34 gnd 0.006397f
C351 output.n35 gnd 0.006041f
C352 output.n36 gnd 0.011243f
C353 output.n37 gnd 0.011243f
C354 output.n38 gnd 0.006041f
C355 output.n39 gnd 0.006397f
C356 output.n40 gnd 0.01428f
C357 output.n41 gnd 0.030913f
C358 output.n42 gnd 0.006397f
C359 output.n43 gnd 0.006041f
C360 output.n44 gnd 0.025987f
C361 output.n45 gnd 0.097665f
C362 output.n46 gnd 0.015803f
C363 output.n47 gnd 0.011243f
C364 output.n48 gnd 0.006041f
C365 output.n49 gnd 0.01428f
C366 output.n50 gnd 0.006397f
C367 output.n51 gnd 0.011243f
C368 output.n52 gnd 0.006041f
C369 output.n53 gnd 0.01428f
C370 output.n54 gnd 0.006397f
C371 output.n55 gnd 0.048111f
C372 output.t0 gnd 0.023274f
C373 output.n56 gnd 0.01071f
C374 output.n57 gnd 0.008435f
C375 output.n58 gnd 0.006041f
C376 output.n59 gnd 0.267512f
C377 output.n60 gnd 0.011243f
C378 output.n61 gnd 0.006041f
C379 output.n62 gnd 0.006397f
C380 output.n63 gnd 0.01428f
C381 output.n64 gnd 0.01428f
C382 output.n65 gnd 0.006397f
C383 output.n66 gnd 0.006041f
C384 output.n67 gnd 0.011243f
C385 output.n68 gnd 0.011243f
C386 output.n69 gnd 0.006041f
C387 output.n70 gnd 0.006397f
C388 output.n71 gnd 0.01428f
C389 output.n72 gnd 0.030913f
C390 output.n73 gnd 0.006397f
C391 output.n74 gnd 0.006041f
C392 output.n75 gnd 0.025987f
C393 output.n76 gnd 0.09306f
C394 output.n77 gnd 1.65264f
C395 output.n78 gnd 0.015803f
C396 output.n79 gnd 0.011243f
C397 output.n80 gnd 0.006041f
C398 output.n81 gnd 0.01428f
C399 output.n82 gnd 0.006397f
C400 output.n83 gnd 0.011243f
C401 output.n84 gnd 0.006041f
C402 output.n85 gnd 0.01428f
C403 output.n86 gnd 0.006397f
C404 output.n87 gnd 0.048111f
C405 output.t2 gnd 0.023274f
C406 output.n88 gnd 0.01071f
C407 output.n89 gnd 0.008435f
C408 output.n90 gnd 0.006041f
C409 output.n91 gnd 0.267512f
C410 output.n92 gnd 0.011243f
C411 output.n93 gnd 0.006041f
C412 output.n94 gnd 0.006397f
C413 output.n95 gnd 0.01428f
C414 output.n96 gnd 0.01428f
C415 output.n97 gnd 0.006397f
C416 output.n98 gnd 0.006041f
C417 output.n99 gnd 0.011243f
C418 output.n100 gnd 0.011243f
C419 output.n101 gnd 0.006041f
C420 output.n102 gnd 0.006397f
C421 output.n103 gnd 0.01428f
C422 output.n104 gnd 0.030913f
C423 output.n105 gnd 0.006397f
C424 output.n106 gnd 0.006041f
C425 output.n107 gnd 0.025987f
C426 output.n108 gnd 0.09306f
C427 output.n109 gnd 0.713089f
C428 output.n110 gnd 0.015803f
C429 output.n111 gnd 0.011243f
C430 output.n112 gnd 0.006041f
C431 output.n113 gnd 0.01428f
C432 output.n114 gnd 0.006397f
C433 output.n115 gnd 0.011243f
C434 output.n116 gnd 0.006041f
C435 output.n117 gnd 0.01428f
C436 output.n118 gnd 0.006397f
C437 output.n119 gnd 0.048111f
C438 output.t19 gnd 0.023274f
C439 output.n120 gnd 0.01071f
C440 output.n121 gnd 0.008435f
C441 output.n122 gnd 0.006041f
C442 output.n123 gnd 0.267512f
C443 output.n124 gnd 0.011243f
C444 output.n125 gnd 0.006041f
C445 output.n126 gnd 0.006397f
C446 output.n127 gnd 0.01428f
C447 output.n128 gnd 0.01428f
C448 output.n129 gnd 0.006397f
C449 output.n130 gnd 0.006041f
C450 output.n131 gnd 0.011243f
C451 output.n132 gnd 0.011243f
C452 output.n133 gnd 0.006041f
C453 output.n134 gnd 0.006397f
C454 output.n135 gnd 0.01428f
C455 output.n136 gnd 0.030913f
C456 output.n137 gnd 0.006397f
C457 output.n138 gnd 0.006041f
C458 output.n139 gnd 0.025987f
C459 output.n140 gnd 0.09306f
C460 output.n141 gnd 1.67353f
C461 a_n2982_8322.t7 gnd 0.100161f
C462 a_n2982_8322.t34 gnd 20.7793f
C463 a_n2982_8322.t33 gnd 20.633598f
C464 a_n2982_8322.t37 gnd 20.633598f
C465 a_n2982_8322.t36 gnd 20.7793f
C466 a_n2982_8322.t35 gnd 20.633598f
C467 a_n2982_8322.t32 gnd 28.9697f
C468 a_n2982_8322.t6 gnd 0.937857f
C469 a_n2982_8322.t19 gnd 0.100161f
C470 a_n2982_8322.t15 gnd 0.100161f
C471 a_n2982_8322.n0 gnd 0.705534f
C472 a_n2982_8322.n1 gnd 0.78833f
C473 a_n2982_8322.t22 gnd 0.100161f
C474 a_n2982_8322.t12 gnd 0.100161f
C475 a_n2982_8322.n2 gnd 0.705534f
C476 a_n2982_8322.n3 gnd 0.40054f
C477 a_n2982_8322.t3 gnd 0.100161f
C478 a_n2982_8322.t2 gnd 0.100161f
C479 a_n2982_8322.n4 gnd 0.705534f
C480 a_n2982_8322.n5 gnd 0.40054f
C481 a_n2982_8322.t16 gnd 0.100161f
C482 a_n2982_8322.t9 gnd 0.100161f
C483 a_n2982_8322.n6 gnd 0.705534f
C484 a_n2982_8322.n7 gnd 0.40054f
C485 a_n2982_8322.t13 gnd 0.100161f
C486 a_n2982_8322.t11 gnd 0.100161f
C487 a_n2982_8322.n8 gnd 0.705534f
C488 a_n2982_8322.n9 gnd 0.40054f
C489 a_n2982_8322.t0 gnd 0.935989f
C490 a_n2982_8322.n10 gnd 1.87142f
C491 a_n2982_8322.t27 gnd 0.937857f
C492 a_n2982_8322.t31 gnd 0.100161f
C493 a_n2982_8322.t30 gnd 0.100161f
C494 a_n2982_8322.n11 gnd 0.705534f
C495 a_n2982_8322.n12 gnd 0.78833f
C496 a_n2982_8322.t25 gnd 0.935989f
C497 a_n2982_8322.n13 gnd 0.396699f
C498 a_n2982_8322.t28 gnd 0.935989f
C499 a_n2982_8322.n14 gnd 0.396699f
C500 a_n2982_8322.t26 gnd 0.100161f
C501 a_n2982_8322.t24 gnd 0.100161f
C502 a_n2982_8322.n15 gnd 0.705534f
C503 a_n2982_8322.n16 gnd 0.40054f
C504 a_n2982_8322.t29 gnd 0.935989f
C505 a_n2982_8322.n17 gnd 1.47143f
C506 a_n2982_8322.n18 gnd 2.35138f
C507 a_n2982_8322.n19 gnd 3.33814f
C508 a_n2982_8322.t1 gnd 0.935989f
C509 a_n2982_8322.n20 gnd 1.11148f
C510 a_n2982_8322.t18 gnd 0.100161f
C511 a_n2982_8322.t17 gnd 0.100161f
C512 a_n2982_8322.n21 gnd 0.705534f
C513 a_n2982_8322.n22 gnd 0.40054f
C514 a_n2982_8322.t5 gnd 0.100161f
C515 a_n2982_8322.t4 gnd 0.100161f
C516 a_n2982_8322.n23 gnd 0.705534f
C517 a_n2982_8322.n24 gnd 0.40054f
C518 a_n2982_8322.t20 gnd 0.100161f
C519 a_n2982_8322.t8 gnd 0.100161f
C520 a_n2982_8322.n25 gnd 0.705534f
C521 a_n2982_8322.n26 gnd 0.40054f
C522 a_n2982_8322.t21 gnd 0.937854f
C523 a_n2982_8322.t14 gnd 0.100161f
C524 a_n2982_8322.t10 gnd 0.100161f
C525 a_n2982_8322.n27 gnd 0.705534f
C526 a_n2982_8322.n28 gnd 0.788332f
C527 a_n2982_8322.n29 gnd 0.400539f
C528 a_n2982_8322.n30 gnd 0.705536f
C529 a_n2982_8322.t23 gnd 0.100161f
C530 a_n2804_13878.t29 gnd 0.194556f
C531 a_n2804_13878.t25 gnd 0.194556f
C532 a_n2804_13878.t31 gnd 0.194556f
C533 a_n2804_13878.n0 gnd 1.53449f
C534 a_n2804_13878.t8 gnd 0.194556f
C535 a_n2804_13878.t20 gnd 0.194556f
C536 a_n2804_13878.n1 gnd 1.53196f
C537 a_n2804_13878.n2 gnd 1.37704f
C538 a_n2804_13878.t12 gnd 0.194556f
C539 a_n2804_13878.t22 gnd 0.194556f
C540 a_n2804_13878.n3 gnd 1.53358f
C541 a_n2804_13878.t27 gnd 0.194556f
C542 a_n2804_13878.t17 gnd 0.194556f
C543 a_n2804_13878.n4 gnd 1.53196f
C544 a_n2804_13878.n5 gnd 2.14061f
C545 a_n2804_13878.t23 gnd 0.194556f
C546 a_n2804_13878.t16 gnd 0.194556f
C547 a_n2804_13878.n6 gnd 1.53196f
C548 a_n2804_13878.n7 gnd 1.04414f
C549 a_n2804_13878.t10 gnd 0.194556f
C550 a_n2804_13878.t13 gnd 0.194556f
C551 a_n2804_13878.n8 gnd 1.53196f
C552 a_n2804_13878.n9 gnd 1.04414f
C553 a_n2804_13878.t26 gnd 0.194556f
C554 a_n2804_13878.t11 gnd 0.194556f
C555 a_n2804_13878.n10 gnd 1.53196f
C556 a_n2804_13878.n11 gnd 1.04414f
C557 a_n2804_13878.t21 gnd 0.194556f
C558 a_n2804_13878.t9 gnd 0.194556f
C559 a_n2804_13878.n12 gnd 1.53196f
C560 a_n2804_13878.n13 gnd 4.90178f
C561 a_n2804_13878.t1 gnd 1.82172f
C562 a_n2804_13878.t4 gnd 0.194556f
C563 a_n2804_13878.t5 gnd 0.194556f
C564 a_n2804_13878.n14 gnd 1.37045f
C565 a_n2804_13878.n15 gnd 1.53128f
C566 a_n2804_13878.t0 gnd 1.81809f
C567 a_n2804_13878.n16 gnd 0.770559f
C568 a_n2804_13878.t3 gnd 1.81809f
C569 a_n2804_13878.n17 gnd 0.770559f
C570 a_n2804_13878.t6 gnd 0.194556f
C571 a_n2804_13878.t7 gnd 0.194556f
C572 a_n2804_13878.n18 gnd 1.37045f
C573 a_n2804_13878.n19 gnd 0.778022f
C574 a_n2804_13878.t2 gnd 1.81809f
C575 a_n2804_13878.n20 gnd 2.85814f
C576 a_n2804_13878.n21 gnd 3.74876f
C577 a_n2804_13878.t15 gnd 0.194556f
C578 a_n2804_13878.t24 gnd 0.194556f
C579 a_n2804_13878.n22 gnd 1.53195f
C580 a_n2804_13878.n23 gnd 2.50239f
C581 a_n2804_13878.t28 gnd 0.194556f
C582 a_n2804_13878.t14 gnd 0.194556f
C583 a_n2804_13878.n24 gnd 1.53196f
C584 a_n2804_13878.n25 gnd 0.678771f
C585 a_n2804_13878.t18 gnd 0.194556f
C586 a_n2804_13878.t19 gnd 0.194556f
C587 a_n2804_13878.n26 gnd 1.53196f
C588 a_n2804_13878.n27 gnd 0.678771f
C589 a_n2804_13878.n28 gnd 0.678768f
C590 a_n2804_13878.n29 gnd 1.53196f
C591 a_n2804_13878.t30 gnd 0.194556f
C592 vdd.t280 gnd 0.037058f
C593 vdd.t261 gnd 0.037058f
C594 vdd.n0 gnd 0.29228f
C595 vdd.t239 gnd 0.037058f
C596 vdd.t276 gnd 0.037058f
C597 vdd.n1 gnd 0.291797f
C598 vdd.n2 gnd 0.269092f
C599 vdd.t257 gnd 0.037058f
C600 vdd.t282 gnd 0.037058f
C601 vdd.n3 gnd 0.291797f
C602 vdd.n4 gnd 0.13609f
C603 vdd.t287 gnd 0.037058f
C604 vdd.t265 gnd 0.037058f
C605 vdd.n5 gnd 0.291797f
C606 vdd.n6 gnd 0.127695f
C607 vdd.t291 gnd 0.037058f
C608 vdd.t255 gnd 0.037058f
C609 vdd.n7 gnd 0.29228f
C610 vdd.t263 gnd 0.037058f
C611 vdd.t285 gnd 0.037058f
C612 vdd.n8 gnd 0.291797f
C613 vdd.n9 gnd 0.269093f
C614 vdd.t272 gnd 0.037058f
C615 vdd.t243 gnd 0.037058f
C616 vdd.n10 gnd 0.291797f
C617 vdd.n11 gnd 0.13609f
C618 vdd.t252 gnd 0.037058f
C619 vdd.t270 gnd 0.037058f
C620 vdd.n12 gnd 0.291797f
C621 vdd.n13 gnd 0.127695f
C622 vdd.n14 gnd 0.090278f
C623 vdd.t300 gnd 0.020588f
C624 vdd.t297 gnd 0.020588f
C625 vdd.n15 gnd 0.1895f
C626 vdd.t301 gnd 0.020588f
C627 vdd.t294 gnd 0.020588f
C628 vdd.n16 gnd 0.188945f
C629 vdd.n17 gnd 0.328824f
C630 vdd.t299 gnd 0.020588f
C631 vdd.t305 gnd 0.020588f
C632 vdd.n18 gnd 0.188945f
C633 vdd.n19 gnd 0.136039f
C634 vdd.t304 gnd 0.020588f
C635 vdd.t295 gnd 0.020588f
C636 vdd.n20 gnd 0.1895f
C637 vdd.t303 gnd 0.020588f
C638 vdd.t306 gnd 0.020588f
C639 vdd.n21 gnd 0.188945f
C640 vdd.n22 gnd 0.328824f
C641 vdd.t296 gnd 0.020588f
C642 vdd.t302 gnd 0.020588f
C643 vdd.n23 gnd 0.188945f
C644 vdd.n24 gnd 0.136039f
C645 vdd.t293 gnd 0.020588f
C646 vdd.t298 gnd 0.020588f
C647 vdd.n25 gnd 0.188945f
C648 vdd.t307 gnd 0.020588f
C649 vdd.t292 gnd 0.020588f
C650 vdd.n26 gnd 0.188945f
C651 vdd.n27 gnd 20.7697f
C652 vdd.n28 gnd 8.3397f
C653 vdd.n29 gnd 0.005615f
C654 vdd.n30 gnd 0.005211f
C655 vdd.n31 gnd 0.002882f
C656 vdd.n32 gnd 0.006618f
C657 vdd.n33 gnd 0.0028f
C658 vdd.n34 gnd 0.002965f
C659 vdd.n35 gnd 0.005211f
C660 vdd.n36 gnd 0.0028f
C661 vdd.n37 gnd 0.006618f
C662 vdd.n38 gnd 0.002965f
C663 vdd.n39 gnd 0.005211f
C664 vdd.n40 gnd 0.0028f
C665 vdd.n41 gnd 0.004963f
C666 vdd.n42 gnd 0.004978f
C667 vdd.t82 gnd 0.014218f
C668 vdd.n43 gnd 0.031635f
C669 vdd.n44 gnd 0.164637f
C670 vdd.n45 gnd 0.0028f
C671 vdd.n46 gnd 0.002965f
C672 vdd.n47 gnd 0.006618f
C673 vdd.n48 gnd 0.006618f
C674 vdd.n49 gnd 0.002965f
C675 vdd.n50 gnd 0.0028f
C676 vdd.n51 gnd 0.005211f
C677 vdd.n52 gnd 0.005211f
C678 vdd.n53 gnd 0.0028f
C679 vdd.n54 gnd 0.002965f
C680 vdd.n55 gnd 0.006618f
C681 vdd.n56 gnd 0.006618f
C682 vdd.n57 gnd 0.002965f
C683 vdd.n58 gnd 0.0028f
C684 vdd.n59 gnd 0.005211f
C685 vdd.n60 gnd 0.005211f
C686 vdd.n61 gnd 0.0028f
C687 vdd.n62 gnd 0.002965f
C688 vdd.n63 gnd 0.006618f
C689 vdd.n64 gnd 0.006618f
C690 vdd.n65 gnd 0.015646f
C691 vdd.n66 gnd 0.002882f
C692 vdd.n67 gnd 0.0028f
C693 vdd.n68 gnd 0.013467f
C694 vdd.n69 gnd 0.009402f
C695 vdd.t51 gnd 0.03294f
C696 vdd.t134 gnd 0.03294f
C697 vdd.n70 gnd 0.226387f
C698 vdd.n71 gnd 0.178019f
C699 vdd.t26 gnd 0.03294f
C700 vdd.t113 gnd 0.03294f
C701 vdd.n72 gnd 0.226387f
C702 vdd.n73 gnd 0.14366f
C703 vdd.t34 gnd 0.03294f
C704 vdd.t127 gnd 0.03294f
C705 vdd.n74 gnd 0.226387f
C706 vdd.n75 gnd 0.14366f
C707 vdd.t65 gnd 0.03294f
C708 vdd.t144 gnd 0.03294f
C709 vdd.n76 gnd 0.226387f
C710 vdd.n77 gnd 0.14366f
C711 vdd.t89 gnd 0.03294f
C712 vdd.t119 gnd 0.03294f
C713 vdd.n78 gnd 0.226387f
C714 vdd.n79 gnd 0.14366f
C715 vdd.t54 gnd 0.03294f
C716 vdd.t136 gnd 0.03294f
C717 vdd.n80 gnd 0.226387f
C718 vdd.n81 gnd 0.14366f
C719 vdd.t75 gnd 0.03294f
C720 vdd.t155 gnd 0.03294f
C721 vdd.n82 gnd 0.226387f
C722 vdd.n83 gnd 0.14366f
C723 vdd.t100 gnd 0.03294f
C724 vdd.t3 gnd 0.03294f
C725 vdd.n84 gnd 0.226387f
C726 vdd.n85 gnd 0.14366f
C727 vdd.t67 gnd 0.03294f
C728 vdd.t145 gnd 0.03294f
C729 vdd.n86 gnd 0.226387f
C730 vdd.n87 gnd 0.14366f
C731 vdd.n88 gnd 0.005615f
C732 vdd.n89 gnd 0.005211f
C733 vdd.n90 gnd 0.002882f
C734 vdd.n91 gnd 0.006618f
C735 vdd.n92 gnd 0.0028f
C736 vdd.n93 gnd 0.002965f
C737 vdd.n94 gnd 0.005211f
C738 vdd.n95 gnd 0.0028f
C739 vdd.n96 gnd 0.006618f
C740 vdd.n97 gnd 0.002965f
C741 vdd.n98 gnd 0.005211f
C742 vdd.n99 gnd 0.0028f
C743 vdd.n100 gnd 0.004963f
C744 vdd.n101 gnd 0.004978f
C745 vdd.t122 gnd 0.014218f
C746 vdd.n102 gnd 0.031635f
C747 vdd.n103 gnd 0.164637f
C748 vdd.n104 gnd 0.0028f
C749 vdd.n105 gnd 0.002965f
C750 vdd.n106 gnd 0.006618f
C751 vdd.n107 gnd 0.006618f
C752 vdd.n108 gnd 0.002965f
C753 vdd.n109 gnd 0.0028f
C754 vdd.n110 gnd 0.005211f
C755 vdd.n111 gnd 0.005211f
C756 vdd.n112 gnd 0.0028f
C757 vdd.n113 gnd 0.002965f
C758 vdd.n114 gnd 0.006618f
C759 vdd.n115 gnd 0.006618f
C760 vdd.n116 gnd 0.002965f
C761 vdd.n117 gnd 0.0028f
C762 vdd.n118 gnd 0.005211f
C763 vdd.n119 gnd 0.005211f
C764 vdd.n120 gnd 0.0028f
C765 vdd.n121 gnd 0.002965f
C766 vdd.n122 gnd 0.006618f
C767 vdd.n123 gnd 0.006618f
C768 vdd.n124 gnd 0.015646f
C769 vdd.n125 gnd 0.002882f
C770 vdd.n126 gnd 0.0028f
C771 vdd.n127 gnd 0.013467f
C772 vdd.n128 gnd 0.009107f
C773 vdd.n129 gnd 0.106884f
C774 vdd.n130 gnd 0.005615f
C775 vdd.n131 gnd 0.005211f
C776 vdd.n132 gnd 0.002882f
C777 vdd.n133 gnd 0.006618f
C778 vdd.n134 gnd 0.0028f
C779 vdd.n135 gnd 0.002965f
C780 vdd.n136 gnd 0.005211f
C781 vdd.n137 gnd 0.0028f
C782 vdd.n138 gnd 0.006618f
C783 vdd.n139 gnd 0.002965f
C784 vdd.n140 gnd 0.005211f
C785 vdd.n141 gnd 0.0028f
C786 vdd.n142 gnd 0.004963f
C787 vdd.n143 gnd 0.004978f
C788 vdd.t141 gnd 0.014218f
C789 vdd.n144 gnd 0.031635f
C790 vdd.n145 gnd 0.164637f
C791 vdd.n146 gnd 0.0028f
C792 vdd.n147 gnd 0.002965f
C793 vdd.n148 gnd 0.006618f
C794 vdd.n149 gnd 0.006618f
C795 vdd.n150 gnd 0.002965f
C796 vdd.n151 gnd 0.0028f
C797 vdd.n152 gnd 0.005211f
C798 vdd.n153 gnd 0.005211f
C799 vdd.n154 gnd 0.0028f
C800 vdd.n155 gnd 0.002965f
C801 vdd.n156 gnd 0.006618f
C802 vdd.n157 gnd 0.006618f
C803 vdd.n158 gnd 0.002965f
C804 vdd.n159 gnd 0.0028f
C805 vdd.n160 gnd 0.005211f
C806 vdd.n161 gnd 0.005211f
C807 vdd.n162 gnd 0.0028f
C808 vdd.n163 gnd 0.002965f
C809 vdd.n164 gnd 0.006618f
C810 vdd.n165 gnd 0.006618f
C811 vdd.n166 gnd 0.015646f
C812 vdd.n167 gnd 0.002882f
C813 vdd.n168 gnd 0.0028f
C814 vdd.n169 gnd 0.013467f
C815 vdd.n170 gnd 0.009402f
C816 vdd.t142 gnd 0.03294f
C817 vdd.t23 gnd 0.03294f
C818 vdd.n171 gnd 0.226387f
C819 vdd.n172 gnd 0.178019f
C820 vdd.t121 gnd 0.03294f
C821 vdd.t133 gnd 0.03294f
C822 vdd.n173 gnd 0.226387f
C823 vdd.n174 gnd 0.14366f
C824 vdd.t17 gnd 0.03294f
C825 vdd.t80 gnd 0.03294f
C826 vdd.n175 gnd 0.226387f
C827 vdd.n176 gnd 0.14366f
C828 vdd.t118 gnd 0.03294f
C829 vdd.t150 gnd 0.03294f
C830 vdd.n177 gnd 0.226387f
C831 vdd.n178 gnd 0.14366f
C832 vdd.t57 gnd 0.03294f
C833 vdd.t117 gnd 0.03294f
C834 vdd.n179 gnd 0.226387f
C835 vdd.n180 gnd 0.14366f
C836 vdd.t158 gnd 0.03294f
C837 vdd.t49 gnd 0.03294f
C838 vdd.n181 gnd 0.226387f
C839 vdd.n182 gnd 0.14366f
C840 vdd.t99 gnd 0.03294f
C841 vdd.t140 gnd 0.03294f
C842 vdd.n183 gnd 0.226387f
C843 vdd.n184 gnd 0.14366f
C844 vdd.t21 gnd 0.03294f
C845 vdd.t47 gnd 0.03294f
C846 vdd.n185 gnd 0.226387f
C847 vdd.n186 gnd 0.14366f
C848 vdd.t132 gnd 0.03294f
C849 vdd.t13 gnd 0.03294f
C850 vdd.n187 gnd 0.226387f
C851 vdd.n188 gnd 0.14366f
C852 vdd.n189 gnd 0.005615f
C853 vdd.n190 gnd 0.005211f
C854 vdd.n191 gnd 0.002882f
C855 vdd.n192 gnd 0.006618f
C856 vdd.n193 gnd 0.0028f
C857 vdd.n194 gnd 0.002965f
C858 vdd.n195 gnd 0.005211f
C859 vdd.n196 gnd 0.0028f
C860 vdd.n197 gnd 0.006618f
C861 vdd.n198 gnd 0.002965f
C862 vdd.n199 gnd 0.005211f
C863 vdd.n200 gnd 0.0028f
C864 vdd.n201 gnd 0.004963f
C865 vdd.n202 gnd 0.004978f
C866 vdd.t15 gnd 0.014218f
C867 vdd.n203 gnd 0.031635f
C868 vdd.n204 gnd 0.164637f
C869 vdd.n205 gnd 0.0028f
C870 vdd.n206 gnd 0.002965f
C871 vdd.n207 gnd 0.006618f
C872 vdd.n208 gnd 0.006618f
C873 vdd.n209 gnd 0.002965f
C874 vdd.n210 gnd 0.0028f
C875 vdd.n211 gnd 0.005211f
C876 vdd.n212 gnd 0.005211f
C877 vdd.n213 gnd 0.0028f
C878 vdd.n214 gnd 0.002965f
C879 vdd.n215 gnd 0.006618f
C880 vdd.n216 gnd 0.006618f
C881 vdd.n217 gnd 0.002965f
C882 vdd.n218 gnd 0.0028f
C883 vdd.n219 gnd 0.005211f
C884 vdd.n220 gnd 0.005211f
C885 vdd.n221 gnd 0.0028f
C886 vdd.n222 gnd 0.002965f
C887 vdd.n223 gnd 0.006618f
C888 vdd.n224 gnd 0.006618f
C889 vdd.n225 gnd 0.015646f
C890 vdd.n226 gnd 0.002882f
C891 vdd.n227 gnd 0.0028f
C892 vdd.n228 gnd 0.013467f
C893 vdd.n229 gnd 0.009107f
C894 vdd.n230 gnd 0.063585f
C895 vdd.n231 gnd 0.229114f
C896 vdd.n232 gnd 0.005615f
C897 vdd.n233 gnd 0.005211f
C898 vdd.n234 gnd 0.002882f
C899 vdd.n235 gnd 0.006618f
C900 vdd.n236 gnd 0.0028f
C901 vdd.n237 gnd 0.002965f
C902 vdd.n238 gnd 0.005211f
C903 vdd.n239 gnd 0.0028f
C904 vdd.n240 gnd 0.006618f
C905 vdd.n241 gnd 0.002965f
C906 vdd.n242 gnd 0.005211f
C907 vdd.n243 gnd 0.0028f
C908 vdd.n244 gnd 0.004963f
C909 vdd.n245 gnd 0.004978f
C910 vdd.t152 gnd 0.014218f
C911 vdd.n246 gnd 0.031635f
C912 vdd.n247 gnd 0.164637f
C913 vdd.n248 gnd 0.0028f
C914 vdd.n249 gnd 0.002965f
C915 vdd.n250 gnd 0.006618f
C916 vdd.n251 gnd 0.006618f
C917 vdd.n252 gnd 0.002965f
C918 vdd.n253 gnd 0.0028f
C919 vdd.n254 gnd 0.005211f
C920 vdd.n255 gnd 0.005211f
C921 vdd.n256 gnd 0.0028f
C922 vdd.n257 gnd 0.002965f
C923 vdd.n258 gnd 0.006618f
C924 vdd.n259 gnd 0.006618f
C925 vdd.n260 gnd 0.002965f
C926 vdd.n261 gnd 0.0028f
C927 vdd.n262 gnd 0.005211f
C928 vdd.n263 gnd 0.005211f
C929 vdd.n264 gnd 0.0028f
C930 vdd.n265 gnd 0.002965f
C931 vdd.n266 gnd 0.006618f
C932 vdd.n267 gnd 0.006618f
C933 vdd.n268 gnd 0.015646f
C934 vdd.n269 gnd 0.002882f
C935 vdd.n270 gnd 0.0028f
C936 vdd.n271 gnd 0.013467f
C937 vdd.n272 gnd 0.009402f
C938 vdd.t154 gnd 0.03294f
C939 vdd.t46 gnd 0.03294f
C940 vdd.n273 gnd 0.226387f
C941 vdd.n274 gnd 0.178019f
C942 vdd.t131 gnd 0.03294f
C943 vdd.t149 gnd 0.03294f
C944 vdd.n275 gnd 0.226387f
C945 vdd.n276 gnd 0.14366f
C946 vdd.t35 gnd 0.03294f
C947 vdd.t101 gnd 0.03294f
C948 vdd.n277 gnd 0.226387f
C949 vdd.n278 gnd 0.14366f
C950 vdd.t130 gnd 0.03294f
C951 vdd.t7 gnd 0.03294f
C952 vdd.n279 gnd 0.226387f
C953 vdd.n280 gnd 0.14366f
C954 vdd.t73 gnd 0.03294f
C955 vdd.t126 gnd 0.03294f
C956 vdd.n281 gnd 0.226387f
C957 vdd.n282 gnd 0.14366f
C958 vdd.t19 gnd 0.03294f
C959 vdd.t71 gnd 0.03294f
C960 vdd.n283 gnd 0.226387f
C961 vdd.n284 gnd 0.14366f
C962 vdd.t109 gnd 0.03294f
C963 vdd.t153 gnd 0.03294f
C964 vdd.n285 gnd 0.226387f
C965 vdd.n286 gnd 0.14366f
C966 vdd.t41 gnd 0.03294f
C967 vdd.t69 gnd 0.03294f
C968 vdd.n287 gnd 0.226387f
C969 vdd.n288 gnd 0.14366f
C970 vdd.t148 gnd 0.03294f
C971 vdd.t31 gnd 0.03294f
C972 vdd.n289 gnd 0.226387f
C973 vdd.n290 gnd 0.14366f
C974 vdd.n291 gnd 0.005615f
C975 vdd.n292 gnd 0.005211f
C976 vdd.n293 gnd 0.002882f
C977 vdd.n294 gnd 0.006618f
C978 vdd.n295 gnd 0.0028f
C979 vdd.n296 gnd 0.002965f
C980 vdd.n297 gnd 0.005211f
C981 vdd.n298 gnd 0.0028f
C982 vdd.n299 gnd 0.006618f
C983 vdd.n300 gnd 0.002965f
C984 vdd.n301 gnd 0.005211f
C985 vdd.n302 gnd 0.0028f
C986 vdd.n303 gnd 0.004963f
C987 vdd.n304 gnd 0.004978f
C988 vdd.t36 gnd 0.014218f
C989 vdd.n305 gnd 0.031635f
C990 vdd.n306 gnd 0.164637f
C991 vdd.n307 gnd 0.0028f
C992 vdd.n308 gnd 0.002965f
C993 vdd.n309 gnd 0.006618f
C994 vdd.n310 gnd 0.006618f
C995 vdd.n311 gnd 0.002965f
C996 vdd.n312 gnd 0.0028f
C997 vdd.n313 gnd 0.005211f
C998 vdd.n314 gnd 0.005211f
C999 vdd.n315 gnd 0.0028f
C1000 vdd.n316 gnd 0.002965f
C1001 vdd.n317 gnd 0.006618f
C1002 vdd.n318 gnd 0.006618f
C1003 vdd.n319 gnd 0.002965f
C1004 vdd.n320 gnd 0.0028f
C1005 vdd.n321 gnd 0.005211f
C1006 vdd.n322 gnd 0.005211f
C1007 vdd.n323 gnd 0.0028f
C1008 vdd.n324 gnd 0.002965f
C1009 vdd.n325 gnd 0.006618f
C1010 vdd.n326 gnd 0.006618f
C1011 vdd.n327 gnd 0.015646f
C1012 vdd.n328 gnd 0.002882f
C1013 vdd.n329 gnd 0.0028f
C1014 vdd.n330 gnd 0.013467f
C1015 vdd.n331 gnd 0.009107f
C1016 vdd.n332 gnd 0.063585f
C1017 vdd.n333 gnd 0.262286f
C1018 vdd.n334 gnd 0.007863f
C1019 vdd.n335 gnd 0.010231f
C1020 vdd.n336 gnd 0.008235f
C1021 vdd.n337 gnd 0.008235f
C1022 vdd.n338 gnd 0.010231f
C1023 vdd.n339 gnd 0.010231f
C1024 vdd.n340 gnd 0.747604f
C1025 vdd.n341 gnd 0.010231f
C1026 vdd.n342 gnd 0.010231f
C1027 vdd.n343 gnd 0.010231f
C1028 vdd.n344 gnd 0.810339f
C1029 vdd.n345 gnd 0.010231f
C1030 vdd.n346 gnd 0.010231f
C1031 vdd.n347 gnd 0.010231f
C1032 vdd.n348 gnd 0.010231f
C1033 vdd.n349 gnd 0.008235f
C1034 vdd.n350 gnd 0.010231f
C1035 vdd.t48 gnd 0.5228f
C1036 vdd.n351 gnd 0.010231f
C1037 vdd.n352 gnd 0.010231f
C1038 vdd.n353 gnd 0.010231f
C1039 vdd.t139 gnd 0.5228f
C1040 vdd.n354 gnd 0.010231f
C1041 vdd.n355 gnd 0.010231f
C1042 vdd.n356 gnd 0.010231f
C1043 vdd.n357 gnd 0.010231f
C1044 vdd.n358 gnd 0.010231f
C1045 vdd.n359 gnd 0.008235f
C1046 vdd.n360 gnd 0.010231f
C1047 vdd.n361 gnd 0.590764f
C1048 vdd.n362 gnd 0.010231f
C1049 vdd.n363 gnd 0.010231f
C1050 vdd.n364 gnd 0.010231f
C1051 vdd.t2 gnd 0.5228f
C1052 vdd.n365 gnd 0.010231f
C1053 vdd.n366 gnd 0.010231f
C1054 vdd.n367 gnd 0.010231f
C1055 vdd.n368 gnd 0.010231f
C1056 vdd.n369 gnd 0.010231f
C1057 vdd.n370 gnd 0.008235f
C1058 vdd.n371 gnd 0.010231f
C1059 vdd.t66 gnd 0.5228f
C1060 vdd.n372 gnd 0.010231f
C1061 vdd.n373 gnd 0.010231f
C1062 vdd.n374 gnd 0.010231f
C1063 vdd.n375 gnd 0.611676f
C1064 vdd.n376 gnd 0.010231f
C1065 vdd.n377 gnd 0.010231f
C1066 vdd.n378 gnd 0.010231f
C1067 vdd.n379 gnd 0.010231f
C1068 vdd.n380 gnd 0.010231f
C1069 vdd.n381 gnd 0.008235f
C1070 vdd.n382 gnd 0.010231f
C1071 vdd.t14 gnd 0.5228f
C1072 vdd.n383 gnd 0.010231f
C1073 vdd.n384 gnd 0.010231f
C1074 vdd.n385 gnd 0.010231f
C1075 vdd.n386 gnd 0.528028f
C1076 vdd.n387 gnd 0.010231f
C1077 vdd.n388 gnd 0.010231f
C1078 vdd.n389 gnd 0.010231f
C1079 vdd.n390 gnd 0.010231f
C1080 vdd.n391 gnd 0.024751f
C1081 vdd.n392 gnd 0.025281f
C1082 vdd.t173 gnd 0.5228f
C1083 vdd.n393 gnd 0.024751f
C1084 vdd.n425 gnd 0.010231f
C1085 vdd.t201 gnd 0.125873f
C1086 vdd.t200 gnd 0.134524f
C1087 vdd.t199 gnd 0.164388f
C1088 vdd.n426 gnd 0.210723f
C1089 vdd.n427 gnd 0.177869f
C1090 vdd.n428 gnd 0.013505f
C1091 vdd.n429 gnd 0.010231f
C1092 vdd.n430 gnd 0.008235f
C1093 vdd.n431 gnd 0.010231f
C1094 vdd.n432 gnd 0.008235f
C1095 vdd.n433 gnd 0.010231f
C1096 vdd.n434 gnd 0.008235f
C1097 vdd.n435 gnd 0.010231f
C1098 vdd.n436 gnd 0.008235f
C1099 vdd.n437 gnd 0.010231f
C1100 vdd.n438 gnd 0.008235f
C1101 vdd.n439 gnd 0.010231f
C1102 vdd.t175 gnd 0.125873f
C1103 vdd.t174 gnd 0.134524f
C1104 vdd.t172 gnd 0.164388f
C1105 vdd.n440 gnd 0.210723f
C1106 vdd.n441 gnd 0.177869f
C1107 vdd.n442 gnd 0.008235f
C1108 vdd.n443 gnd 0.010231f
C1109 vdd.n444 gnd 0.008235f
C1110 vdd.n445 gnd 0.010231f
C1111 vdd.n446 gnd 0.008235f
C1112 vdd.n447 gnd 0.010231f
C1113 vdd.n448 gnd 0.008235f
C1114 vdd.n449 gnd 0.010231f
C1115 vdd.n450 gnd 0.008235f
C1116 vdd.n451 gnd 0.010231f
C1117 vdd.t181 gnd 0.125873f
C1118 vdd.t180 gnd 0.134524f
C1119 vdd.t179 gnd 0.164388f
C1120 vdd.n452 gnd 0.210723f
C1121 vdd.n453 gnd 0.177869f
C1122 vdd.n454 gnd 0.017623f
C1123 vdd.n455 gnd 0.010231f
C1124 vdd.n456 gnd 0.008235f
C1125 vdd.n457 gnd 0.010231f
C1126 vdd.n458 gnd 0.008235f
C1127 vdd.n459 gnd 0.010231f
C1128 vdd.n460 gnd 0.008235f
C1129 vdd.n461 gnd 0.010231f
C1130 vdd.n462 gnd 0.008235f
C1131 vdd.n463 gnd 0.010231f
C1132 vdd.n464 gnd 0.025281f
C1133 vdd.n465 gnd 0.006835f
C1134 vdd.n466 gnd 0.008235f
C1135 vdd.n467 gnd 0.010231f
C1136 vdd.n468 gnd 0.010231f
C1137 vdd.n469 gnd 0.008235f
C1138 vdd.n470 gnd 0.010231f
C1139 vdd.n471 gnd 0.010231f
C1140 vdd.n472 gnd 0.010231f
C1141 vdd.n473 gnd 0.010231f
C1142 vdd.n474 gnd 0.010231f
C1143 vdd.n475 gnd 0.008235f
C1144 vdd.n476 gnd 0.008235f
C1145 vdd.n477 gnd 0.010231f
C1146 vdd.n478 gnd 0.010231f
C1147 vdd.n479 gnd 0.008235f
C1148 vdd.n480 gnd 0.010231f
C1149 vdd.n481 gnd 0.010231f
C1150 vdd.n482 gnd 0.010231f
C1151 vdd.n483 gnd 0.010231f
C1152 vdd.n484 gnd 0.010231f
C1153 vdd.n485 gnd 0.008235f
C1154 vdd.n486 gnd 0.008235f
C1155 vdd.n487 gnd 0.010231f
C1156 vdd.n488 gnd 0.010231f
C1157 vdd.n489 gnd 0.008235f
C1158 vdd.n490 gnd 0.010231f
C1159 vdd.n491 gnd 0.010231f
C1160 vdd.n492 gnd 0.010231f
C1161 vdd.n493 gnd 0.010231f
C1162 vdd.n494 gnd 0.010231f
C1163 vdd.n495 gnd 0.008235f
C1164 vdd.n496 gnd 0.008235f
C1165 vdd.n497 gnd 0.010231f
C1166 vdd.n498 gnd 0.010231f
C1167 vdd.n499 gnd 0.008235f
C1168 vdd.n500 gnd 0.010231f
C1169 vdd.n501 gnd 0.010231f
C1170 vdd.n502 gnd 0.010231f
C1171 vdd.n503 gnd 0.010231f
C1172 vdd.n504 gnd 0.010231f
C1173 vdd.n505 gnd 0.008235f
C1174 vdd.n506 gnd 0.008235f
C1175 vdd.n507 gnd 0.010231f
C1176 vdd.n508 gnd 0.010231f
C1177 vdd.n509 gnd 0.006876f
C1178 vdd.n510 gnd 0.010231f
C1179 vdd.n511 gnd 0.010231f
C1180 vdd.n512 gnd 0.010231f
C1181 vdd.n513 gnd 0.010231f
C1182 vdd.n514 gnd 0.010231f
C1183 vdd.n515 gnd 0.006876f
C1184 vdd.n516 gnd 0.008235f
C1185 vdd.n517 gnd 0.010231f
C1186 vdd.n518 gnd 0.010231f
C1187 vdd.n519 gnd 0.008235f
C1188 vdd.n520 gnd 0.010231f
C1189 vdd.n521 gnd 0.010231f
C1190 vdd.n522 gnd 0.010231f
C1191 vdd.n523 gnd 0.010231f
C1192 vdd.n524 gnd 0.010231f
C1193 vdd.n525 gnd 0.008235f
C1194 vdd.n526 gnd 0.008235f
C1195 vdd.n527 gnd 0.010231f
C1196 vdd.n528 gnd 0.010231f
C1197 vdd.n529 gnd 0.008235f
C1198 vdd.n530 gnd 0.010231f
C1199 vdd.n531 gnd 0.010231f
C1200 vdd.n532 gnd 0.010231f
C1201 vdd.n533 gnd 0.010231f
C1202 vdd.n534 gnd 0.010231f
C1203 vdd.n535 gnd 0.008235f
C1204 vdd.n536 gnd 0.008235f
C1205 vdd.n537 gnd 0.010231f
C1206 vdd.n538 gnd 0.010231f
C1207 vdd.n539 gnd 0.008235f
C1208 vdd.n540 gnd 0.010231f
C1209 vdd.n541 gnd 0.010231f
C1210 vdd.n542 gnd 0.010231f
C1211 vdd.n543 gnd 0.010231f
C1212 vdd.n544 gnd 0.010231f
C1213 vdd.n545 gnd 0.008235f
C1214 vdd.n546 gnd 0.008235f
C1215 vdd.n547 gnd 0.010231f
C1216 vdd.n548 gnd 0.010231f
C1217 vdd.n549 gnd 0.008235f
C1218 vdd.n550 gnd 0.010231f
C1219 vdd.n551 gnd 0.010231f
C1220 vdd.n552 gnd 0.010231f
C1221 vdd.n553 gnd 0.010231f
C1222 vdd.n554 gnd 0.010231f
C1223 vdd.n555 gnd 0.008235f
C1224 vdd.n556 gnd 0.008235f
C1225 vdd.n557 gnd 0.010231f
C1226 vdd.n558 gnd 0.010231f
C1227 vdd.n559 gnd 0.008235f
C1228 vdd.n560 gnd 0.010231f
C1229 vdd.n561 gnd 0.010231f
C1230 vdd.n562 gnd 0.010231f
C1231 vdd.n563 gnd 0.010231f
C1232 vdd.n564 gnd 0.010231f
C1233 vdd.n565 gnd 0.0056f
C1234 vdd.n566 gnd 0.017623f
C1235 vdd.n567 gnd 0.010231f
C1236 vdd.n568 gnd 0.010231f
C1237 vdd.n569 gnd 0.008153f
C1238 vdd.n570 gnd 0.010231f
C1239 vdd.n571 gnd 0.010231f
C1240 vdd.n572 gnd 0.010231f
C1241 vdd.n573 gnd 0.010231f
C1242 vdd.n574 gnd 0.010231f
C1243 vdd.n575 gnd 0.008235f
C1244 vdd.n576 gnd 0.008235f
C1245 vdd.n577 gnd 0.010231f
C1246 vdd.n578 gnd 0.010231f
C1247 vdd.n579 gnd 0.008235f
C1248 vdd.n580 gnd 0.010231f
C1249 vdd.n581 gnd 0.010231f
C1250 vdd.n582 gnd 0.010231f
C1251 vdd.n583 gnd 0.010231f
C1252 vdd.n584 gnd 0.010231f
C1253 vdd.n585 gnd 0.008235f
C1254 vdd.n586 gnd 0.008235f
C1255 vdd.n587 gnd 0.010231f
C1256 vdd.n588 gnd 0.010231f
C1257 vdd.n589 gnd 0.008235f
C1258 vdd.n590 gnd 0.010231f
C1259 vdd.n591 gnd 0.010231f
C1260 vdd.n592 gnd 0.010231f
C1261 vdd.n593 gnd 0.010231f
C1262 vdd.n594 gnd 0.010231f
C1263 vdd.n595 gnd 0.008235f
C1264 vdd.n596 gnd 0.008235f
C1265 vdd.n597 gnd 0.010231f
C1266 vdd.n598 gnd 0.010231f
C1267 vdd.n599 gnd 0.008235f
C1268 vdd.n600 gnd 0.010231f
C1269 vdd.n601 gnd 0.010231f
C1270 vdd.n602 gnd 0.010231f
C1271 vdd.n603 gnd 0.010231f
C1272 vdd.n604 gnd 0.010231f
C1273 vdd.n605 gnd 0.008235f
C1274 vdd.n606 gnd 0.008235f
C1275 vdd.n607 gnd 0.010231f
C1276 vdd.n608 gnd 0.010231f
C1277 vdd.n609 gnd 0.008235f
C1278 vdd.n610 gnd 0.010231f
C1279 vdd.n611 gnd 0.010231f
C1280 vdd.n612 gnd 0.010231f
C1281 vdd.n613 gnd 0.010231f
C1282 vdd.n614 gnd 0.010231f
C1283 vdd.n615 gnd 0.008235f
C1284 vdd.n616 gnd 0.010231f
C1285 vdd.n617 gnd 0.008235f
C1286 vdd.n618 gnd 0.004323f
C1287 vdd.n619 gnd 0.010231f
C1288 vdd.n620 gnd 0.010231f
C1289 vdd.n621 gnd 0.008235f
C1290 vdd.n622 gnd 0.010231f
C1291 vdd.n623 gnd 0.008235f
C1292 vdd.n624 gnd 0.010231f
C1293 vdd.n625 gnd 0.008235f
C1294 vdd.n626 gnd 0.010231f
C1295 vdd.n627 gnd 0.008235f
C1296 vdd.n628 gnd 0.010231f
C1297 vdd.n629 gnd 0.008235f
C1298 vdd.n630 gnd 0.010231f
C1299 vdd.n631 gnd 0.008235f
C1300 vdd.n632 gnd 0.010231f
C1301 vdd.n633 gnd 0.569852f
C1302 vdd.t56 gnd 0.5228f
C1303 vdd.n634 gnd 0.010231f
C1304 vdd.n635 gnd 0.008235f
C1305 vdd.n636 gnd 0.010231f
C1306 vdd.n637 gnd 0.008235f
C1307 vdd.n638 gnd 0.010231f
C1308 vdd.t64 gnd 0.5228f
C1309 vdd.n639 gnd 0.010231f
C1310 vdd.n640 gnd 0.008235f
C1311 vdd.n641 gnd 0.010231f
C1312 vdd.n642 gnd 0.008235f
C1313 vdd.n643 gnd 0.010231f
C1314 vdd.t79 gnd 0.5228f
C1315 vdd.n644 gnd 0.6535f
C1316 vdd.n645 gnd 0.010231f
C1317 vdd.n646 gnd 0.008235f
C1318 vdd.n647 gnd 0.010231f
C1319 vdd.n648 gnd 0.008235f
C1320 vdd.n649 gnd 0.010231f
C1321 vdd.t16 gnd 0.5228f
C1322 vdd.n650 gnd 0.010231f
C1323 vdd.n651 gnd 0.008235f
C1324 vdd.n652 gnd 0.010231f
C1325 vdd.n653 gnd 0.008235f
C1326 vdd.n654 gnd 0.010231f
C1327 vdd.n655 gnd 0.726692f
C1328 vdd.n656 gnd 0.867847f
C1329 vdd.t112 gnd 0.5228f
C1330 vdd.n657 gnd 0.010231f
C1331 vdd.n658 gnd 0.008235f
C1332 vdd.n659 gnd 0.010231f
C1333 vdd.n660 gnd 0.008235f
C1334 vdd.n661 gnd 0.010231f
C1335 vdd.n662 gnd 0.54894f
C1336 vdd.n663 gnd 0.010231f
C1337 vdd.n664 gnd 0.008235f
C1338 vdd.n665 gnd 0.010231f
C1339 vdd.n666 gnd 0.008235f
C1340 vdd.n667 gnd 0.010231f
C1341 vdd.t50 gnd 0.5228f
C1342 vdd.t22 gnd 0.5228f
C1343 vdd.n668 gnd 0.010231f
C1344 vdd.n669 gnd 0.008235f
C1345 vdd.n670 gnd 0.010231f
C1346 vdd.n671 gnd 0.008235f
C1347 vdd.n672 gnd 0.010231f
C1348 vdd.t81 gnd 0.5228f
C1349 vdd.n673 gnd 0.010231f
C1350 vdd.n674 gnd 0.008235f
C1351 vdd.n675 gnd 0.010231f
C1352 vdd.n676 gnd 0.008235f
C1353 vdd.n677 gnd 0.010231f
C1354 vdd.n678 gnd 1.0456f
C1355 vdd.n679 gnd 0.852163f
C1356 vdd.n680 gnd 0.010231f
C1357 vdd.n681 gnd 0.008235f
C1358 vdd.n682 gnd 0.024751f
C1359 vdd.n683 gnd 0.006835f
C1360 vdd.n684 gnd 0.024751f
C1361 vdd.t186 gnd 0.5228f
C1362 vdd.n685 gnd 0.024751f
C1363 vdd.n686 gnd 0.006835f
C1364 vdd.n687 gnd 0.008799f
C1365 vdd.t187 gnd 0.125873f
C1366 vdd.t188 gnd 0.134524f
C1367 vdd.t185 gnd 0.164388f
C1368 vdd.n688 gnd 0.210723f
C1369 vdd.n689 gnd 0.177045f
C1370 vdd.n690 gnd 0.012682f
C1371 vdd.n691 gnd 0.010231f
C1372 vdd.n692 gnd 12.3485f
C1373 vdd.n723 gnd 1.4377f
C1374 vdd.n724 gnd 0.010231f
C1375 vdd.n725 gnd 0.010231f
C1376 vdd.n726 gnd 0.025281f
C1377 vdd.n727 gnd 0.008799f
C1378 vdd.n728 gnd 0.010231f
C1379 vdd.n729 gnd 0.008235f
C1380 vdd.n730 gnd 0.006548f
C1381 vdd.n731 gnd 0.042961f
C1382 vdd.n732 gnd 0.008235f
C1383 vdd.n733 gnd 0.010231f
C1384 vdd.n734 gnd 0.010231f
C1385 vdd.n735 gnd 0.010231f
C1386 vdd.n736 gnd 0.010231f
C1387 vdd.n737 gnd 0.010231f
C1388 vdd.n738 gnd 0.010231f
C1389 vdd.n739 gnd 0.010231f
C1390 vdd.n740 gnd 0.010231f
C1391 vdd.n741 gnd 0.010231f
C1392 vdd.n742 gnd 0.010231f
C1393 vdd.n743 gnd 0.010231f
C1394 vdd.n744 gnd 0.010231f
C1395 vdd.n745 gnd 0.010231f
C1396 vdd.n746 gnd 0.010231f
C1397 vdd.n747 gnd 0.006876f
C1398 vdd.n748 gnd 0.010231f
C1399 vdd.n749 gnd 0.010231f
C1400 vdd.n750 gnd 0.010231f
C1401 vdd.n751 gnd 0.010231f
C1402 vdd.n752 gnd 0.010231f
C1403 vdd.n753 gnd 0.010231f
C1404 vdd.n754 gnd 0.010231f
C1405 vdd.n755 gnd 0.010231f
C1406 vdd.n756 gnd 0.010231f
C1407 vdd.n757 gnd 0.010231f
C1408 vdd.n758 gnd 0.010231f
C1409 vdd.n759 gnd 0.010231f
C1410 vdd.n760 gnd 0.010231f
C1411 vdd.n761 gnd 0.010231f
C1412 vdd.n762 gnd 0.010231f
C1413 vdd.n763 gnd 0.010231f
C1414 vdd.n764 gnd 0.010231f
C1415 vdd.n765 gnd 0.010231f
C1416 vdd.n766 gnd 0.010231f
C1417 vdd.n767 gnd 0.008153f
C1418 vdd.t197 gnd 0.125873f
C1419 vdd.t198 gnd 0.134524f
C1420 vdd.t196 gnd 0.164388f
C1421 vdd.n768 gnd 0.210723f
C1422 vdd.n769 gnd 0.177045f
C1423 vdd.n770 gnd 0.010231f
C1424 vdd.n771 gnd 0.010231f
C1425 vdd.n772 gnd 0.010231f
C1426 vdd.n773 gnd 0.010231f
C1427 vdd.n774 gnd 0.010231f
C1428 vdd.n775 gnd 0.010231f
C1429 vdd.n776 gnd 0.010231f
C1430 vdd.n777 gnd 0.010231f
C1431 vdd.n778 gnd 0.010231f
C1432 vdd.n779 gnd 0.010231f
C1433 vdd.n780 gnd 0.010231f
C1434 vdd.n781 gnd 0.010231f
C1435 vdd.n782 gnd 0.010231f
C1436 vdd.n783 gnd 0.006548f
C1437 vdd.n785 gnd 0.006957f
C1438 vdd.n786 gnd 0.006957f
C1439 vdd.n787 gnd 0.006957f
C1440 vdd.n788 gnd 0.006957f
C1441 vdd.n789 gnd 0.006957f
C1442 vdd.n790 gnd 0.006957f
C1443 vdd.n792 gnd 0.006957f
C1444 vdd.n793 gnd 0.006957f
C1445 vdd.n795 gnd 0.006957f
C1446 vdd.n796 gnd 0.005065f
C1447 vdd.n798 gnd 0.006957f
C1448 vdd.t163 gnd 0.281145f
C1449 vdd.t162 gnd 0.287787f
C1450 vdd.t160 gnd 0.183542f
C1451 vdd.n799 gnd 0.099195f
C1452 vdd.n800 gnd 0.056266f
C1453 vdd.n801 gnd 0.009943f
C1454 vdd.n802 gnd 0.015797f
C1455 vdd.n804 gnd 0.006957f
C1456 vdd.n805 gnd 0.711008f
C1457 vdd.n806 gnd 0.014897f
C1458 vdd.n807 gnd 0.014897f
C1459 vdd.n808 gnd 0.006957f
C1460 vdd.n809 gnd 0.015797f
C1461 vdd.n810 gnd 0.006957f
C1462 vdd.n811 gnd 0.006957f
C1463 vdd.n812 gnd 0.006957f
C1464 vdd.n813 gnd 0.006957f
C1465 vdd.n814 gnd 0.006957f
C1466 vdd.n816 gnd 0.006957f
C1467 vdd.n817 gnd 0.006957f
C1468 vdd.n819 gnd 0.006957f
C1469 vdd.n820 gnd 0.006957f
C1470 vdd.n822 gnd 0.006957f
C1471 vdd.n823 gnd 0.006957f
C1472 vdd.n825 gnd 0.006957f
C1473 vdd.n826 gnd 0.006957f
C1474 vdd.n828 gnd 0.006957f
C1475 vdd.n829 gnd 0.006957f
C1476 vdd.n831 gnd 0.006957f
C1477 vdd.t184 gnd 0.281145f
C1478 vdd.t183 gnd 0.287787f
C1479 vdd.t182 gnd 0.183542f
C1480 vdd.n832 gnd 0.099195f
C1481 vdd.n833 gnd 0.056266f
C1482 vdd.n834 gnd 0.006957f
C1483 vdd.n836 gnd 0.006957f
C1484 vdd.n837 gnd 0.006957f
C1485 vdd.t161 gnd 0.355504f
C1486 vdd.n838 gnd 0.006957f
C1487 vdd.n839 gnd 0.006957f
C1488 vdd.n840 gnd 0.006957f
C1489 vdd.n841 gnd 0.006957f
C1490 vdd.n842 gnd 0.006957f
C1491 vdd.n843 gnd 0.711008f
C1492 vdd.n844 gnd 0.006957f
C1493 vdd.n845 gnd 0.006957f
C1494 vdd.n846 gnd 0.559396f
C1495 vdd.n847 gnd 0.006957f
C1496 vdd.n848 gnd 0.006957f
C1497 vdd.n849 gnd 0.006957f
C1498 vdd.n850 gnd 0.006957f
C1499 vdd.n851 gnd 0.711008f
C1500 vdd.n852 gnd 0.006957f
C1501 vdd.n853 gnd 0.006957f
C1502 vdd.n854 gnd 0.006957f
C1503 vdd.n855 gnd 0.006957f
C1504 vdd.n856 gnd 0.006957f
C1505 vdd.t250 gnd 0.355504f
C1506 vdd.n857 gnd 0.006957f
C1507 vdd.n858 gnd 0.006957f
C1508 vdd.n859 gnd 0.006957f
C1509 vdd.n860 gnd 0.006957f
C1510 vdd.n861 gnd 0.006957f
C1511 vdd.t267 gnd 0.355504f
C1512 vdd.n862 gnd 0.006957f
C1513 vdd.n863 gnd 0.006957f
C1514 vdd.n864 gnd 0.684868f
C1515 vdd.n865 gnd 0.006957f
C1516 vdd.n866 gnd 0.006957f
C1517 vdd.n867 gnd 0.006957f
C1518 vdd.t266 gnd 0.355504f
C1519 vdd.n868 gnd 0.006957f
C1520 vdd.n869 gnd 0.006957f
C1521 vdd.n870 gnd 0.528028f
C1522 vdd.n871 gnd 0.006957f
C1523 vdd.n872 gnd 0.006957f
C1524 vdd.n873 gnd 0.006957f
C1525 vdd.n874 gnd 0.49666f
C1526 vdd.n875 gnd 0.006957f
C1527 vdd.n876 gnd 0.006957f
C1528 vdd.n877 gnd 0.371188f
C1529 vdd.n878 gnd 0.006957f
C1530 vdd.n879 gnd 0.006957f
C1531 vdd.n880 gnd 0.006957f
C1532 vdd.n881 gnd 0.6535f
C1533 vdd.n882 gnd 0.006957f
C1534 vdd.n883 gnd 0.006957f
C1535 vdd.t273 gnd 0.355504f
C1536 vdd.n884 gnd 0.006957f
C1537 vdd.n885 gnd 0.006957f
C1538 vdd.n886 gnd 0.006957f
C1539 vdd.n887 gnd 0.711008f
C1540 vdd.n888 gnd 0.006957f
C1541 vdd.n889 gnd 0.006957f
C1542 vdd.t274 gnd 0.355504f
C1543 vdd.n890 gnd 0.006957f
C1544 vdd.n891 gnd 0.006957f
C1545 vdd.n892 gnd 0.006957f
C1546 vdd.t244 gnd 0.355504f
C1547 vdd.n893 gnd 0.006957f
C1548 vdd.n894 gnd 0.006957f
C1549 vdd.n895 gnd 0.006957f
C1550 vdd.t191 gnd 0.287787f
C1551 vdd.t189 gnd 0.183542f
C1552 vdd.t192 gnd 0.287787f
C1553 vdd.n896 gnd 0.161748f
C1554 vdd.n897 gnd 0.020155f
C1555 vdd.n898 gnd 0.006957f
C1556 vdd.t190 gnd 0.256172f
C1557 vdd.n899 gnd 0.006957f
C1558 vdd.n900 gnd 0.006957f
C1559 vdd.n901 gnd 0.611676f
C1560 vdd.n902 gnd 0.006957f
C1561 vdd.n903 gnd 0.006957f
C1562 vdd.n904 gnd 0.006957f
C1563 vdd.n905 gnd 0.413012f
C1564 vdd.n906 gnd 0.006957f
C1565 vdd.n907 gnd 0.006957f
C1566 vdd.t245 gnd 0.146384f
C1567 vdd.n908 gnd 0.454836f
C1568 vdd.n909 gnd 0.006957f
C1569 vdd.n910 gnd 0.006957f
C1570 vdd.n911 gnd 0.006957f
C1571 vdd.n912 gnd 0.569852f
C1572 vdd.n913 gnd 0.006957f
C1573 vdd.n914 gnd 0.006957f
C1574 vdd.t258 gnd 0.355504f
C1575 vdd.n915 gnd 0.006957f
C1576 vdd.n916 gnd 0.006957f
C1577 vdd.n917 gnd 0.006957f
C1578 vdd.t254 gnd 0.355504f
C1579 vdd.n918 gnd 0.006957f
C1580 vdd.n919 gnd 0.006957f
C1581 vdd.t277 gnd 0.355504f
C1582 vdd.n920 gnd 0.006957f
C1583 vdd.n921 gnd 0.006957f
C1584 vdd.n922 gnd 0.006957f
C1585 vdd.t236 gnd 0.240488f
C1586 vdd.n923 gnd 0.006957f
C1587 vdd.n924 gnd 0.006957f
C1588 vdd.n925 gnd 0.62736f
C1589 vdd.n926 gnd 0.006957f
C1590 vdd.n927 gnd 0.006957f
C1591 vdd.n928 gnd 0.006957f
C1592 vdd.t278 gnd 0.355504f
C1593 vdd.n929 gnd 0.006957f
C1594 vdd.n930 gnd 0.006957f
C1595 vdd.t290 gnd 0.33982f
C1596 vdd.n931 gnd 0.47052f
C1597 vdd.n932 gnd 0.006957f
C1598 vdd.n933 gnd 0.006957f
C1599 vdd.n934 gnd 0.006957f
C1600 vdd.t240 gnd 0.355504f
C1601 vdd.n935 gnd 0.006957f
C1602 vdd.n936 gnd 0.006957f
C1603 vdd.t284 gnd 0.355504f
C1604 vdd.n937 gnd 0.006957f
C1605 vdd.n938 gnd 0.006957f
C1606 vdd.n939 gnd 0.006957f
C1607 vdd.n940 gnd 0.711008f
C1608 vdd.n941 gnd 0.006957f
C1609 vdd.n942 gnd 0.006957f
C1610 vdd.t262 gnd 0.355504f
C1611 vdd.n943 gnd 0.006957f
C1612 vdd.n944 gnd 0.006957f
C1613 vdd.n945 gnd 0.006957f
C1614 vdd.n946 gnd 0.491432f
C1615 vdd.n947 gnd 0.006957f
C1616 vdd.n948 gnd 0.006957f
C1617 vdd.n949 gnd 0.006957f
C1618 vdd.n950 gnd 0.006957f
C1619 vdd.n951 gnd 0.006957f
C1620 vdd.t213 gnd 0.355504f
C1621 vdd.n952 gnd 0.006957f
C1622 vdd.n953 gnd 0.006957f
C1623 vdd.t242 gnd 0.355504f
C1624 vdd.n954 gnd 0.006957f
C1625 vdd.n955 gnd 0.014897f
C1626 vdd.n956 gnd 0.014897f
C1627 vdd.n957 gnd 0.805111f
C1628 vdd.n958 gnd 0.006957f
C1629 vdd.n959 gnd 0.006957f
C1630 vdd.t271 gnd 0.355504f
C1631 vdd.n960 gnd 0.014897f
C1632 vdd.n961 gnd 0.006957f
C1633 vdd.n962 gnd 0.006957f
C1634 vdd.t286 gnd 0.606448f
C1635 vdd.n980 gnd 0.015797f
C1636 vdd.n998 gnd 0.014897f
C1637 vdd.n999 gnd 0.006957f
C1638 vdd.n1000 gnd 0.014897f
C1639 vdd.t229 gnd 0.281145f
C1640 vdd.t228 gnd 0.287787f
C1641 vdd.t227 gnd 0.183542f
C1642 vdd.n1001 gnd 0.099195f
C1643 vdd.n1002 gnd 0.056266f
C1644 vdd.n1003 gnd 0.015797f
C1645 vdd.n1004 gnd 0.006957f
C1646 vdd.n1005 gnd 0.41824f
C1647 vdd.n1006 gnd 0.014897f
C1648 vdd.n1007 gnd 0.006957f
C1649 vdd.n1008 gnd 0.015797f
C1650 vdd.n1009 gnd 0.006957f
C1651 vdd.t208 gnd 0.281145f
C1652 vdd.t207 gnd 0.287787f
C1653 vdd.t205 gnd 0.183542f
C1654 vdd.n1010 gnd 0.099195f
C1655 vdd.n1011 gnd 0.056266f
C1656 vdd.n1012 gnd 0.009943f
C1657 vdd.n1013 gnd 0.006957f
C1658 vdd.n1014 gnd 0.006957f
C1659 vdd.t206 gnd 0.355504f
C1660 vdd.n1015 gnd 0.006957f
C1661 vdd.t281 gnd 0.355504f
C1662 vdd.n1016 gnd 0.006957f
C1663 vdd.n1017 gnd 0.006957f
C1664 vdd.n1018 gnd 0.006957f
C1665 vdd.n1019 gnd 0.006957f
C1666 vdd.n1020 gnd 0.006957f
C1667 vdd.n1021 gnd 0.711008f
C1668 vdd.n1022 gnd 0.006957f
C1669 vdd.n1023 gnd 0.006957f
C1670 vdd.t256 gnd 0.355504f
C1671 vdd.n1024 gnd 0.006957f
C1672 vdd.n1025 gnd 0.006957f
C1673 vdd.n1026 gnd 0.006957f
C1674 vdd.n1027 gnd 0.006957f
C1675 vdd.n1028 gnd 0.512344f
C1676 vdd.n1029 gnd 0.006957f
C1677 vdd.n1030 gnd 0.006957f
C1678 vdd.n1031 gnd 0.006957f
C1679 vdd.n1032 gnd 0.006957f
C1680 vdd.n1033 gnd 0.006957f
C1681 vdd.t237 gnd 0.355504f
C1682 vdd.n1034 gnd 0.006957f
C1683 vdd.n1035 gnd 0.006957f
C1684 vdd.t275 gnd 0.355504f
C1685 vdd.n1036 gnd 0.006957f
C1686 vdd.n1037 gnd 0.006957f
C1687 vdd.n1038 gnd 0.006957f
C1688 vdd.t259 gnd 0.355504f
C1689 vdd.n1039 gnd 0.006957f
C1690 vdd.n1040 gnd 0.006957f
C1691 vdd.t238 gnd 0.355504f
C1692 vdd.n1041 gnd 0.006957f
C1693 vdd.n1042 gnd 0.006957f
C1694 vdd.n1043 gnd 0.006957f
C1695 vdd.t260 gnd 0.33982f
C1696 vdd.n1044 gnd 0.006957f
C1697 vdd.n1045 gnd 0.006957f
C1698 vdd.n1046 gnd 0.528028f
C1699 vdd.n1047 gnd 0.006957f
C1700 vdd.n1048 gnd 0.006957f
C1701 vdd.n1049 gnd 0.006957f
C1702 vdd.t279 gnd 0.355504f
C1703 vdd.n1050 gnd 0.006957f
C1704 vdd.n1051 gnd 0.006957f
C1705 vdd.t247 gnd 0.240488f
C1706 vdd.n1052 gnd 0.371188f
C1707 vdd.n1053 gnd 0.006957f
C1708 vdd.n1054 gnd 0.006957f
C1709 vdd.n1055 gnd 0.006957f
C1710 vdd.n1056 gnd 0.6535f
C1711 vdd.n1057 gnd 0.006957f
C1712 vdd.n1058 gnd 0.006957f
C1713 vdd.t288 gnd 0.355504f
C1714 vdd.n1059 gnd 0.006957f
C1715 vdd.n1060 gnd 0.006957f
C1716 vdd.n1061 gnd 0.006957f
C1717 vdd.n1062 gnd 0.711008f
C1718 vdd.n1063 gnd 0.006957f
C1719 vdd.n1064 gnd 0.006957f
C1720 vdd.t253 gnd 0.355504f
C1721 vdd.n1065 gnd 0.006957f
C1722 vdd.n1066 gnd 0.006957f
C1723 vdd.n1067 gnd 0.006957f
C1724 vdd.t246 gnd 0.146384f
C1725 vdd.n1068 gnd 0.006957f
C1726 vdd.n1069 gnd 0.006957f
C1727 vdd.n1070 gnd 0.006957f
C1728 vdd.t218 gnd 0.287787f
C1729 vdd.t216 gnd 0.183542f
C1730 vdd.t219 gnd 0.287787f
C1731 vdd.n1071 gnd 0.161748f
C1732 vdd.n1072 gnd 0.006957f
C1733 vdd.n1073 gnd 0.006957f
C1734 vdd.t268 gnd 0.355504f
C1735 vdd.n1074 gnd 0.006957f
C1736 vdd.n1075 gnd 0.006957f
C1737 vdd.t217 gnd 0.256172f
C1738 vdd.n1076 gnd 0.564624f
C1739 vdd.n1077 gnd 0.006957f
C1740 vdd.n1078 gnd 0.006957f
C1741 vdd.n1079 gnd 0.006957f
C1742 vdd.n1080 gnd 0.413012f
C1743 vdd.n1081 gnd 0.006957f
C1744 vdd.n1082 gnd 0.006957f
C1745 vdd.n1083 gnd 0.454836f
C1746 vdd.n1084 gnd 0.006957f
C1747 vdd.n1085 gnd 0.006957f
C1748 vdd.n1086 gnd 0.006957f
C1749 vdd.n1087 gnd 0.569852f
C1750 vdd.n1088 gnd 0.006957f
C1751 vdd.n1089 gnd 0.006957f
C1752 vdd.t248 gnd 0.355504f
C1753 vdd.n1090 gnd 0.006957f
C1754 vdd.n1091 gnd 0.006957f
C1755 vdd.n1092 gnd 0.006957f
C1756 vdd.n1093 gnd 0.711008f
C1757 vdd.n1094 gnd 0.006957f
C1758 vdd.n1095 gnd 0.006957f
C1759 vdd.t249 gnd 0.355504f
C1760 vdd.n1096 gnd 0.006957f
C1761 vdd.n1097 gnd 0.006957f
C1762 vdd.n1098 gnd 0.006957f
C1763 vdd.t289 gnd 0.355504f
C1764 vdd.n1099 gnd 0.006957f
C1765 vdd.n1100 gnd 0.006957f
C1766 vdd.n1101 gnd 0.006957f
C1767 vdd.n1102 gnd 0.006957f
C1768 vdd.n1103 gnd 0.006957f
C1769 vdd.t283 gnd 0.355504f
C1770 vdd.n1104 gnd 0.006957f
C1771 vdd.n1105 gnd 0.006957f
C1772 vdd.n1106 gnd 0.695324f
C1773 vdd.n1107 gnd 0.006957f
C1774 vdd.n1108 gnd 0.006957f
C1775 vdd.n1109 gnd 0.006957f
C1776 vdd.t241 gnd 0.355504f
C1777 vdd.n1110 gnd 0.006957f
C1778 vdd.n1111 gnd 0.006957f
C1779 vdd.n1112 gnd 0.538484f
C1780 vdd.n1113 gnd 0.006957f
C1781 vdd.n1114 gnd 0.006957f
C1782 vdd.n1115 gnd 0.006957f
C1783 vdd.n1116 gnd 0.711008f
C1784 vdd.n1117 gnd 0.006957f
C1785 vdd.n1118 gnd 0.006957f
C1786 vdd.n1119 gnd 0.381644f
C1787 vdd.n1120 gnd 0.006957f
C1788 vdd.n1121 gnd 0.006957f
C1789 vdd.n1122 gnd 0.006957f
C1790 vdd.n1123 gnd 0.711008f
C1791 vdd.n1124 gnd 0.006957f
C1792 vdd.n1125 gnd 0.006957f
C1793 vdd.n1126 gnd 0.006957f
C1794 vdd.n1127 gnd 0.006957f
C1795 vdd.n1128 gnd 0.006957f
C1796 vdd.t165 gnd 0.355504f
C1797 vdd.n1129 gnd 0.006957f
C1798 vdd.n1130 gnd 0.006957f
C1799 vdd.n1131 gnd 0.006957f
C1800 vdd.n1132 gnd 0.014897f
C1801 vdd.n1133 gnd 0.014897f
C1802 vdd.n1134 gnd 0.961951f
C1803 vdd.n1135 gnd 0.006957f
C1804 vdd.n1136 gnd 0.006957f
C1805 vdd.n1137 gnd 0.507116f
C1806 vdd.n1138 gnd 0.014897f
C1807 vdd.n1139 gnd 0.006957f
C1808 vdd.n1140 gnd 0.006957f
C1809 vdd.n1141 gnd 12.7668f
C1810 vdd.n1175 gnd 0.015797f
C1811 vdd.n1176 gnd 0.006957f
C1812 vdd.n1177 gnd 0.006957f
C1813 vdd.n1178 gnd 0.006548f
C1814 vdd.n1181 gnd 0.025281f
C1815 vdd.n1182 gnd 0.006835f
C1816 vdd.n1183 gnd 0.008235f
C1817 vdd.n1185 gnd 0.010231f
C1818 vdd.n1186 gnd 0.010231f
C1819 vdd.n1187 gnd 0.008235f
C1820 vdd.n1189 gnd 0.010231f
C1821 vdd.n1190 gnd 0.010231f
C1822 vdd.n1191 gnd 0.010231f
C1823 vdd.n1192 gnd 0.010231f
C1824 vdd.n1193 gnd 0.010231f
C1825 vdd.n1194 gnd 0.008235f
C1826 vdd.n1196 gnd 0.010231f
C1827 vdd.n1197 gnd 0.010231f
C1828 vdd.n1198 gnd 0.010231f
C1829 vdd.n1199 gnd 0.010231f
C1830 vdd.n1200 gnd 0.010231f
C1831 vdd.n1201 gnd 0.008235f
C1832 vdd.n1203 gnd 0.010231f
C1833 vdd.n1204 gnd 0.010231f
C1834 vdd.n1205 gnd 0.010231f
C1835 vdd.n1206 gnd 0.010231f
C1836 vdd.n1207 gnd 0.006876f
C1837 vdd.t178 gnd 0.125873f
C1838 vdd.t177 gnd 0.134524f
C1839 vdd.t176 gnd 0.164388f
C1840 vdd.n1208 gnd 0.210723f
C1841 vdd.n1209 gnd 0.177045f
C1842 vdd.n1211 gnd 0.010231f
C1843 vdd.n1212 gnd 0.010231f
C1844 vdd.n1213 gnd 0.008235f
C1845 vdd.n1214 gnd 0.010231f
C1846 vdd.n1216 gnd 0.010231f
C1847 vdd.n1217 gnd 0.010231f
C1848 vdd.n1218 gnd 0.010231f
C1849 vdd.n1219 gnd 0.010231f
C1850 vdd.n1220 gnd 0.008235f
C1851 vdd.n1222 gnd 0.010231f
C1852 vdd.n1223 gnd 0.010231f
C1853 vdd.n1224 gnd 0.010231f
C1854 vdd.n1225 gnd 0.010231f
C1855 vdd.n1226 gnd 0.010231f
C1856 vdd.n1227 gnd 0.008235f
C1857 vdd.n1229 gnd 0.010231f
C1858 vdd.n1230 gnd 0.010231f
C1859 vdd.n1231 gnd 0.010231f
C1860 vdd.n1232 gnd 0.010231f
C1861 vdd.n1233 gnd 0.010231f
C1862 vdd.n1234 gnd 0.008235f
C1863 vdd.n1236 gnd 0.010231f
C1864 vdd.n1237 gnd 0.010231f
C1865 vdd.n1238 gnd 0.010231f
C1866 vdd.n1239 gnd 0.010231f
C1867 vdd.n1240 gnd 0.010231f
C1868 vdd.n1241 gnd 0.008235f
C1869 vdd.n1243 gnd 0.010231f
C1870 vdd.n1244 gnd 0.010231f
C1871 vdd.n1245 gnd 0.010231f
C1872 vdd.n1246 gnd 0.010231f
C1873 vdd.n1247 gnd 0.008153f
C1874 vdd.t171 gnd 0.125873f
C1875 vdd.t170 gnd 0.134524f
C1876 vdd.t168 gnd 0.164388f
C1877 vdd.n1248 gnd 0.210723f
C1878 vdd.n1249 gnd 0.177045f
C1879 vdd.n1251 gnd 0.010231f
C1880 vdd.n1252 gnd 0.010231f
C1881 vdd.n1253 gnd 0.008235f
C1882 vdd.n1254 gnd 0.010231f
C1883 vdd.n1256 gnd 0.010231f
C1884 vdd.n1257 gnd 0.010231f
C1885 vdd.n1258 gnd 0.010231f
C1886 vdd.n1259 gnd 0.010231f
C1887 vdd.n1260 gnd 0.008235f
C1888 vdd.n1262 gnd 0.010231f
C1889 vdd.n1263 gnd 0.010231f
C1890 vdd.n1264 gnd 0.010231f
C1891 vdd.n1265 gnd 0.010231f
C1892 vdd.n1266 gnd 0.010231f
C1893 vdd.n1267 gnd 0.008235f
C1894 vdd.n1269 gnd 0.010231f
C1895 vdd.n1270 gnd 0.010231f
C1896 vdd.n1271 gnd 0.010231f
C1897 vdd.n1272 gnd 0.010231f
C1898 vdd.n1273 gnd 0.010231f
C1899 vdd.n1274 gnd 0.008235f
C1900 vdd.n1276 gnd 0.010231f
C1901 vdd.n1277 gnd 0.010231f
C1902 vdd.n1278 gnd 0.006548f
C1903 vdd.n1279 gnd 0.008235f
C1904 vdd.n1280 gnd 0.015797f
C1905 vdd.n1281 gnd 0.015797f
C1906 vdd.n1282 gnd 0.006957f
C1907 vdd.n1283 gnd 0.006957f
C1908 vdd.n1284 gnd 0.006957f
C1909 vdd.n1285 gnd 0.006957f
C1910 vdd.n1286 gnd 0.006957f
C1911 vdd.n1287 gnd 0.006957f
C1912 vdd.n1288 gnd 0.006957f
C1913 vdd.n1289 gnd 0.006957f
C1914 vdd.n1290 gnd 0.006957f
C1915 vdd.n1291 gnd 0.006957f
C1916 vdd.n1292 gnd 0.006957f
C1917 vdd.n1293 gnd 0.006957f
C1918 vdd.n1294 gnd 0.006957f
C1919 vdd.n1295 gnd 0.006957f
C1920 vdd.n1296 gnd 0.006957f
C1921 vdd.n1297 gnd 0.006957f
C1922 vdd.n1298 gnd 0.006957f
C1923 vdd.n1299 gnd 0.006957f
C1924 vdd.n1300 gnd 0.006957f
C1925 vdd.n1301 gnd 0.006957f
C1926 vdd.n1302 gnd 0.006957f
C1927 vdd.n1303 gnd 0.006957f
C1928 vdd.n1304 gnd 0.006957f
C1929 vdd.n1305 gnd 0.006957f
C1930 vdd.n1306 gnd 0.006957f
C1931 vdd.n1307 gnd 0.006957f
C1932 vdd.n1308 gnd 0.006957f
C1933 vdd.n1309 gnd 0.006957f
C1934 vdd.n1310 gnd 0.006957f
C1935 vdd.n1311 gnd 0.006957f
C1936 vdd.n1312 gnd 0.006957f
C1937 vdd.n1313 gnd 0.006957f
C1938 vdd.n1314 gnd 0.006957f
C1939 vdd.t166 gnd 0.281145f
C1940 vdd.t167 gnd 0.287787f
C1941 vdd.t164 gnd 0.183542f
C1942 vdd.n1315 gnd 0.099195f
C1943 vdd.n1316 gnd 0.056266f
C1944 vdd.n1317 gnd 0.009943f
C1945 vdd.n1318 gnd 0.006957f
C1946 vdd.t203 gnd 0.281145f
C1947 vdd.t204 gnd 0.287787f
C1948 vdd.t202 gnd 0.183542f
C1949 vdd.n1319 gnd 0.099195f
C1950 vdd.n1320 gnd 0.056266f
C1951 vdd.n1321 gnd 0.006957f
C1952 vdd.n1322 gnd 0.006957f
C1953 vdd.n1323 gnd 0.006957f
C1954 vdd.n1324 gnd 0.006957f
C1955 vdd.n1325 gnd 0.006957f
C1956 vdd.n1326 gnd 0.006957f
C1957 vdd.n1327 gnd 0.006957f
C1958 vdd.n1328 gnd 0.006957f
C1959 vdd.n1329 gnd 0.006957f
C1960 vdd.n1330 gnd 0.006957f
C1961 vdd.n1331 gnd 0.006957f
C1962 vdd.n1332 gnd 0.006957f
C1963 vdd.n1333 gnd 0.006957f
C1964 vdd.n1334 gnd 0.006957f
C1965 vdd.n1335 gnd 0.006957f
C1966 vdd.n1336 gnd 0.006957f
C1967 vdd.n1337 gnd 0.006957f
C1968 vdd.n1338 gnd 0.006957f
C1969 vdd.n1339 gnd 0.006957f
C1970 vdd.n1340 gnd 0.006957f
C1971 vdd.n1341 gnd 0.006957f
C1972 vdd.n1342 gnd 0.006957f
C1973 vdd.n1343 gnd 0.006957f
C1974 vdd.n1344 gnd 0.006957f
C1975 vdd.n1345 gnd 0.006957f
C1976 vdd.n1346 gnd 0.006957f
C1977 vdd.n1347 gnd 0.005065f
C1978 vdd.n1348 gnd 0.009943f
C1979 vdd.n1349 gnd 0.005371f
C1980 vdd.n1350 gnd 0.006957f
C1981 vdd.n1351 gnd 0.006957f
C1982 vdd.n1352 gnd 0.006957f
C1983 vdd.n1353 gnd 0.015797f
C1984 vdd.n1354 gnd 0.015797f
C1985 vdd.n1355 gnd 0.014897f
C1986 vdd.n1356 gnd 0.014897f
C1987 vdd.n1357 gnd 0.006957f
C1988 vdd.n1358 gnd 0.006957f
C1989 vdd.n1359 gnd 0.006957f
C1990 vdd.n1360 gnd 0.006957f
C1991 vdd.n1361 gnd 0.006957f
C1992 vdd.n1362 gnd 0.006957f
C1993 vdd.n1363 gnd 0.006957f
C1994 vdd.n1364 gnd 0.006957f
C1995 vdd.n1365 gnd 0.006957f
C1996 vdd.n1366 gnd 0.006957f
C1997 vdd.n1367 gnd 0.006957f
C1998 vdd.n1368 gnd 0.006957f
C1999 vdd.n1369 gnd 0.006957f
C2000 vdd.n1370 gnd 0.006957f
C2001 vdd.n1371 gnd 0.006957f
C2002 vdd.n1372 gnd 0.006957f
C2003 vdd.n1373 gnd 0.006957f
C2004 vdd.n1374 gnd 0.006957f
C2005 vdd.n1375 gnd 0.006957f
C2006 vdd.n1376 gnd 0.006957f
C2007 vdd.n1377 gnd 0.006957f
C2008 vdd.n1378 gnd 0.006957f
C2009 vdd.n1379 gnd 0.006957f
C2010 vdd.n1380 gnd 0.006957f
C2011 vdd.n1381 gnd 0.006957f
C2012 vdd.n1382 gnd 0.006957f
C2013 vdd.n1383 gnd 0.006957f
C2014 vdd.n1384 gnd 0.006957f
C2015 vdd.n1385 gnd 0.006957f
C2016 vdd.n1386 gnd 0.006957f
C2017 vdd.n1387 gnd 0.006957f
C2018 vdd.n1388 gnd 0.006957f
C2019 vdd.n1389 gnd 0.006957f
C2020 vdd.n1390 gnd 0.006957f
C2021 vdd.n1391 gnd 0.006957f
C2022 vdd.n1392 gnd 0.006957f
C2023 vdd.n1393 gnd 0.006957f
C2024 vdd.n1394 gnd 0.006957f
C2025 vdd.n1395 gnd 0.006957f
C2026 vdd.n1396 gnd 0.006957f
C2027 vdd.n1397 gnd 0.006957f
C2028 vdd.n1398 gnd 0.006957f
C2029 vdd.n1399 gnd 0.423468f
C2030 vdd.n1400 gnd 0.006957f
C2031 vdd.n1401 gnd 0.006957f
C2032 vdd.n1402 gnd 0.006957f
C2033 vdd.n1403 gnd 0.006957f
C2034 vdd.n1404 gnd 0.006957f
C2035 vdd.n1405 gnd 0.006957f
C2036 vdd.n1406 gnd 0.006957f
C2037 vdd.n1407 gnd 0.006957f
C2038 vdd.n1408 gnd 0.006957f
C2039 vdd.n1409 gnd 0.006957f
C2040 vdd.n1410 gnd 0.006957f
C2041 vdd.n1411 gnd 0.006957f
C2042 vdd.n1412 gnd 0.006957f
C2043 vdd.n1413 gnd 0.006957f
C2044 vdd.n1414 gnd 0.006957f
C2045 vdd.n1415 gnd 0.006957f
C2046 vdd.n1416 gnd 0.006957f
C2047 vdd.n1417 gnd 0.006957f
C2048 vdd.n1418 gnd 0.006957f
C2049 vdd.n1419 gnd 0.006957f
C2050 vdd.n1420 gnd 0.006957f
C2051 vdd.n1421 gnd 0.006957f
C2052 vdd.n1422 gnd 0.006957f
C2053 vdd.n1423 gnd 0.006957f
C2054 vdd.n1424 gnd 0.006957f
C2055 vdd.n1425 gnd 0.643044f
C2056 vdd.n1426 gnd 0.006957f
C2057 vdd.n1427 gnd 0.006957f
C2058 vdd.n1428 gnd 0.006957f
C2059 vdd.n1429 gnd 0.006957f
C2060 vdd.n1430 gnd 0.006957f
C2061 vdd.n1431 gnd 0.006957f
C2062 vdd.n1432 gnd 0.006957f
C2063 vdd.n1433 gnd 0.006957f
C2064 vdd.n1434 gnd 0.006957f
C2065 vdd.n1435 gnd 0.006957f
C2066 vdd.n1436 gnd 0.006957f
C2067 vdd.n1437 gnd 0.224804f
C2068 vdd.n1438 gnd 0.006957f
C2069 vdd.n1439 gnd 0.006957f
C2070 vdd.n1440 gnd 0.006957f
C2071 vdd.n1441 gnd 0.006957f
C2072 vdd.n1442 gnd 0.006957f
C2073 vdd.n1443 gnd 0.006957f
C2074 vdd.n1444 gnd 0.006957f
C2075 vdd.n1445 gnd 0.006957f
C2076 vdd.n1446 gnd 0.006957f
C2077 vdd.n1447 gnd 0.006957f
C2078 vdd.n1448 gnd 0.006957f
C2079 vdd.n1449 gnd 0.006957f
C2080 vdd.n1450 gnd 0.006957f
C2081 vdd.n1451 gnd 0.006957f
C2082 vdd.n1452 gnd 0.006957f
C2083 vdd.n1453 gnd 0.006957f
C2084 vdd.n1454 gnd 0.006957f
C2085 vdd.n1455 gnd 0.006957f
C2086 vdd.n1456 gnd 0.006957f
C2087 vdd.n1457 gnd 0.006957f
C2088 vdd.n1458 gnd 0.006957f
C2089 vdd.n1459 gnd 0.006957f
C2090 vdd.n1460 gnd 0.006957f
C2091 vdd.n1461 gnd 0.006957f
C2092 vdd.n1462 gnd 0.006957f
C2093 vdd.n1463 gnd 0.006957f
C2094 vdd.n1464 gnd 0.006957f
C2095 vdd.n1465 gnd 0.006957f
C2096 vdd.n1466 gnd 0.006957f
C2097 vdd.n1467 gnd 0.006957f
C2098 vdd.n1468 gnd 0.006957f
C2099 vdd.n1469 gnd 0.006957f
C2100 vdd.n1470 gnd 0.006957f
C2101 vdd.n1471 gnd 0.006957f
C2102 vdd.n1472 gnd 0.006957f
C2103 vdd.n1473 gnd 0.006957f
C2104 vdd.n1474 gnd 0.006957f
C2105 vdd.n1475 gnd 0.006957f
C2106 vdd.n1476 gnd 0.006957f
C2107 vdd.n1477 gnd 0.006957f
C2108 vdd.n1478 gnd 0.006957f
C2109 vdd.n1479 gnd 0.006957f
C2110 vdd.n1480 gnd 0.014897f
C2111 vdd.n1481 gnd 0.014897f
C2112 vdd.n1482 gnd 0.015797f
C2113 vdd.n1483 gnd 0.006957f
C2114 vdd.n1484 gnd 0.006957f
C2115 vdd.n1485 gnd 0.005371f
C2116 vdd.n1486 gnd 0.006957f
C2117 vdd.n1487 gnd 0.006957f
C2118 vdd.n1488 gnd 0.005065f
C2119 vdd.n1489 gnd 0.006957f
C2120 vdd.n1490 gnd 0.006957f
C2121 vdd.n1491 gnd 0.006957f
C2122 vdd.n1492 gnd 0.006957f
C2123 vdd.n1493 gnd 0.006957f
C2124 vdd.n1494 gnd 0.006957f
C2125 vdd.n1495 gnd 0.006957f
C2126 vdd.n1496 gnd 0.006957f
C2127 vdd.n1497 gnd 0.006957f
C2128 vdd.n1498 gnd 0.006957f
C2129 vdd.n1499 gnd 0.006957f
C2130 vdd.n1500 gnd 0.006957f
C2131 vdd.n1501 gnd 0.006957f
C2132 vdd.n1502 gnd 0.006957f
C2133 vdd.n1503 gnd 0.006957f
C2134 vdd.n1504 gnd 0.006957f
C2135 vdd.n1505 gnd 0.006957f
C2136 vdd.n1506 gnd 0.006957f
C2137 vdd.n1507 gnd 0.006957f
C2138 vdd.n1508 gnd 0.006957f
C2139 vdd.n1509 gnd 0.006957f
C2140 vdd.n1510 gnd 0.006957f
C2141 vdd.n1511 gnd 0.006957f
C2142 vdd.n1512 gnd 0.006957f
C2143 vdd.n1513 gnd 0.006957f
C2144 vdd.n1514 gnd 0.006957f
C2145 vdd.n1515 gnd 0.046868f
C2146 vdd.n1517 gnd 0.025281f
C2147 vdd.n1518 gnd 0.008235f
C2148 vdd.n1520 gnd 0.010231f
C2149 vdd.n1521 gnd 0.008235f
C2150 vdd.n1522 gnd 0.010231f
C2151 vdd.n1524 gnd 0.010231f
C2152 vdd.n1525 gnd 0.010231f
C2153 vdd.n1527 gnd 0.010231f
C2154 vdd.n1528 gnd 0.006835f
C2155 vdd.t169 gnd 0.5228f
C2156 vdd.n1529 gnd 0.010231f
C2157 vdd.n1530 gnd 0.025281f
C2158 vdd.n1531 gnd 0.008235f
C2159 vdd.n1532 gnd 0.010231f
C2160 vdd.n1533 gnd 0.008235f
C2161 vdd.n1534 gnd 0.010231f
C2162 vdd.n1535 gnd 1.0456f
C2163 vdd.n1536 gnd 0.010231f
C2164 vdd.n1537 gnd 0.008235f
C2165 vdd.n1538 gnd 0.008235f
C2166 vdd.n1539 gnd 0.010231f
C2167 vdd.n1540 gnd 0.008235f
C2168 vdd.n1541 gnd 0.010231f
C2169 vdd.t42 gnd 0.5228f
C2170 vdd.n1542 gnd 0.010231f
C2171 vdd.n1543 gnd 0.008235f
C2172 vdd.n1544 gnd 0.010231f
C2173 vdd.n1545 gnd 0.008235f
C2174 vdd.n1546 gnd 0.010231f
C2175 vdd.t92 gnd 0.5228f
C2176 vdd.n1547 gnd 0.010231f
C2177 vdd.n1548 gnd 0.008235f
C2178 vdd.n1549 gnd 0.010231f
C2179 vdd.n1550 gnd 0.008235f
C2180 vdd.n1551 gnd 0.010231f
C2181 vdd.n1552 gnd 0.841707f
C2182 vdd.n1553 gnd 0.867847f
C2183 vdd.t96 gnd 0.5228f
C2184 vdd.n1554 gnd 0.010231f
C2185 vdd.n1555 gnd 0.008235f
C2186 vdd.n1556 gnd 0.010231f
C2187 vdd.n1557 gnd 0.008235f
C2188 vdd.n1558 gnd 0.010231f
C2189 vdd.n1559 gnd 0.663956f
C2190 vdd.n1560 gnd 0.010231f
C2191 vdd.n1561 gnd 0.008235f
C2192 vdd.n1562 gnd 0.010231f
C2193 vdd.n1563 gnd 0.008235f
C2194 vdd.n1564 gnd 0.010231f
C2195 vdd.t39 gnd 0.5228f
C2196 vdd.t37 gnd 0.5228f
C2197 vdd.n1565 gnd 0.010231f
C2198 vdd.n1566 gnd 0.008235f
C2199 vdd.n1567 gnd 0.010231f
C2200 vdd.n1568 gnd 0.008235f
C2201 vdd.n1569 gnd 0.010231f
C2202 vdd.t4 gnd 0.5228f
C2203 vdd.n1570 gnd 0.010231f
C2204 vdd.n1571 gnd 0.008235f
C2205 vdd.n1572 gnd 0.010231f
C2206 vdd.n1573 gnd 0.008235f
C2207 vdd.n1574 gnd 0.010231f
C2208 vdd.t8 gnd 0.5228f
C2209 vdd.n1575 gnd 0.737148f
C2210 vdd.n1576 gnd 0.010231f
C2211 vdd.n1577 gnd 0.008235f
C2212 vdd.n1578 gnd 0.010231f
C2213 vdd.n1579 gnd 0.008235f
C2214 vdd.n1580 gnd 0.010231f
C2215 vdd.n1581 gnd 0.820795f
C2216 vdd.n1582 gnd 0.010231f
C2217 vdd.n1583 gnd 0.008235f
C2218 vdd.n1584 gnd 0.010231f
C2219 vdd.n1585 gnd 0.008235f
C2220 vdd.n1586 gnd 0.010231f
C2221 vdd.n1587 gnd 0.643044f
C2222 vdd.t90 gnd 0.5228f
C2223 vdd.n1588 gnd 0.010231f
C2224 vdd.n1589 gnd 0.008235f
C2225 vdd.n1590 gnd 0.010231f
C2226 vdd.n1591 gnd 0.008235f
C2227 vdd.n1592 gnd 0.010231f
C2228 vdd.t52 gnd 0.5228f
C2229 vdd.n1593 gnd 0.010231f
C2230 vdd.n1594 gnd 0.008235f
C2231 vdd.n1595 gnd 0.010231f
C2232 vdd.n1596 gnd 0.008235f
C2233 vdd.n1597 gnd 0.010231f
C2234 vdd.t110 gnd 0.5228f
C2235 vdd.n1598 gnd 0.580308f
C2236 vdd.n1599 gnd 0.010231f
C2237 vdd.n1600 gnd 0.008235f
C2238 vdd.n1601 gnd 0.010231f
C2239 vdd.n1602 gnd 0.008235f
C2240 vdd.n1603 gnd 0.010231f
C2241 vdd.t76 gnd 0.5228f
C2242 vdd.n1604 gnd 0.010231f
C2243 vdd.n1605 gnd 0.008235f
C2244 vdd.n1606 gnd 0.010231f
C2245 vdd.n1607 gnd 0.008235f
C2246 vdd.n1608 gnd 0.010231f
C2247 vdd.n1609 gnd 0.799883f
C2248 vdd.n1610 gnd 0.867847f
C2249 vdd.t44 gnd 0.5228f
C2250 vdd.n1611 gnd 0.010231f
C2251 vdd.n1612 gnd 0.008235f
C2252 vdd.n1613 gnd 0.010231f
C2253 vdd.n1614 gnd 0.008235f
C2254 vdd.n1615 gnd 0.010231f
C2255 vdd.n1616 gnd 0.622132f
C2256 vdd.n1617 gnd 0.010231f
C2257 vdd.n1618 gnd 0.008235f
C2258 vdd.n1619 gnd 0.010231f
C2259 vdd.n1620 gnd 0.008235f
C2260 vdd.n1621 gnd 0.010231f
C2261 vdd.t32 gnd 0.5228f
C2262 vdd.t128 gnd 0.5228f
C2263 vdd.n1622 gnd 0.010231f
C2264 vdd.n1623 gnd 0.008235f
C2265 vdd.n1624 gnd 0.010231f
C2266 vdd.n1625 gnd 0.008235f
C2267 vdd.n1626 gnd 0.010231f
C2268 vdd.t84 gnd 0.5228f
C2269 vdd.n1627 gnd 0.010231f
C2270 vdd.n1628 gnd 0.008235f
C2271 vdd.n1629 gnd 0.010231f
C2272 vdd.n1630 gnd 0.008235f
C2273 vdd.n1631 gnd 0.010231f
C2274 vdd.t87 gnd 0.5228f
C2275 vdd.n1632 gnd 0.778971f
C2276 vdd.n1633 gnd 0.010231f
C2277 vdd.n1634 gnd 0.008235f
C2278 vdd.n1635 gnd 0.010231f
C2279 vdd.n1636 gnd 0.008235f
C2280 vdd.n1637 gnd 0.010231f
C2281 vdd.n1638 gnd 1.0456f
C2282 vdd.n1639 gnd 0.010231f
C2283 vdd.n1640 gnd 0.008235f
C2284 vdd.n1641 gnd 0.024751f
C2285 vdd.n1642 gnd 0.006835f
C2286 vdd.n1643 gnd 0.024751f
C2287 vdd.t224 gnd 0.5228f
C2288 vdd.n1644 gnd 0.024751f
C2289 vdd.n1645 gnd 0.006835f
C2290 vdd.n1646 gnd 0.010231f
C2291 vdd.n1647 gnd 0.008235f
C2292 vdd.n1648 gnd 0.010231f
C2293 vdd.n1679 gnd 0.025281f
C2294 vdd.n1680 gnd 1.54226f
C2295 vdd.n1681 gnd 0.010231f
C2296 vdd.n1682 gnd 0.008235f
C2297 vdd.n1683 gnd 0.010231f
C2298 vdd.n1684 gnd 0.010231f
C2299 vdd.n1685 gnd 0.010231f
C2300 vdd.n1686 gnd 0.010231f
C2301 vdd.n1687 gnd 0.010231f
C2302 vdd.n1688 gnd 0.008235f
C2303 vdd.n1689 gnd 0.010231f
C2304 vdd.n1690 gnd 0.010231f
C2305 vdd.n1691 gnd 0.010231f
C2306 vdd.n1692 gnd 0.010231f
C2307 vdd.n1693 gnd 0.010231f
C2308 vdd.n1694 gnd 0.008235f
C2309 vdd.n1695 gnd 0.010231f
C2310 vdd.n1696 gnd 0.010231f
C2311 vdd.n1697 gnd 0.010231f
C2312 vdd.n1698 gnd 0.010231f
C2313 vdd.n1699 gnd 0.010231f
C2314 vdd.n1700 gnd 0.008235f
C2315 vdd.n1701 gnd 0.010231f
C2316 vdd.n1702 gnd 0.010231f
C2317 vdd.n1703 gnd 0.010231f
C2318 vdd.n1704 gnd 0.010231f
C2319 vdd.n1705 gnd 0.010231f
C2320 vdd.t234 gnd 0.125873f
C2321 vdd.t235 gnd 0.134524f
C2322 vdd.t233 gnd 0.164388f
C2323 vdd.n1706 gnd 0.210723f
C2324 vdd.n1707 gnd 0.177869f
C2325 vdd.n1708 gnd 0.017623f
C2326 vdd.n1709 gnd 0.010231f
C2327 vdd.n1710 gnd 0.010231f
C2328 vdd.n1711 gnd 0.010231f
C2329 vdd.n1712 gnd 0.010231f
C2330 vdd.n1713 gnd 0.010231f
C2331 vdd.n1714 gnd 0.008235f
C2332 vdd.n1715 gnd 0.010231f
C2333 vdd.n1716 gnd 0.010231f
C2334 vdd.n1717 gnd 0.010231f
C2335 vdd.n1718 gnd 0.010231f
C2336 vdd.n1719 gnd 0.010231f
C2337 vdd.n1720 gnd 0.008235f
C2338 vdd.n1721 gnd 0.010231f
C2339 vdd.n1722 gnd 0.010231f
C2340 vdd.n1723 gnd 0.010231f
C2341 vdd.n1724 gnd 0.010231f
C2342 vdd.n1725 gnd 0.010231f
C2343 vdd.n1726 gnd 0.008235f
C2344 vdd.n1727 gnd 0.010231f
C2345 vdd.n1728 gnd 0.010231f
C2346 vdd.n1729 gnd 0.010231f
C2347 vdd.n1730 gnd 0.010231f
C2348 vdd.n1731 gnd 0.010231f
C2349 vdd.n1732 gnd 0.008235f
C2350 vdd.n1733 gnd 0.010231f
C2351 vdd.n1734 gnd 0.010231f
C2352 vdd.n1735 gnd 0.010231f
C2353 vdd.n1736 gnd 0.010231f
C2354 vdd.n1737 gnd 0.010231f
C2355 vdd.n1738 gnd 0.008235f
C2356 vdd.n1739 gnd 0.010231f
C2357 vdd.n1740 gnd 0.010231f
C2358 vdd.n1741 gnd 0.010231f
C2359 vdd.n1742 gnd 0.010231f
C2360 vdd.n1743 gnd 0.008235f
C2361 vdd.n1744 gnd 0.010231f
C2362 vdd.n1745 gnd 0.010231f
C2363 vdd.n1746 gnd 0.010231f
C2364 vdd.n1747 gnd 0.010231f
C2365 vdd.n1748 gnd 0.010231f
C2366 vdd.n1749 gnd 0.008235f
C2367 vdd.n1750 gnd 0.010231f
C2368 vdd.n1751 gnd 0.010231f
C2369 vdd.n1752 gnd 0.010231f
C2370 vdd.n1753 gnd 0.010231f
C2371 vdd.n1754 gnd 0.010231f
C2372 vdd.n1755 gnd 0.008235f
C2373 vdd.n1756 gnd 0.010231f
C2374 vdd.n1757 gnd 0.010231f
C2375 vdd.n1758 gnd 0.010231f
C2376 vdd.n1759 gnd 0.010231f
C2377 vdd.n1760 gnd 0.010231f
C2378 vdd.n1761 gnd 0.008235f
C2379 vdd.n1762 gnd 0.010231f
C2380 vdd.n1763 gnd 0.010231f
C2381 vdd.n1764 gnd 0.010231f
C2382 vdd.n1765 gnd 0.010231f
C2383 vdd.n1766 gnd 0.010231f
C2384 vdd.n1767 gnd 0.008235f
C2385 vdd.n1768 gnd 0.010231f
C2386 vdd.n1769 gnd 0.010231f
C2387 vdd.n1770 gnd 0.010231f
C2388 vdd.n1771 gnd 0.010231f
C2389 vdd.t231 gnd 0.125873f
C2390 vdd.t232 gnd 0.134524f
C2391 vdd.t230 gnd 0.164388f
C2392 vdd.n1772 gnd 0.210723f
C2393 vdd.n1773 gnd 0.177869f
C2394 vdd.n1774 gnd 0.013505f
C2395 vdd.n1775 gnd 0.003912f
C2396 vdd.n1776 gnd 0.025281f
C2397 vdd.n1777 gnd 0.010231f
C2398 vdd.n1778 gnd 0.004323f
C2399 vdd.n1779 gnd 0.008235f
C2400 vdd.n1780 gnd 0.008235f
C2401 vdd.n1781 gnd 0.010231f
C2402 vdd.n1782 gnd 0.010231f
C2403 vdd.n1783 gnd 0.010231f
C2404 vdd.n1784 gnd 0.008235f
C2405 vdd.n1785 gnd 0.008235f
C2406 vdd.n1786 gnd 0.008235f
C2407 vdd.n1787 gnd 0.010231f
C2408 vdd.n1788 gnd 0.010231f
C2409 vdd.n1789 gnd 0.010231f
C2410 vdd.n1790 gnd 0.008235f
C2411 vdd.n1791 gnd 0.008235f
C2412 vdd.n1792 gnd 0.008235f
C2413 vdd.n1793 gnd 0.010231f
C2414 vdd.n1794 gnd 0.010231f
C2415 vdd.n1795 gnd 0.010231f
C2416 vdd.n1796 gnd 0.008235f
C2417 vdd.n1797 gnd 0.008235f
C2418 vdd.n1798 gnd 0.008235f
C2419 vdd.n1799 gnd 0.010231f
C2420 vdd.n1800 gnd 0.010231f
C2421 vdd.n1801 gnd 0.010231f
C2422 vdd.n1802 gnd 0.008235f
C2423 vdd.n1803 gnd 0.008235f
C2424 vdd.n1804 gnd 0.008235f
C2425 vdd.n1805 gnd 0.010231f
C2426 vdd.n1806 gnd 0.010231f
C2427 vdd.n1807 gnd 0.010231f
C2428 vdd.n1808 gnd 0.008153f
C2429 vdd.n1809 gnd 0.010231f
C2430 vdd.t225 gnd 0.125873f
C2431 vdd.t226 gnd 0.134524f
C2432 vdd.t223 gnd 0.164388f
C2433 vdd.n1810 gnd 0.210723f
C2434 vdd.n1811 gnd 0.177869f
C2435 vdd.n1812 gnd 0.017623f
C2436 vdd.n1813 gnd 0.0056f
C2437 vdd.n1814 gnd 0.010231f
C2438 vdd.n1815 gnd 0.010231f
C2439 vdd.n1816 gnd 0.010231f
C2440 vdd.n1817 gnd 0.008235f
C2441 vdd.n1818 gnd 0.008235f
C2442 vdd.n1819 gnd 0.008235f
C2443 vdd.n1820 gnd 0.010231f
C2444 vdd.n1821 gnd 0.010231f
C2445 vdd.n1822 gnd 0.010231f
C2446 vdd.n1823 gnd 0.008235f
C2447 vdd.n1824 gnd 0.008235f
C2448 vdd.n1825 gnd 0.008235f
C2449 vdd.n1826 gnd 0.010231f
C2450 vdd.n1827 gnd 0.010231f
C2451 vdd.n1828 gnd 0.010231f
C2452 vdd.n1829 gnd 0.008235f
C2453 vdd.n1830 gnd 0.008235f
C2454 vdd.n1831 gnd 0.008235f
C2455 vdd.n1832 gnd 0.010231f
C2456 vdd.n1833 gnd 0.010231f
C2457 vdd.n1834 gnd 0.010231f
C2458 vdd.n1835 gnd 0.008235f
C2459 vdd.n1836 gnd 0.008235f
C2460 vdd.n1837 gnd 0.008235f
C2461 vdd.n1838 gnd 0.010231f
C2462 vdd.n1839 gnd 0.010231f
C2463 vdd.n1840 gnd 0.010231f
C2464 vdd.n1841 gnd 0.008235f
C2465 vdd.n1842 gnd 0.008235f
C2466 vdd.n1843 gnd 0.006876f
C2467 vdd.n1844 gnd 0.010231f
C2468 vdd.n1845 gnd 0.010231f
C2469 vdd.n1846 gnd 0.010231f
C2470 vdd.n1847 gnd 0.006876f
C2471 vdd.n1848 gnd 0.008235f
C2472 vdd.n1849 gnd 0.008235f
C2473 vdd.n1850 gnd 0.010231f
C2474 vdd.n1851 gnd 0.010231f
C2475 vdd.n1852 gnd 0.010231f
C2476 vdd.n1853 gnd 0.008235f
C2477 vdd.n1854 gnd 0.008235f
C2478 vdd.n1855 gnd 0.008235f
C2479 vdd.n1856 gnd 0.010231f
C2480 vdd.n1857 gnd 0.010231f
C2481 vdd.n1858 gnd 0.010231f
C2482 vdd.n1859 gnd 0.008235f
C2483 vdd.n1860 gnd 0.008235f
C2484 vdd.n1861 gnd 0.008235f
C2485 vdd.n1862 gnd 0.010231f
C2486 vdd.n1863 gnd 0.010231f
C2487 vdd.n1864 gnd 0.010231f
C2488 vdd.n1865 gnd 0.008235f
C2489 vdd.n1866 gnd 0.008235f
C2490 vdd.n1867 gnd 0.008235f
C2491 vdd.n1868 gnd 0.010231f
C2492 vdd.n1869 gnd 0.010231f
C2493 vdd.n1870 gnd 0.010231f
C2494 vdd.n1871 gnd 0.008235f
C2495 vdd.n1872 gnd 0.010231f
C2496 vdd.n1873 gnd 2.47807f
C2497 vdd.n1875 gnd 0.025281f
C2498 vdd.n1876 gnd 0.006835f
C2499 vdd.n1877 gnd 0.025281f
C2500 vdd.n1878 gnd 0.024751f
C2501 vdd.n1879 gnd 0.010231f
C2502 vdd.n1880 gnd 0.008235f
C2503 vdd.n1881 gnd 0.010231f
C2504 vdd.n1882 gnd 0.528028f
C2505 vdd.n1883 gnd 0.010231f
C2506 vdd.n1884 gnd 0.008235f
C2507 vdd.n1885 gnd 0.010231f
C2508 vdd.n1886 gnd 0.010231f
C2509 vdd.n1887 gnd 0.010231f
C2510 vdd.n1888 gnd 0.008235f
C2511 vdd.n1889 gnd 0.010231f
C2512 vdd.n1890 gnd 0.956723f
C2513 vdd.n1891 gnd 1.0456f
C2514 vdd.n1892 gnd 0.010231f
C2515 vdd.n1893 gnd 0.008235f
C2516 vdd.n1894 gnd 0.010231f
C2517 vdd.n1895 gnd 0.010231f
C2518 vdd.n1896 gnd 0.010231f
C2519 vdd.n1897 gnd 0.008235f
C2520 vdd.n1898 gnd 0.010231f
C2521 vdd.n1899 gnd 0.611676f
C2522 vdd.n1900 gnd 0.010231f
C2523 vdd.n1901 gnd 0.008235f
C2524 vdd.n1902 gnd 0.010231f
C2525 vdd.n1903 gnd 0.010231f
C2526 vdd.n1904 gnd 0.010231f
C2527 vdd.n1905 gnd 0.008235f
C2528 vdd.n1906 gnd 0.010231f
C2529 vdd.n1907 gnd 0.60122f
C2530 vdd.n1908 gnd 0.789427f
C2531 vdd.n1909 gnd 0.010231f
C2532 vdd.n1910 gnd 0.008235f
C2533 vdd.n1911 gnd 0.010231f
C2534 vdd.n1912 gnd 0.010231f
C2535 vdd.n1913 gnd 0.010231f
C2536 vdd.n1914 gnd 0.008235f
C2537 vdd.n1915 gnd 0.010231f
C2538 vdd.n1916 gnd 0.867847f
C2539 vdd.n1917 gnd 0.010231f
C2540 vdd.n1918 gnd 0.008235f
C2541 vdd.n1919 gnd 0.010231f
C2542 vdd.n1920 gnd 0.010231f
C2543 vdd.n1921 gnd 0.010231f
C2544 vdd.n1922 gnd 0.008235f
C2545 vdd.n1923 gnd 0.010231f
C2546 vdd.t94 gnd 0.5228f
C2547 vdd.n1924 gnd 0.768516f
C2548 vdd.n1925 gnd 0.010231f
C2549 vdd.n1926 gnd 0.008235f
C2550 vdd.n1927 gnd 0.010231f
C2551 vdd.n1928 gnd 0.010231f
C2552 vdd.n1929 gnd 0.010231f
C2553 vdd.n1930 gnd 0.008235f
C2554 vdd.n1931 gnd 0.010231f
C2555 vdd.n1932 gnd 0.590764f
C2556 vdd.n1933 gnd 0.010231f
C2557 vdd.n1934 gnd 0.008235f
C2558 vdd.n1935 gnd 0.010231f
C2559 vdd.n1936 gnd 0.010231f
C2560 vdd.n1937 gnd 0.010231f
C2561 vdd.n1938 gnd 0.008235f
C2562 vdd.n1939 gnd 0.010231f
C2563 vdd.n1940 gnd 0.75806f
C2564 vdd.n1941 gnd 0.632588f
C2565 vdd.n1942 gnd 0.010231f
C2566 vdd.n1943 gnd 0.008235f
C2567 vdd.n1944 gnd 0.010231f
C2568 vdd.n1945 gnd 0.010231f
C2569 vdd.n1946 gnd 0.010231f
C2570 vdd.n1947 gnd 0.008235f
C2571 vdd.n1948 gnd 0.010231f
C2572 vdd.n1949 gnd 0.810339f
C2573 vdd.n1950 gnd 0.010231f
C2574 vdd.n1951 gnd 0.008235f
C2575 vdd.n1952 gnd 0.010231f
C2576 vdd.n1953 gnd 0.010231f
C2577 vdd.n1954 gnd 0.010231f
C2578 vdd.n1955 gnd 0.008235f
C2579 vdd.n1956 gnd 0.010231f
C2580 vdd.t0 gnd 0.5228f
C2581 vdd.n1957 gnd 0.867847f
C2582 vdd.n1958 gnd 0.010231f
C2583 vdd.n1959 gnd 0.008235f
C2584 vdd.n1960 gnd 0.010231f
C2585 vdd.n1961 gnd 0.007863f
C2586 vdd.n1962 gnd 0.005615f
C2587 vdd.n1963 gnd 0.005211f
C2588 vdd.n1964 gnd 0.002882f
C2589 vdd.n1965 gnd 0.006618f
C2590 vdd.n1966 gnd 0.0028f
C2591 vdd.n1967 gnd 0.002965f
C2592 vdd.n1968 gnd 0.005211f
C2593 vdd.n1969 gnd 0.0028f
C2594 vdd.n1970 gnd 0.006618f
C2595 vdd.n1971 gnd 0.002965f
C2596 vdd.n1972 gnd 0.005211f
C2597 vdd.n1973 gnd 0.0028f
C2598 vdd.n1974 gnd 0.004963f
C2599 vdd.n1975 gnd 0.004978f
C2600 vdd.t83 gnd 0.014218f
C2601 vdd.n1976 gnd 0.031635f
C2602 vdd.n1977 gnd 0.164637f
C2603 vdd.n1978 gnd 0.0028f
C2604 vdd.n1979 gnd 0.002965f
C2605 vdd.n1980 gnd 0.006618f
C2606 vdd.n1981 gnd 0.006618f
C2607 vdd.n1982 gnd 0.002965f
C2608 vdd.n1983 gnd 0.0028f
C2609 vdd.n1984 gnd 0.005211f
C2610 vdd.n1985 gnd 0.005211f
C2611 vdd.n1986 gnd 0.0028f
C2612 vdd.n1987 gnd 0.002965f
C2613 vdd.n1988 gnd 0.006618f
C2614 vdd.n1989 gnd 0.006618f
C2615 vdd.n1990 gnd 0.002965f
C2616 vdd.n1991 gnd 0.0028f
C2617 vdd.n1992 gnd 0.005211f
C2618 vdd.n1993 gnd 0.005211f
C2619 vdd.n1994 gnd 0.0028f
C2620 vdd.n1995 gnd 0.002965f
C2621 vdd.n1996 gnd 0.006618f
C2622 vdd.n1997 gnd 0.006618f
C2623 vdd.n1998 gnd 0.015646f
C2624 vdd.n1999 gnd 0.002882f
C2625 vdd.n2000 gnd 0.0028f
C2626 vdd.n2001 gnd 0.013467f
C2627 vdd.n2002 gnd 0.009402f
C2628 vdd.t135 gnd 0.03294f
C2629 vdd.t159 gnd 0.03294f
C2630 vdd.n2003 gnd 0.226387f
C2631 vdd.n2004 gnd 0.178019f
C2632 vdd.t114 gnd 0.03294f
C2633 vdd.t27 gnd 0.03294f
C2634 vdd.n2005 gnd 0.226387f
C2635 vdd.n2006 gnd 0.14366f
C2636 vdd.t98 gnd 0.03294f
C2637 vdd.t40 gnd 0.03294f
C2638 vdd.n2007 gnd 0.226387f
C2639 vdd.n2008 gnd 0.14366f
C2640 vdd.t146 gnd 0.03294f
C2641 vdd.t68 gnd 0.03294f
C2642 vdd.n2009 gnd 0.226387f
C2643 vdd.n2010 gnd 0.14366f
C2644 vdd.t120 gnd 0.03294f
C2645 vdd.t91 gnd 0.03294f
C2646 vdd.n2011 gnd 0.226387f
C2647 vdd.n2012 gnd 0.14366f
C2648 vdd.t137 gnd 0.03294f
C2649 vdd.t53 gnd 0.03294f
C2650 vdd.n2013 gnd 0.226387f
C2651 vdd.n2014 gnd 0.14366f
C2652 vdd.t156 gnd 0.03294f
C2653 vdd.t77 gnd 0.03294f
C2654 vdd.n2015 gnd 0.226387f
C2655 vdd.n2016 gnd 0.14366f
C2656 vdd.t129 gnd 0.03294f
C2657 vdd.t102 gnd 0.03294f
C2658 vdd.n2017 gnd 0.226387f
C2659 vdd.n2018 gnd 0.14366f
C2660 vdd.t147 gnd 0.03294f
C2661 vdd.t70 gnd 0.03294f
C2662 vdd.n2019 gnd 0.226387f
C2663 vdd.n2020 gnd 0.14366f
C2664 vdd.n2021 gnd 0.005615f
C2665 vdd.n2022 gnd 0.005211f
C2666 vdd.n2023 gnd 0.002882f
C2667 vdd.n2024 gnd 0.006618f
C2668 vdd.n2025 gnd 0.0028f
C2669 vdd.n2026 gnd 0.002965f
C2670 vdd.n2027 gnd 0.005211f
C2671 vdd.n2028 gnd 0.0028f
C2672 vdd.n2029 gnd 0.006618f
C2673 vdd.n2030 gnd 0.002965f
C2674 vdd.n2031 gnd 0.005211f
C2675 vdd.n2032 gnd 0.0028f
C2676 vdd.n2033 gnd 0.004963f
C2677 vdd.n2034 gnd 0.004978f
C2678 vdd.t124 gnd 0.014218f
C2679 vdd.n2035 gnd 0.031635f
C2680 vdd.n2036 gnd 0.164637f
C2681 vdd.n2037 gnd 0.0028f
C2682 vdd.n2038 gnd 0.002965f
C2683 vdd.n2039 gnd 0.006618f
C2684 vdd.n2040 gnd 0.006618f
C2685 vdd.n2041 gnd 0.002965f
C2686 vdd.n2042 gnd 0.0028f
C2687 vdd.n2043 gnd 0.005211f
C2688 vdd.n2044 gnd 0.005211f
C2689 vdd.n2045 gnd 0.0028f
C2690 vdd.n2046 gnd 0.002965f
C2691 vdd.n2047 gnd 0.006618f
C2692 vdd.n2048 gnd 0.006618f
C2693 vdd.n2049 gnd 0.002965f
C2694 vdd.n2050 gnd 0.0028f
C2695 vdd.n2051 gnd 0.005211f
C2696 vdd.n2052 gnd 0.005211f
C2697 vdd.n2053 gnd 0.0028f
C2698 vdd.n2054 gnd 0.002965f
C2699 vdd.n2055 gnd 0.006618f
C2700 vdd.n2056 gnd 0.006618f
C2701 vdd.n2057 gnd 0.015646f
C2702 vdd.n2058 gnd 0.002882f
C2703 vdd.n2059 gnd 0.0028f
C2704 vdd.n2060 gnd 0.013467f
C2705 vdd.n2061 gnd 0.009107f
C2706 vdd.n2062 gnd 0.106884f
C2707 vdd.n2063 gnd 0.005615f
C2708 vdd.n2064 gnd 0.005211f
C2709 vdd.n2065 gnd 0.002882f
C2710 vdd.n2066 gnd 0.006618f
C2711 vdd.n2067 gnd 0.0028f
C2712 vdd.n2068 gnd 0.002965f
C2713 vdd.n2069 gnd 0.005211f
C2714 vdd.n2070 gnd 0.0028f
C2715 vdd.n2071 gnd 0.006618f
C2716 vdd.n2072 gnd 0.002965f
C2717 vdd.n2073 gnd 0.005211f
C2718 vdd.n2074 gnd 0.0028f
C2719 vdd.n2075 gnd 0.004963f
C2720 vdd.n2076 gnd 0.004978f
C2721 vdd.t43 gnd 0.014218f
C2722 vdd.n2077 gnd 0.031635f
C2723 vdd.n2078 gnd 0.164637f
C2724 vdd.n2079 gnd 0.0028f
C2725 vdd.n2080 gnd 0.002965f
C2726 vdd.n2081 gnd 0.006618f
C2727 vdd.n2082 gnd 0.006618f
C2728 vdd.n2083 gnd 0.002965f
C2729 vdd.n2084 gnd 0.0028f
C2730 vdd.n2085 gnd 0.005211f
C2731 vdd.n2086 gnd 0.005211f
C2732 vdd.n2087 gnd 0.0028f
C2733 vdd.n2088 gnd 0.002965f
C2734 vdd.n2089 gnd 0.006618f
C2735 vdd.n2090 gnd 0.006618f
C2736 vdd.n2091 gnd 0.002965f
C2737 vdd.n2092 gnd 0.0028f
C2738 vdd.n2093 gnd 0.005211f
C2739 vdd.n2094 gnd 0.005211f
C2740 vdd.n2095 gnd 0.0028f
C2741 vdd.n2096 gnd 0.002965f
C2742 vdd.n2097 gnd 0.006618f
C2743 vdd.n2098 gnd 0.006618f
C2744 vdd.n2099 gnd 0.015646f
C2745 vdd.n2100 gnd 0.002882f
C2746 vdd.n2101 gnd 0.0028f
C2747 vdd.n2102 gnd 0.013467f
C2748 vdd.n2103 gnd 0.009402f
C2749 vdd.t97 gnd 0.03294f
C2750 vdd.t93 gnd 0.03294f
C2751 vdd.n2104 gnd 0.226387f
C2752 vdd.n2105 gnd 0.178019f
C2753 vdd.t38 gnd 0.03294f
C2754 vdd.t11 gnd 0.03294f
C2755 vdd.n2106 gnd 0.226387f
C2756 vdd.n2107 gnd 0.14366f
C2757 vdd.t5 gnd 0.03294f
C2758 vdd.t86 gnd 0.03294f
C2759 vdd.n2108 gnd 0.226387f
C2760 vdd.n2109 gnd 0.14366f
C2761 vdd.t61 gnd 0.03294f
C2762 vdd.t9 gnd 0.03294f
C2763 vdd.n2110 gnd 0.226387f
C2764 vdd.n2111 gnd 0.14366f
C2765 vdd.t1 gnd 0.03294f
C2766 vdd.t115 gnd 0.03294f
C2767 vdd.n2112 gnd 0.226387f
C2768 vdd.n2113 gnd 0.14366f
C2769 vdd.t111 gnd 0.03294f
C2770 vdd.t55 gnd 0.03294f
C2771 vdd.n2114 gnd 0.226387f
C2772 vdd.n2115 gnd 0.14366f
C2773 vdd.t45 gnd 0.03294f
C2774 vdd.t143 gnd 0.03294f
C2775 vdd.n2116 gnd 0.226387f
C2776 vdd.n2117 gnd 0.14366f
C2777 vdd.t138 gnd 0.03294f
C2778 vdd.t95 gnd 0.03294f
C2779 vdd.n2118 gnd 0.226387f
C2780 vdd.n2119 gnd 0.14366f
C2781 vdd.t85 gnd 0.03294f
C2782 vdd.t33 gnd 0.03294f
C2783 vdd.n2120 gnd 0.226387f
C2784 vdd.n2121 gnd 0.14366f
C2785 vdd.n2122 gnd 0.005615f
C2786 vdd.n2123 gnd 0.005211f
C2787 vdd.n2124 gnd 0.002882f
C2788 vdd.n2125 gnd 0.006618f
C2789 vdd.n2126 gnd 0.0028f
C2790 vdd.n2127 gnd 0.002965f
C2791 vdd.n2128 gnd 0.005211f
C2792 vdd.n2129 gnd 0.0028f
C2793 vdd.n2130 gnd 0.006618f
C2794 vdd.n2131 gnd 0.002965f
C2795 vdd.n2132 gnd 0.005211f
C2796 vdd.n2133 gnd 0.0028f
C2797 vdd.n2134 gnd 0.004963f
C2798 vdd.n2135 gnd 0.004978f
C2799 vdd.t88 gnd 0.014218f
C2800 vdd.n2136 gnd 0.031635f
C2801 vdd.n2137 gnd 0.164637f
C2802 vdd.n2138 gnd 0.0028f
C2803 vdd.n2139 gnd 0.002965f
C2804 vdd.n2140 gnd 0.006618f
C2805 vdd.n2141 gnd 0.006618f
C2806 vdd.n2142 gnd 0.002965f
C2807 vdd.n2143 gnd 0.0028f
C2808 vdd.n2144 gnd 0.005211f
C2809 vdd.n2145 gnd 0.005211f
C2810 vdd.n2146 gnd 0.0028f
C2811 vdd.n2147 gnd 0.002965f
C2812 vdd.n2148 gnd 0.006618f
C2813 vdd.n2149 gnd 0.006618f
C2814 vdd.n2150 gnd 0.002965f
C2815 vdd.n2151 gnd 0.0028f
C2816 vdd.n2152 gnd 0.005211f
C2817 vdd.n2153 gnd 0.005211f
C2818 vdd.n2154 gnd 0.0028f
C2819 vdd.n2155 gnd 0.002965f
C2820 vdd.n2156 gnd 0.006618f
C2821 vdd.n2157 gnd 0.006618f
C2822 vdd.n2158 gnd 0.015646f
C2823 vdd.n2159 gnd 0.002882f
C2824 vdd.n2160 gnd 0.0028f
C2825 vdd.n2161 gnd 0.013467f
C2826 vdd.n2162 gnd 0.009107f
C2827 vdd.n2163 gnd 0.063585f
C2828 vdd.n2164 gnd 0.229114f
C2829 vdd.n2165 gnd 0.005615f
C2830 vdd.n2166 gnd 0.005211f
C2831 vdd.n2167 gnd 0.002882f
C2832 vdd.n2168 gnd 0.006618f
C2833 vdd.n2169 gnd 0.0028f
C2834 vdd.n2170 gnd 0.002965f
C2835 vdd.n2171 gnd 0.005211f
C2836 vdd.n2172 gnd 0.0028f
C2837 vdd.n2173 gnd 0.006618f
C2838 vdd.n2174 gnd 0.002965f
C2839 vdd.n2175 gnd 0.005211f
C2840 vdd.n2176 gnd 0.0028f
C2841 vdd.n2177 gnd 0.004963f
C2842 vdd.n2178 gnd 0.004978f
C2843 vdd.t62 gnd 0.014218f
C2844 vdd.n2179 gnd 0.031635f
C2845 vdd.n2180 gnd 0.164637f
C2846 vdd.n2181 gnd 0.0028f
C2847 vdd.n2182 gnd 0.002965f
C2848 vdd.n2183 gnd 0.006618f
C2849 vdd.n2184 gnd 0.006618f
C2850 vdd.n2185 gnd 0.002965f
C2851 vdd.n2186 gnd 0.0028f
C2852 vdd.n2187 gnd 0.005211f
C2853 vdd.n2188 gnd 0.005211f
C2854 vdd.n2189 gnd 0.0028f
C2855 vdd.n2190 gnd 0.002965f
C2856 vdd.n2191 gnd 0.006618f
C2857 vdd.n2192 gnd 0.006618f
C2858 vdd.n2193 gnd 0.002965f
C2859 vdd.n2194 gnd 0.0028f
C2860 vdd.n2195 gnd 0.005211f
C2861 vdd.n2196 gnd 0.005211f
C2862 vdd.n2197 gnd 0.0028f
C2863 vdd.n2198 gnd 0.002965f
C2864 vdd.n2199 gnd 0.006618f
C2865 vdd.n2200 gnd 0.006618f
C2866 vdd.n2201 gnd 0.015646f
C2867 vdd.n2202 gnd 0.002882f
C2868 vdd.n2203 gnd 0.0028f
C2869 vdd.n2204 gnd 0.013467f
C2870 vdd.n2205 gnd 0.009402f
C2871 vdd.t108 gnd 0.03294f
C2872 vdd.t106 gnd 0.03294f
C2873 vdd.n2206 gnd 0.226387f
C2874 vdd.n2207 gnd 0.178019f
C2875 vdd.t59 gnd 0.03294f
C2876 vdd.t30 gnd 0.03294f
C2877 vdd.n2208 gnd 0.226387f
C2878 vdd.n2209 gnd 0.14366f
C2879 vdd.t28 gnd 0.03294f
C2880 vdd.t104 gnd 0.03294f
C2881 vdd.n2210 gnd 0.226387f
C2882 vdd.n2211 gnd 0.14366f
C2883 vdd.t78 gnd 0.03294f
C2884 vdd.t29 gnd 0.03294f
C2885 vdd.n2212 gnd 0.226387f
C2886 vdd.n2213 gnd 0.14366f
C2887 vdd.t24 gnd 0.03294f
C2888 vdd.t125 gnd 0.03294f
C2889 vdd.n2214 gnd 0.226387f
C2890 vdd.n2215 gnd 0.14366f
C2891 vdd.t123 gnd 0.03294f
C2892 vdd.t72 gnd 0.03294f
C2893 vdd.n2216 gnd 0.226387f
C2894 vdd.n2217 gnd 0.14366f
C2895 vdd.t63 gnd 0.03294f
C2896 vdd.t157 gnd 0.03294f
C2897 vdd.n2218 gnd 0.226387f
C2898 vdd.n2219 gnd 0.14366f
C2899 vdd.t151 gnd 0.03294f
C2900 vdd.t107 gnd 0.03294f
C2901 vdd.n2220 gnd 0.226387f
C2902 vdd.n2221 gnd 0.14366f
C2903 vdd.t103 gnd 0.03294f
C2904 vdd.t58 gnd 0.03294f
C2905 vdd.n2222 gnd 0.226387f
C2906 vdd.n2223 gnd 0.14366f
C2907 vdd.n2224 gnd 0.005615f
C2908 vdd.n2225 gnd 0.005211f
C2909 vdd.n2226 gnd 0.002882f
C2910 vdd.n2227 gnd 0.006618f
C2911 vdd.n2228 gnd 0.0028f
C2912 vdd.n2229 gnd 0.002965f
C2913 vdd.n2230 gnd 0.005211f
C2914 vdd.n2231 gnd 0.0028f
C2915 vdd.n2232 gnd 0.006618f
C2916 vdd.n2233 gnd 0.002965f
C2917 vdd.n2234 gnd 0.005211f
C2918 vdd.n2235 gnd 0.0028f
C2919 vdd.n2236 gnd 0.004963f
C2920 vdd.n2237 gnd 0.004978f
C2921 vdd.t105 gnd 0.014218f
C2922 vdd.n2238 gnd 0.031635f
C2923 vdd.n2239 gnd 0.164637f
C2924 vdd.n2240 gnd 0.0028f
C2925 vdd.n2241 gnd 0.002965f
C2926 vdd.n2242 gnd 0.006618f
C2927 vdd.n2243 gnd 0.006618f
C2928 vdd.n2244 gnd 0.002965f
C2929 vdd.n2245 gnd 0.0028f
C2930 vdd.n2246 gnd 0.005211f
C2931 vdd.n2247 gnd 0.005211f
C2932 vdd.n2248 gnd 0.0028f
C2933 vdd.n2249 gnd 0.002965f
C2934 vdd.n2250 gnd 0.006618f
C2935 vdd.n2251 gnd 0.006618f
C2936 vdd.n2252 gnd 0.002965f
C2937 vdd.n2253 gnd 0.0028f
C2938 vdd.n2254 gnd 0.005211f
C2939 vdd.n2255 gnd 0.005211f
C2940 vdd.n2256 gnd 0.0028f
C2941 vdd.n2257 gnd 0.002965f
C2942 vdd.n2258 gnd 0.006618f
C2943 vdd.n2259 gnd 0.006618f
C2944 vdd.n2260 gnd 0.015646f
C2945 vdd.n2261 gnd 0.002882f
C2946 vdd.n2262 gnd 0.0028f
C2947 vdd.n2263 gnd 0.013467f
C2948 vdd.n2264 gnd 0.009107f
C2949 vdd.n2265 gnd 0.063585f
C2950 vdd.n2266 gnd 0.262286f
C2951 vdd.n2267 gnd 2.99909f
C2952 vdd.n2268 gnd 0.603486f
C2953 vdd.n2269 gnd 0.007863f
C2954 vdd.n2270 gnd 0.008235f
C2955 vdd.n2271 gnd 0.010231f
C2956 vdd.n2272 gnd 0.747604f
C2957 vdd.n2273 gnd 0.010231f
C2958 vdd.n2274 gnd 0.008235f
C2959 vdd.n2275 gnd 0.010231f
C2960 vdd.n2276 gnd 0.010231f
C2961 vdd.n2277 gnd 0.010231f
C2962 vdd.n2278 gnd 0.008235f
C2963 vdd.n2279 gnd 0.010231f
C2964 vdd.n2280 gnd 0.867847f
C2965 vdd.t60 gnd 0.5228f
C2966 vdd.n2281 gnd 0.569852f
C2967 vdd.n2282 gnd 0.010231f
C2968 vdd.n2283 gnd 0.008235f
C2969 vdd.n2284 gnd 0.010231f
C2970 vdd.n2285 gnd 0.010231f
C2971 vdd.n2286 gnd 0.010231f
C2972 vdd.n2287 gnd 0.008235f
C2973 vdd.n2288 gnd 0.010231f
C2974 vdd.n2289 gnd 0.6535f
C2975 vdd.n2290 gnd 0.010231f
C2976 vdd.n2291 gnd 0.008235f
C2977 vdd.n2292 gnd 0.010231f
C2978 vdd.n2293 gnd 0.010231f
C2979 vdd.n2294 gnd 0.010231f
C2980 vdd.n2295 gnd 0.008235f
C2981 vdd.n2296 gnd 0.010231f
C2982 vdd.n2297 gnd 0.559396f
C2983 vdd.n2298 gnd 0.831251f
C2984 vdd.n2299 gnd 0.010231f
C2985 vdd.n2300 gnd 0.008235f
C2986 vdd.n2301 gnd 0.010231f
C2987 vdd.n2302 gnd 0.010231f
C2988 vdd.n2303 gnd 0.010231f
C2989 vdd.n2304 gnd 0.008235f
C2990 vdd.n2305 gnd 0.010231f
C2991 vdd.n2306 gnd 0.867847f
C2992 vdd.n2307 gnd 0.010231f
C2993 vdd.n2308 gnd 0.008235f
C2994 vdd.n2309 gnd 0.010231f
C2995 vdd.n2310 gnd 0.010231f
C2996 vdd.n2311 gnd 0.010231f
C2997 vdd.n2312 gnd 0.008235f
C2998 vdd.n2313 gnd 0.010231f
C2999 vdd.t10 gnd 0.5228f
C3000 vdd.n2314 gnd 0.726692f
C3001 vdd.n2315 gnd 0.010231f
C3002 vdd.n2316 gnd 0.008235f
C3003 vdd.n2317 gnd 0.010231f
C3004 vdd.n2318 gnd 0.010231f
C3005 vdd.n2319 gnd 0.010231f
C3006 vdd.n2320 gnd 0.008235f
C3007 vdd.n2321 gnd 0.010231f
C3008 vdd.n2322 gnd 0.54894f
C3009 vdd.n2323 gnd 0.010231f
C3010 vdd.n2324 gnd 0.008235f
C3011 vdd.n2325 gnd 0.010231f
C3012 vdd.n2326 gnd 0.010231f
C3013 vdd.n2327 gnd 0.010231f
C3014 vdd.n2328 gnd 0.008235f
C3015 vdd.n2329 gnd 0.010231f
C3016 vdd.n2330 gnd 0.716236f
C3017 vdd.n2331 gnd 0.674412f
C3018 vdd.n2332 gnd 0.010231f
C3019 vdd.n2333 gnd 0.008235f
C3020 vdd.n2334 gnd 0.010231f
C3021 vdd.n2335 gnd 0.010231f
C3022 vdd.n2336 gnd 0.010231f
C3023 vdd.n2337 gnd 0.008235f
C3024 vdd.n2338 gnd 0.010231f
C3025 vdd.n2339 gnd 0.852163f
C3026 vdd.n2340 gnd 0.010231f
C3027 vdd.n2341 gnd 0.008235f
C3028 vdd.n2342 gnd 0.010231f
C3029 vdd.n2343 gnd 0.010231f
C3030 vdd.n2344 gnd 0.024751f
C3031 vdd.n2345 gnd 0.010231f
C3032 vdd.n2346 gnd 0.010231f
C3033 vdd.n2347 gnd 0.008235f
C3034 vdd.n2348 gnd 0.010231f
C3035 vdd.n2349 gnd 0.632588f
C3036 vdd.n2350 gnd 1.0456f
C3037 vdd.n2351 gnd 0.010231f
C3038 vdd.n2352 gnd 0.008235f
C3039 vdd.n2353 gnd 0.010231f
C3040 vdd.n2354 gnd 0.010231f
C3041 vdd.n2355 gnd 0.024751f
C3042 vdd.n2356 gnd 0.006835f
C3043 vdd.n2357 gnd 0.024751f
C3044 vdd.n2358 gnd 1.4377f
C3045 vdd.n2359 gnd 0.024751f
C3046 vdd.n2360 gnd 0.025281f
C3047 vdd.n2361 gnd 0.003912f
C3048 vdd.t195 gnd 0.125873f
C3049 vdd.t194 gnd 0.134524f
C3050 vdd.t193 gnd 0.164388f
C3051 vdd.n2362 gnd 0.210723f
C3052 vdd.n2363 gnd 0.177045f
C3053 vdd.n2364 gnd 0.012682f
C3054 vdd.n2365 gnd 0.004323f
C3055 vdd.n2366 gnd 0.008799f
C3056 vdd.n2367 gnd 1.08617f
C3057 vdd.n2369 gnd 0.008235f
C3058 vdd.n2370 gnd 0.008235f
C3059 vdd.n2371 gnd 0.010231f
C3060 vdd.n2373 gnd 0.010231f
C3061 vdd.n2374 gnd 0.010231f
C3062 vdd.n2375 gnd 0.008235f
C3063 vdd.n2376 gnd 0.008235f
C3064 vdd.n2377 gnd 0.008235f
C3065 vdd.n2378 gnd 0.010231f
C3066 vdd.n2380 gnd 0.010231f
C3067 vdd.n2381 gnd 0.010231f
C3068 vdd.n2382 gnd 0.008235f
C3069 vdd.n2383 gnd 0.008235f
C3070 vdd.n2384 gnd 0.008235f
C3071 vdd.n2385 gnd 0.010231f
C3072 vdd.n2387 gnd 0.010231f
C3073 vdd.n2388 gnd 0.010231f
C3074 vdd.n2389 gnd 0.008235f
C3075 vdd.n2390 gnd 0.008235f
C3076 vdd.n2391 gnd 0.008235f
C3077 vdd.n2392 gnd 0.010231f
C3078 vdd.n2394 gnd 0.010231f
C3079 vdd.n2395 gnd 0.010231f
C3080 vdd.n2396 gnd 0.008235f
C3081 vdd.n2397 gnd 0.010231f
C3082 vdd.n2398 gnd 0.010231f
C3083 vdd.n2399 gnd 0.010231f
C3084 vdd.n2400 gnd 0.016799f
C3085 vdd.n2401 gnd 0.0056f
C3086 vdd.n2402 gnd 0.008235f
C3087 vdd.n2403 gnd 0.010231f
C3088 vdd.n2405 gnd 0.010231f
C3089 vdd.n2406 gnd 0.010231f
C3090 vdd.n2407 gnd 0.008235f
C3091 vdd.n2408 gnd 0.008235f
C3092 vdd.n2409 gnd 0.008235f
C3093 vdd.n2410 gnd 0.010231f
C3094 vdd.n2412 gnd 0.010231f
C3095 vdd.n2413 gnd 0.010231f
C3096 vdd.n2414 gnd 0.008235f
C3097 vdd.n2415 gnd 0.008235f
C3098 vdd.n2416 gnd 0.008235f
C3099 vdd.n2417 gnd 0.010231f
C3100 vdd.n2419 gnd 0.010231f
C3101 vdd.n2420 gnd 0.010231f
C3102 vdd.n2421 gnd 0.008235f
C3103 vdd.n2422 gnd 0.008235f
C3104 vdd.n2423 gnd 0.008235f
C3105 vdd.n2424 gnd 0.010231f
C3106 vdd.n2426 gnd 0.010231f
C3107 vdd.n2427 gnd 0.010231f
C3108 vdd.n2428 gnd 0.008235f
C3109 vdd.n2429 gnd 0.008235f
C3110 vdd.n2430 gnd 0.008235f
C3111 vdd.n2431 gnd 0.010231f
C3112 vdd.n2433 gnd 0.010231f
C3113 vdd.n2434 gnd 0.010231f
C3114 vdd.n2435 gnd 0.008235f
C3115 vdd.n2436 gnd 0.010231f
C3116 vdd.n2437 gnd 0.010231f
C3117 vdd.n2438 gnd 0.010231f
C3118 vdd.n2439 gnd 0.016799f
C3119 vdd.n2440 gnd 0.006876f
C3120 vdd.n2441 gnd 0.008235f
C3121 vdd.n2442 gnd 0.010231f
C3122 vdd.n2444 gnd 0.010231f
C3123 vdd.n2445 gnd 0.010231f
C3124 vdd.n2446 gnd 0.008235f
C3125 vdd.n2447 gnd 0.008235f
C3126 vdd.n2448 gnd 0.008235f
C3127 vdd.n2449 gnd 0.010231f
C3128 vdd.n2451 gnd 0.010231f
C3129 vdd.n2452 gnd 0.010231f
C3130 vdd.n2453 gnd 0.008235f
C3131 vdd.n2454 gnd 0.008235f
C3132 vdd.n2455 gnd 0.008235f
C3133 vdd.n2456 gnd 0.010231f
C3134 vdd.n2458 gnd 0.010231f
C3135 vdd.n2459 gnd 0.010231f
C3136 vdd.n2460 gnd 0.008235f
C3137 vdd.n2461 gnd 0.008235f
C3138 vdd.n2462 gnd 0.008235f
C3139 vdd.n2463 gnd 0.010231f
C3140 vdd.n2465 gnd 0.010231f
C3141 vdd.n2466 gnd 0.008235f
C3142 vdd.n2467 gnd 0.008235f
C3143 vdd.n2468 gnd 0.010231f
C3144 vdd.n2470 gnd 0.010231f
C3145 vdd.n2471 gnd 0.010231f
C3146 vdd.n2472 gnd 0.008235f
C3147 vdd.n2473 gnd 0.008799f
C3148 vdd.n2474 gnd 1.08617f
C3149 vdd.n2475 gnd 0.046868f
C3150 vdd.n2476 gnd 0.006957f
C3151 vdd.n2477 gnd 0.006957f
C3152 vdd.n2478 gnd 0.006957f
C3153 vdd.n2479 gnd 0.006957f
C3154 vdd.n2480 gnd 0.006957f
C3155 vdd.n2481 gnd 0.006957f
C3156 vdd.n2482 gnd 0.006957f
C3157 vdd.n2483 gnd 0.006957f
C3158 vdd.n2484 gnd 0.006957f
C3159 vdd.n2485 gnd 0.006957f
C3160 vdd.n2486 gnd 0.006957f
C3161 vdd.n2487 gnd 0.006957f
C3162 vdd.n2488 gnd 0.006957f
C3163 vdd.n2489 gnd 0.006957f
C3164 vdd.n2490 gnd 0.006957f
C3165 vdd.n2491 gnd 0.006957f
C3166 vdd.n2492 gnd 0.006957f
C3167 vdd.n2493 gnd 0.006957f
C3168 vdd.n2494 gnd 0.006957f
C3169 vdd.n2495 gnd 0.006957f
C3170 vdd.n2496 gnd 0.006957f
C3171 vdd.n2497 gnd 0.006957f
C3172 vdd.n2498 gnd 0.006957f
C3173 vdd.n2499 gnd 0.006957f
C3174 vdd.n2500 gnd 0.006957f
C3175 vdd.n2501 gnd 0.006957f
C3176 vdd.n2502 gnd 0.006957f
C3177 vdd.n2503 gnd 0.006957f
C3178 vdd.n2504 gnd 0.006957f
C3179 vdd.n2505 gnd 0.006957f
C3180 vdd.n2506 gnd 12.3485f
C3181 vdd.n2508 gnd 0.015797f
C3182 vdd.n2509 gnd 0.015797f
C3183 vdd.n2510 gnd 0.014897f
C3184 vdd.n2511 gnd 0.006957f
C3185 vdd.n2512 gnd 0.006957f
C3186 vdd.n2513 gnd 0.711008f
C3187 vdd.n2514 gnd 0.006957f
C3188 vdd.n2515 gnd 0.006957f
C3189 vdd.n2516 gnd 0.006957f
C3190 vdd.n2517 gnd 0.006957f
C3191 vdd.n2518 gnd 0.006957f
C3192 vdd.n2519 gnd 0.559396f
C3193 vdd.n2520 gnd 0.006957f
C3194 vdd.n2521 gnd 0.006957f
C3195 vdd.n2522 gnd 0.006957f
C3196 vdd.n2523 gnd 0.006957f
C3197 vdd.n2524 gnd 0.006957f
C3198 vdd.n2525 gnd 0.711008f
C3199 vdd.n2526 gnd 0.006957f
C3200 vdd.n2527 gnd 0.006957f
C3201 vdd.n2528 gnd 0.006957f
C3202 vdd.n2529 gnd 0.006957f
C3203 vdd.n2530 gnd 0.006957f
C3204 vdd.n2531 gnd 0.711008f
C3205 vdd.n2532 gnd 0.006957f
C3206 vdd.n2533 gnd 0.006957f
C3207 vdd.n2534 gnd 0.006957f
C3208 vdd.n2535 gnd 0.006957f
C3209 vdd.n2536 gnd 0.006957f
C3210 vdd.n2537 gnd 0.684868f
C3211 vdd.n2538 gnd 0.006957f
C3212 vdd.n2539 gnd 0.006957f
C3213 vdd.n2540 gnd 0.006957f
C3214 vdd.n2541 gnd 0.006957f
C3215 vdd.n2542 gnd 0.006957f
C3216 vdd.n2543 gnd 0.528028f
C3217 vdd.n2544 gnd 0.006957f
C3218 vdd.n2545 gnd 0.006957f
C3219 vdd.n2546 gnd 0.006957f
C3220 vdd.n2547 gnd 0.006957f
C3221 vdd.n2548 gnd 0.006957f
C3222 vdd.n2549 gnd 0.371188f
C3223 vdd.n2550 gnd 0.006957f
C3224 vdd.n2551 gnd 0.006957f
C3225 vdd.n2552 gnd 0.006957f
C3226 vdd.n2553 gnd 0.006957f
C3227 vdd.n2554 gnd 0.006957f
C3228 vdd.n2555 gnd 0.49666f
C3229 vdd.n2556 gnd 0.006957f
C3230 vdd.n2557 gnd 0.006957f
C3231 vdd.n2558 gnd 0.006957f
C3232 vdd.n2559 gnd 0.006957f
C3233 vdd.n2560 gnd 0.006957f
C3234 vdd.n2561 gnd 0.6535f
C3235 vdd.n2562 gnd 0.006957f
C3236 vdd.n2563 gnd 0.006957f
C3237 vdd.n2564 gnd 0.006957f
C3238 vdd.n2565 gnd 0.006957f
C3239 vdd.n2566 gnd 0.006957f
C3240 vdd.n2567 gnd 0.711008f
C3241 vdd.n2568 gnd 0.006957f
C3242 vdd.n2569 gnd 0.006957f
C3243 vdd.n2570 gnd 0.006957f
C3244 vdd.n2571 gnd 0.006957f
C3245 vdd.n2572 gnd 0.006957f
C3246 vdd.n2573 gnd 0.611676f
C3247 vdd.n2574 gnd 0.006957f
C3248 vdd.n2575 gnd 0.006957f
C3249 vdd.n2576 gnd 0.005525f
C3250 vdd.n2577 gnd 0.020155f
C3251 vdd.n2578 gnd 0.004911f
C3252 vdd.n2579 gnd 0.006957f
C3253 vdd.n2580 gnd 0.454836f
C3254 vdd.n2581 gnd 0.006957f
C3255 vdd.n2582 gnd 0.006957f
C3256 vdd.n2583 gnd 0.006957f
C3257 vdd.n2584 gnd 0.006957f
C3258 vdd.n2585 gnd 0.006957f
C3259 vdd.n2586 gnd 0.413012f
C3260 vdd.n2587 gnd 0.006957f
C3261 vdd.n2588 gnd 0.006957f
C3262 vdd.n2589 gnd 0.006957f
C3263 vdd.n2590 gnd 0.006957f
C3264 vdd.n2591 gnd 0.006957f
C3265 vdd.n2592 gnd 0.569852f
C3266 vdd.n2593 gnd 0.006957f
C3267 vdd.n2594 gnd 0.006957f
C3268 vdd.n2595 gnd 0.006957f
C3269 vdd.n2596 gnd 0.006957f
C3270 vdd.n2597 gnd 0.006957f
C3271 vdd.n2598 gnd 0.62736f
C3272 vdd.n2599 gnd 0.006957f
C3273 vdd.n2600 gnd 0.006957f
C3274 vdd.n2601 gnd 0.006957f
C3275 vdd.n2602 gnd 0.006957f
C3276 vdd.n2603 gnd 0.006957f
C3277 vdd.n2604 gnd 0.47052f
C3278 vdd.n2605 gnd 0.006957f
C3279 vdd.n2606 gnd 0.006957f
C3280 vdd.n2607 gnd 0.006957f
C3281 vdd.n2608 gnd 0.006957f
C3282 vdd.n2609 gnd 0.006957f
C3283 vdd.n2610 gnd 0.224804f
C3284 vdd.n2611 gnd 0.006957f
C3285 vdd.n2612 gnd 0.006957f
C3286 vdd.n2613 gnd 0.006957f
C3287 vdd.n2614 gnd 0.006957f
C3288 vdd.n2615 gnd 0.006957f
C3289 vdd.n2616 gnd 0.224804f
C3290 vdd.n2617 gnd 0.006957f
C3291 vdd.n2618 gnd 0.006957f
C3292 vdd.n2619 gnd 0.006957f
C3293 vdd.n2620 gnd 0.006957f
C3294 vdd.n2621 gnd 0.006957f
C3295 vdd.n2622 gnd 0.711008f
C3296 vdd.n2623 gnd 0.006957f
C3297 vdd.n2624 gnd 0.006957f
C3298 vdd.n2625 gnd 0.006957f
C3299 vdd.n2626 gnd 0.006957f
C3300 vdd.n2627 gnd 0.006957f
C3301 vdd.n2628 gnd 0.006957f
C3302 vdd.n2629 gnd 0.006957f
C3303 vdd.n2630 gnd 0.491432f
C3304 vdd.n2631 gnd 0.006957f
C3305 vdd.n2632 gnd 0.006957f
C3306 vdd.n2633 gnd 0.006957f
C3307 vdd.n2634 gnd 0.006957f
C3308 vdd.n2635 gnd 0.006957f
C3309 vdd.n2636 gnd 0.006957f
C3310 vdd.n2637 gnd 0.44438f
C3311 vdd.n2638 gnd 0.006957f
C3312 vdd.n2639 gnd 0.006957f
C3313 vdd.n2640 gnd 0.006957f
C3314 vdd.n2641 gnd 0.015797f
C3315 vdd.n2642 gnd 0.014897f
C3316 vdd.n2643 gnd 0.006957f
C3317 vdd.n2644 gnd 0.006957f
C3318 vdd.n2645 gnd 0.005371f
C3319 vdd.n2646 gnd 0.006957f
C3320 vdd.n2647 gnd 0.006957f
C3321 vdd.n2648 gnd 0.005065f
C3322 vdd.n2649 gnd 0.006957f
C3323 vdd.n2650 gnd 0.006957f
C3324 vdd.n2651 gnd 0.006957f
C3325 vdd.n2652 gnd 0.006957f
C3326 vdd.n2653 gnd 0.006957f
C3327 vdd.n2654 gnd 0.006957f
C3328 vdd.n2655 gnd 0.006957f
C3329 vdd.n2656 gnd 0.006957f
C3330 vdd.n2657 gnd 0.006957f
C3331 vdd.n2658 gnd 0.006957f
C3332 vdd.n2659 gnd 0.006957f
C3333 vdd.n2660 gnd 0.006957f
C3334 vdd.n2661 gnd 0.006957f
C3335 vdd.n2662 gnd 0.006957f
C3336 vdd.n2663 gnd 0.006957f
C3337 vdd.n2664 gnd 0.006957f
C3338 vdd.n2665 gnd 0.006957f
C3339 vdd.n2666 gnd 0.006957f
C3340 vdd.n2667 gnd 0.006957f
C3341 vdd.n2668 gnd 0.006957f
C3342 vdd.n2669 gnd 0.006957f
C3343 vdd.n2670 gnd 0.006957f
C3344 vdd.n2671 gnd 0.006957f
C3345 vdd.n2672 gnd 0.006957f
C3346 vdd.n2673 gnd 0.006957f
C3347 vdd.n2674 gnd 0.006957f
C3348 vdd.n2675 gnd 0.006957f
C3349 vdd.n2676 gnd 0.006957f
C3350 vdd.n2677 gnd 0.006957f
C3351 vdd.n2678 gnd 0.006957f
C3352 vdd.n2679 gnd 0.006957f
C3353 vdd.n2680 gnd 0.006957f
C3354 vdd.n2681 gnd 0.006957f
C3355 vdd.n2682 gnd 0.006957f
C3356 vdd.n2683 gnd 0.006957f
C3357 vdd.n2684 gnd 0.006957f
C3358 vdd.n2685 gnd 0.006957f
C3359 vdd.n2686 gnd 0.006957f
C3360 vdd.n2687 gnd 0.006957f
C3361 vdd.n2688 gnd 0.006957f
C3362 vdd.n2689 gnd 0.006957f
C3363 vdd.n2690 gnd 0.006957f
C3364 vdd.n2691 gnd 0.006957f
C3365 vdd.n2692 gnd 0.006957f
C3366 vdd.n2693 gnd 0.006957f
C3367 vdd.n2694 gnd 0.006957f
C3368 vdd.n2695 gnd 0.006957f
C3369 vdd.n2696 gnd 0.006957f
C3370 vdd.n2697 gnd 0.006957f
C3371 vdd.n2698 gnd 0.006957f
C3372 vdd.n2699 gnd 0.006957f
C3373 vdd.n2700 gnd 0.006957f
C3374 vdd.n2701 gnd 0.006957f
C3375 vdd.n2702 gnd 0.006957f
C3376 vdd.n2703 gnd 0.006957f
C3377 vdd.n2704 gnd 0.006957f
C3378 vdd.n2705 gnd 0.006957f
C3379 vdd.n2706 gnd 0.006957f
C3380 vdd.n2707 gnd 0.006957f
C3381 vdd.n2708 gnd 0.006957f
C3382 vdd.n2709 gnd 0.015797f
C3383 vdd.n2710 gnd 0.014897f
C3384 vdd.n2711 gnd 0.014897f
C3385 vdd.n2712 gnd 0.805111f
C3386 vdd.n2713 gnd 0.014897f
C3387 vdd.n2714 gnd 0.015797f
C3388 vdd.n2715 gnd 0.014897f
C3389 vdd.n2716 gnd 0.006957f
C3390 vdd.n2717 gnd 0.006957f
C3391 vdd.n2718 gnd 0.006957f
C3392 vdd.n2719 gnd 0.005371f
C3393 vdd.n2720 gnd 0.009943f
C3394 vdd.n2721 gnd 0.005065f
C3395 vdd.n2722 gnd 0.006957f
C3396 vdd.n2723 gnd 0.006957f
C3397 vdd.n2724 gnd 0.006957f
C3398 vdd.n2725 gnd 0.006957f
C3399 vdd.n2726 gnd 0.006957f
C3400 vdd.n2727 gnd 0.006957f
C3401 vdd.n2728 gnd 0.006957f
C3402 vdd.n2729 gnd 0.006957f
C3403 vdd.n2730 gnd 0.006957f
C3404 vdd.n2731 gnd 0.006957f
C3405 vdd.n2732 gnd 0.006957f
C3406 vdd.n2733 gnd 0.006957f
C3407 vdd.n2734 gnd 0.006957f
C3408 vdd.n2735 gnd 0.006957f
C3409 vdd.n2736 gnd 0.006957f
C3410 vdd.n2737 gnd 0.006957f
C3411 vdd.n2738 gnd 0.006957f
C3412 vdd.n2739 gnd 0.006957f
C3413 vdd.n2740 gnd 0.006957f
C3414 vdd.n2741 gnd 0.006957f
C3415 vdd.n2742 gnd 0.006957f
C3416 vdd.n2743 gnd 0.006957f
C3417 vdd.n2744 gnd 0.006957f
C3418 vdd.n2745 gnd 0.006957f
C3419 vdd.n2746 gnd 0.006957f
C3420 vdd.n2747 gnd 0.006957f
C3421 vdd.n2748 gnd 0.006957f
C3422 vdd.n2749 gnd 0.006957f
C3423 vdd.n2750 gnd 0.006957f
C3424 vdd.n2751 gnd 0.006957f
C3425 vdd.n2752 gnd 0.006957f
C3426 vdd.n2753 gnd 0.006957f
C3427 vdd.n2754 gnd 0.006957f
C3428 vdd.n2755 gnd 0.006957f
C3429 vdd.n2756 gnd 0.006957f
C3430 vdd.n2757 gnd 0.006957f
C3431 vdd.n2758 gnd 0.006957f
C3432 vdd.n2759 gnd 0.006957f
C3433 vdd.n2760 gnd 0.006957f
C3434 vdd.n2761 gnd 0.006957f
C3435 vdd.n2762 gnd 0.006957f
C3436 vdd.n2763 gnd 0.006957f
C3437 vdd.n2764 gnd 0.006957f
C3438 vdd.n2765 gnd 0.006957f
C3439 vdd.n2766 gnd 0.006957f
C3440 vdd.n2767 gnd 0.006957f
C3441 vdd.n2768 gnd 0.006957f
C3442 vdd.n2769 gnd 0.006957f
C3443 vdd.n2770 gnd 0.006957f
C3444 vdd.n2771 gnd 0.006957f
C3445 vdd.n2772 gnd 0.006957f
C3446 vdd.n2773 gnd 0.006957f
C3447 vdd.n2774 gnd 0.006957f
C3448 vdd.n2775 gnd 0.006957f
C3449 vdd.n2776 gnd 0.006957f
C3450 vdd.n2777 gnd 0.006957f
C3451 vdd.n2778 gnd 0.006957f
C3452 vdd.n2779 gnd 0.006957f
C3453 vdd.n2780 gnd 0.006957f
C3454 vdd.n2781 gnd 0.006957f
C3455 vdd.n2782 gnd 0.015797f
C3456 vdd.n2783 gnd 0.015797f
C3457 vdd.n2784 gnd 0.867847f
C3458 vdd.t264 gnd 3.08452f
C3459 vdd.t251 gnd 3.08452f
C3460 vdd.n2818 gnd 0.015797f
C3461 vdd.t269 gnd 0.606448f
C3462 vdd.n2819 gnd 0.006957f
C3463 vdd.t214 gnd 0.281145f
C3464 vdd.t215 gnd 0.287787f
C3465 vdd.t212 gnd 0.183542f
C3466 vdd.n2820 gnd 0.099195f
C3467 vdd.n2821 gnd 0.056266f
C3468 vdd.n2822 gnd 0.006957f
C3469 vdd.t221 gnd 0.281145f
C3470 vdd.t222 gnd 0.287787f
C3471 vdd.t220 gnd 0.183542f
C3472 vdd.n2823 gnd 0.099195f
C3473 vdd.n2824 gnd 0.056266f
C3474 vdd.n2825 gnd 0.009943f
C3475 vdd.n2826 gnd 0.015797f
C3476 vdd.n2827 gnd 0.015797f
C3477 vdd.n2828 gnd 0.006957f
C3478 vdd.n2829 gnd 0.006957f
C3479 vdd.n2830 gnd 0.006957f
C3480 vdd.n2831 gnd 0.006957f
C3481 vdd.n2832 gnd 0.006957f
C3482 vdd.n2833 gnd 0.006957f
C3483 vdd.n2834 gnd 0.006957f
C3484 vdd.n2835 gnd 0.006957f
C3485 vdd.n2836 gnd 0.006957f
C3486 vdd.n2837 gnd 0.006957f
C3487 vdd.n2838 gnd 0.006957f
C3488 vdd.n2839 gnd 0.006957f
C3489 vdd.n2840 gnd 0.006957f
C3490 vdd.n2841 gnd 0.006957f
C3491 vdd.n2842 gnd 0.006957f
C3492 vdd.n2843 gnd 0.006957f
C3493 vdd.n2844 gnd 0.006957f
C3494 vdd.n2845 gnd 0.006957f
C3495 vdd.n2846 gnd 0.006957f
C3496 vdd.n2847 gnd 0.006957f
C3497 vdd.n2848 gnd 0.006957f
C3498 vdd.n2849 gnd 0.006957f
C3499 vdd.n2850 gnd 0.006957f
C3500 vdd.n2851 gnd 0.006957f
C3501 vdd.n2852 gnd 0.006957f
C3502 vdd.n2853 gnd 0.006957f
C3503 vdd.n2854 gnd 0.006957f
C3504 vdd.n2855 gnd 0.006957f
C3505 vdd.n2856 gnd 0.006957f
C3506 vdd.n2857 gnd 0.006957f
C3507 vdd.n2858 gnd 0.006957f
C3508 vdd.n2859 gnd 0.006957f
C3509 vdd.n2860 gnd 0.006957f
C3510 vdd.n2861 gnd 0.006957f
C3511 vdd.n2862 gnd 0.006957f
C3512 vdd.n2863 gnd 0.006957f
C3513 vdd.n2864 gnd 0.006957f
C3514 vdd.n2865 gnd 0.006957f
C3515 vdd.n2866 gnd 0.006957f
C3516 vdd.n2867 gnd 0.006957f
C3517 vdd.n2868 gnd 0.006957f
C3518 vdd.n2869 gnd 0.006957f
C3519 vdd.n2870 gnd 0.006957f
C3520 vdd.n2871 gnd 0.006957f
C3521 vdd.n2872 gnd 0.006957f
C3522 vdd.n2873 gnd 0.006957f
C3523 vdd.n2874 gnd 0.006957f
C3524 vdd.n2875 gnd 0.006957f
C3525 vdd.n2876 gnd 0.006957f
C3526 vdd.n2877 gnd 0.006957f
C3527 vdd.n2878 gnd 0.006957f
C3528 vdd.n2879 gnd 0.006957f
C3529 vdd.n2880 gnd 0.006957f
C3530 vdd.n2881 gnd 0.006957f
C3531 vdd.n2882 gnd 0.006957f
C3532 vdd.n2883 gnd 0.006957f
C3533 vdd.n2884 gnd 0.006957f
C3534 vdd.n2885 gnd 0.006957f
C3535 vdd.n2886 gnd 0.006957f
C3536 vdd.n2887 gnd 0.006957f
C3537 vdd.n2888 gnd 0.005065f
C3538 vdd.n2889 gnd 0.006957f
C3539 vdd.n2890 gnd 0.006957f
C3540 vdd.n2891 gnd 0.005371f
C3541 vdd.n2892 gnd 0.006957f
C3542 vdd.n2893 gnd 0.006957f
C3543 vdd.n2894 gnd 0.015797f
C3544 vdd.n2895 gnd 0.014897f
C3545 vdd.n2896 gnd 0.014897f
C3546 vdd.n2897 gnd 0.006957f
C3547 vdd.n2898 gnd 0.006957f
C3548 vdd.n2899 gnd 0.006957f
C3549 vdd.n2900 gnd 0.006957f
C3550 vdd.n2901 gnd 0.006957f
C3551 vdd.n2902 gnd 0.006957f
C3552 vdd.n2903 gnd 0.006957f
C3553 vdd.n2904 gnd 0.006957f
C3554 vdd.n2905 gnd 0.006957f
C3555 vdd.n2906 gnd 0.006957f
C3556 vdd.n2907 gnd 0.006957f
C3557 vdd.n2908 gnd 0.006957f
C3558 vdd.n2909 gnd 0.006957f
C3559 vdd.n2910 gnd 0.006957f
C3560 vdd.n2911 gnd 0.006957f
C3561 vdd.n2912 gnd 0.006957f
C3562 vdd.n2913 gnd 0.006957f
C3563 vdd.n2914 gnd 0.006957f
C3564 vdd.n2915 gnd 0.006957f
C3565 vdd.n2916 gnd 0.006957f
C3566 vdd.n2917 gnd 0.006957f
C3567 vdd.n2918 gnd 0.006957f
C3568 vdd.n2919 gnd 0.006957f
C3569 vdd.n2920 gnd 0.006957f
C3570 vdd.n2921 gnd 0.006957f
C3571 vdd.n2922 gnd 0.006957f
C3572 vdd.n2923 gnd 0.006957f
C3573 vdd.n2924 gnd 0.006957f
C3574 vdd.n2925 gnd 0.006957f
C3575 vdd.n2926 gnd 0.006957f
C3576 vdd.n2927 gnd 0.006957f
C3577 vdd.n2928 gnd 0.006957f
C3578 vdd.n2929 gnd 0.006957f
C3579 vdd.n2930 gnd 0.006957f
C3580 vdd.n2931 gnd 0.006957f
C3581 vdd.n2932 gnd 0.006957f
C3582 vdd.n2933 gnd 0.006957f
C3583 vdd.n2934 gnd 0.006957f
C3584 vdd.n2935 gnd 0.006957f
C3585 vdd.n2936 gnd 0.006957f
C3586 vdd.n2937 gnd 0.006957f
C3587 vdd.n2938 gnd 0.006957f
C3588 vdd.n2939 gnd 0.006957f
C3589 vdd.n2940 gnd 0.006957f
C3590 vdd.n2941 gnd 0.006957f
C3591 vdd.n2942 gnd 0.006957f
C3592 vdd.n2943 gnd 0.006957f
C3593 vdd.n2944 gnd 0.006957f
C3594 vdd.n2945 gnd 0.006957f
C3595 vdd.n2946 gnd 0.006957f
C3596 vdd.n2947 gnd 0.006957f
C3597 vdd.n2948 gnd 0.006957f
C3598 vdd.n2949 gnd 0.006957f
C3599 vdd.n2950 gnd 0.006957f
C3600 vdd.n2951 gnd 0.006957f
C3601 vdd.n2952 gnd 0.006957f
C3602 vdd.n2953 gnd 0.006957f
C3603 vdd.n2954 gnd 0.006957f
C3604 vdd.n2955 gnd 0.006957f
C3605 vdd.n2956 gnd 0.006957f
C3606 vdd.n2957 gnd 0.006957f
C3607 vdd.n2958 gnd 0.006957f
C3608 vdd.n2959 gnd 0.006957f
C3609 vdd.n2960 gnd 0.006957f
C3610 vdd.n2961 gnd 0.006957f
C3611 vdd.n2962 gnd 0.006957f
C3612 vdd.n2963 gnd 0.006957f
C3613 vdd.n2964 gnd 0.006957f
C3614 vdd.n2965 gnd 0.006957f
C3615 vdd.n2966 gnd 0.006957f
C3616 vdd.n2967 gnd 0.006957f
C3617 vdd.n2968 gnd 0.006957f
C3618 vdd.n2969 gnd 0.006957f
C3619 vdd.n2970 gnd 0.006957f
C3620 vdd.n2971 gnd 0.006957f
C3621 vdd.n2972 gnd 0.006957f
C3622 vdd.n2973 gnd 0.006957f
C3623 vdd.n2974 gnd 0.006957f
C3624 vdd.n2975 gnd 0.006957f
C3625 vdd.n2976 gnd 0.006957f
C3626 vdd.n2977 gnd 0.006957f
C3627 vdd.n2978 gnd 0.006957f
C3628 vdd.n2979 gnd 0.006957f
C3629 vdd.n2980 gnd 0.006957f
C3630 vdd.n2981 gnd 0.006957f
C3631 vdd.n2982 gnd 0.006957f
C3632 vdd.n2983 gnd 0.006957f
C3633 vdd.n2984 gnd 0.006957f
C3634 vdd.n2985 gnd 0.006957f
C3635 vdd.n2986 gnd 0.006957f
C3636 vdd.n2987 gnd 0.006957f
C3637 vdd.n2988 gnd 0.006957f
C3638 vdd.n2989 gnd 0.006957f
C3639 vdd.n2990 gnd 0.006957f
C3640 vdd.n2991 gnd 0.006957f
C3641 vdd.n2992 gnd 0.006957f
C3642 vdd.n2993 gnd 0.006957f
C3643 vdd.n2994 gnd 0.006957f
C3644 vdd.n2995 gnd 0.006957f
C3645 vdd.n2996 gnd 0.006957f
C3646 vdd.n2997 gnd 0.006957f
C3647 vdd.n2998 gnd 0.224804f
C3648 vdd.n2999 gnd 0.006957f
C3649 vdd.n3000 gnd 0.006957f
C3650 vdd.n3001 gnd 0.006957f
C3651 vdd.n3002 gnd 0.006957f
C3652 vdd.n3003 gnd 0.006957f
C3653 vdd.n3004 gnd 0.224804f
C3654 vdd.n3005 gnd 0.006957f
C3655 vdd.n3006 gnd 0.006957f
C3656 vdd.n3007 gnd 0.006957f
C3657 vdd.n3008 gnd 0.006957f
C3658 vdd.n3009 gnd 0.006957f
C3659 vdd.n3010 gnd 0.006957f
C3660 vdd.n3011 gnd 0.006957f
C3661 vdd.n3012 gnd 0.006957f
C3662 vdd.n3013 gnd 0.006957f
C3663 vdd.n3014 gnd 0.006957f
C3664 vdd.n3015 gnd 0.006957f
C3665 vdd.n3016 gnd 0.44438f
C3666 vdd.n3017 gnd 0.006957f
C3667 vdd.n3018 gnd 0.006957f
C3668 vdd.n3019 gnd 0.006957f
C3669 vdd.n3020 gnd 0.014897f
C3670 vdd.n3021 gnd 0.014897f
C3671 vdd.n3022 gnd 0.015797f
C3672 vdd.n3023 gnd 0.015797f
C3673 vdd.n3024 gnd 0.006957f
C3674 vdd.n3025 gnd 0.006957f
C3675 vdd.n3026 gnd 0.006957f
C3676 vdd.n3027 gnd 0.005371f
C3677 vdd.n3028 gnd 0.009943f
C3678 vdd.n3029 gnd 0.005065f
C3679 vdd.n3030 gnd 0.006957f
C3680 vdd.n3031 gnd 0.006957f
C3681 vdd.n3032 gnd 0.006957f
C3682 vdd.n3033 gnd 0.006957f
C3683 vdd.n3034 gnd 0.006957f
C3684 vdd.n3035 gnd 0.006957f
C3685 vdd.n3036 gnd 0.006957f
C3686 vdd.n3037 gnd 0.006957f
C3687 vdd.n3038 gnd 0.006957f
C3688 vdd.n3039 gnd 0.006957f
C3689 vdd.n3040 gnd 0.006957f
C3690 vdd.n3041 gnd 0.006957f
C3691 vdd.n3042 gnd 0.006957f
C3692 vdd.n3043 gnd 0.006957f
C3693 vdd.n3044 gnd 0.006957f
C3694 vdd.n3045 gnd 0.006957f
C3695 vdd.n3046 gnd 0.006957f
C3696 vdd.n3047 gnd 0.006957f
C3697 vdd.n3048 gnd 0.006957f
C3698 vdd.n3049 gnd 0.006957f
C3699 vdd.n3050 gnd 0.006957f
C3700 vdd.n3051 gnd 0.006957f
C3701 vdd.n3052 gnd 0.006957f
C3702 vdd.n3053 gnd 0.006957f
C3703 vdd.n3054 gnd 0.006957f
C3704 vdd.n3055 gnd 0.006957f
C3705 vdd.n3056 gnd 0.006957f
C3706 vdd.n3057 gnd 0.006957f
C3707 vdd.n3058 gnd 0.006957f
C3708 vdd.n3059 gnd 0.006957f
C3709 vdd.n3060 gnd 0.006957f
C3710 vdd.n3061 gnd 0.006957f
C3711 vdd.n3062 gnd 0.006957f
C3712 vdd.n3063 gnd 0.006957f
C3713 vdd.n3064 gnd 0.006957f
C3714 vdd.n3065 gnd 0.006957f
C3715 vdd.n3066 gnd 0.006957f
C3716 vdd.n3067 gnd 0.006957f
C3717 vdd.n3068 gnd 0.006957f
C3718 vdd.n3069 gnd 0.006957f
C3719 vdd.n3070 gnd 0.006957f
C3720 vdd.n3071 gnd 0.006957f
C3721 vdd.n3072 gnd 0.006957f
C3722 vdd.n3073 gnd 0.006957f
C3723 vdd.n3074 gnd 0.006957f
C3724 vdd.n3075 gnd 0.006957f
C3725 vdd.n3076 gnd 0.006957f
C3726 vdd.n3077 gnd 0.006957f
C3727 vdd.n3078 gnd 0.006957f
C3728 vdd.n3079 gnd 0.006957f
C3729 vdd.n3080 gnd 0.006957f
C3730 vdd.n3081 gnd 0.006957f
C3731 vdd.n3082 gnd 0.006957f
C3732 vdd.n3083 gnd 0.006957f
C3733 vdd.n3084 gnd 0.006957f
C3734 vdd.n3085 gnd 0.006957f
C3735 vdd.n3086 gnd 0.006957f
C3736 vdd.n3087 gnd 0.006957f
C3737 vdd.n3088 gnd 0.867847f
C3738 vdd.n3090 gnd 0.015797f
C3739 vdd.n3091 gnd 0.015797f
C3740 vdd.n3092 gnd 0.014897f
C3741 vdd.n3093 gnd 0.006957f
C3742 vdd.n3094 gnd 0.006957f
C3743 vdd.n3095 gnd 0.41824f
C3744 vdd.n3096 gnd 0.006957f
C3745 vdd.n3097 gnd 0.006957f
C3746 vdd.n3098 gnd 0.006957f
C3747 vdd.n3099 gnd 0.006957f
C3748 vdd.n3100 gnd 0.006957f
C3749 vdd.n3101 gnd 0.423468f
C3750 vdd.n3102 gnd 0.006957f
C3751 vdd.n3103 gnd 0.006957f
C3752 vdd.n3104 gnd 0.006957f
C3753 vdd.n3105 gnd 0.006957f
C3754 vdd.n3106 gnd 0.006957f
C3755 vdd.n3107 gnd 0.711008f
C3756 vdd.n3108 gnd 0.006957f
C3757 vdd.n3109 gnd 0.006957f
C3758 vdd.n3110 gnd 0.006957f
C3759 vdd.n3111 gnd 0.006957f
C3760 vdd.n3112 gnd 0.006957f
C3761 vdd.n3113 gnd 0.512344f
C3762 vdd.n3114 gnd 0.006957f
C3763 vdd.n3115 gnd 0.006957f
C3764 vdd.n3116 gnd 0.006957f
C3765 vdd.n3117 gnd 0.006957f
C3766 vdd.n3118 gnd 0.006957f
C3767 vdd.n3119 gnd 0.643044f
C3768 vdd.n3120 gnd 0.006957f
C3769 vdd.n3121 gnd 0.006957f
C3770 vdd.n3122 gnd 0.006957f
C3771 vdd.n3123 gnd 0.006957f
C3772 vdd.n3124 gnd 0.006957f
C3773 vdd.n3125 gnd 0.528028f
C3774 vdd.n3126 gnd 0.006957f
C3775 vdd.n3127 gnd 0.006957f
C3776 vdd.n3128 gnd 0.006957f
C3777 vdd.n3129 gnd 0.006957f
C3778 vdd.n3130 gnd 0.006957f
C3779 vdd.n3131 gnd 0.371188f
C3780 vdd.n3132 gnd 0.006957f
C3781 vdd.n3133 gnd 0.006957f
C3782 vdd.n3134 gnd 0.006957f
C3783 vdd.n3135 gnd 0.006957f
C3784 vdd.n3136 gnd 0.006957f
C3785 vdd.n3137 gnd 0.224804f
C3786 vdd.n3138 gnd 0.006957f
C3787 vdd.n3139 gnd 0.006957f
C3788 vdd.n3140 gnd 0.006957f
C3789 vdd.n3141 gnd 0.006957f
C3790 vdd.n3142 gnd 0.006957f
C3791 vdd.n3143 gnd 0.6535f
C3792 vdd.n3144 gnd 0.006957f
C3793 vdd.n3145 gnd 0.006957f
C3794 vdd.n3146 gnd 0.006957f
C3795 vdd.n3147 gnd 0.004911f
C3796 vdd.n3148 gnd 0.006957f
C3797 vdd.n3149 gnd 0.006957f
C3798 vdd.n3150 gnd 0.711008f
C3799 vdd.n3151 gnd 0.006957f
C3800 vdd.n3152 gnd 0.006957f
C3801 vdd.n3153 gnd 0.006957f
C3802 vdd.n3154 gnd 0.006957f
C3803 vdd.n3155 gnd 0.006957f
C3804 vdd.n3156 gnd 0.564624f
C3805 vdd.n3157 gnd 0.006957f
C3806 vdd.n3158 gnd 0.005525f
C3807 vdd.n3159 gnd 0.006957f
C3808 vdd.n3160 gnd 0.006957f
C3809 vdd.n3161 gnd 0.006957f
C3810 vdd.n3162 gnd 0.454836f
C3811 vdd.n3163 gnd 0.006957f
C3812 vdd.n3164 gnd 0.006957f
C3813 vdd.n3165 gnd 0.006957f
C3814 vdd.n3166 gnd 0.006957f
C3815 vdd.n3167 gnd 0.006957f
C3816 vdd.n3168 gnd 0.413012f
C3817 vdd.n3169 gnd 0.006957f
C3818 vdd.n3170 gnd 0.006957f
C3819 vdd.n3171 gnd 0.006957f
C3820 vdd.n3172 gnd 0.006957f
C3821 vdd.n3173 gnd 0.006957f
C3822 vdd.n3174 gnd 0.569852f
C3823 vdd.n3175 gnd 0.006957f
C3824 vdd.n3176 gnd 0.006957f
C3825 vdd.n3177 gnd 0.006957f
C3826 vdd.n3178 gnd 0.006957f
C3827 vdd.n3179 gnd 0.006957f
C3828 vdd.n3180 gnd 0.711008f
C3829 vdd.n3181 gnd 0.006957f
C3830 vdd.n3182 gnd 0.006957f
C3831 vdd.n3183 gnd 0.006957f
C3832 vdd.n3184 gnd 0.006957f
C3833 vdd.n3185 gnd 0.006957f
C3834 vdd.n3186 gnd 0.695324f
C3835 vdd.n3187 gnd 0.006957f
C3836 vdd.n3188 gnd 0.006957f
C3837 vdd.n3189 gnd 0.006957f
C3838 vdd.n3190 gnd 0.006957f
C3839 vdd.n3191 gnd 0.006957f
C3840 vdd.n3192 gnd 0.538484f
C3841 vdd.n3193 gnd 0.006957f
C3842 vdd.n3194 gnd 0.006957f
C3843 vdd.n3195 gnd 0.006957f
C3844 vdd.n3196 gnd 0.006957f
C3845 vdd.n3197 gnd 0.006957f
C3846 vdd.n3198 gnd 0.381644f
C3847 vdd.n3199 gnd 0.006957f
C3848 vdd.n3200 gnd 0.006957f
C3849 vdd.n3201 gnd 0.006957f
C3850 vdd.n3202 gnd 0.006957f
C3851 vdd.n3203 gnd 0.006957f
C3852 vdd.n3204 gnd 0.711008f
C3853 vdd.n3205 gnd 0.006957f
C3854 vdd.n3206 gnd 0.006957f
C3855 vdd.n3207 gnd 0.006957f
C3856 vdd.n3208 gnd 0.006957f
C3857 vdd.n3209 gnd 0.006957f
C3858 vdd.n3210 gnd 0.006957f
C3859 vdd.n3212 gnd 0.006957f
C3860 vdd.n3213 gnd 0.006957f
C3861 vdd.n3215 gnd 0.006957f
C3862 vdd.n3216 gnd 0.006957f
C3863 vdd.n3219 gnd 0.006957f
C3864 vdd.n3220 gnd 0.006957f
C3865 vdd.n3221 gnd 0.006957f
C3866 vdd.n3222 gnd 0.006957f
C3867 vdd.n3224 gnd 0.006957f
C3868 vdd.n3225 gnd 0.006957f
C3869 vdd.n3226 gnd 0.006957f
C3870 vdd.n3227 gnd 0.006957f
C3871 vdd.n3228 gnd 0.006957f
C3872 vdd.n3229 gnd 0.006957f
C3873 vdd.n3231 gnd 0.006957f
C3874 vdd.n3232 gnd 0.006957f
C3875 vdd.n3233 gnd 0.006957f
C3876 vdd.n3234 gnd 0.006957f
C3877 vdd.n3235 gnd 0.006957f
C3878 vdd.n3236 gnd 0.006957f
C3879 vdd.n3238 gnd 0.006957f
C3880 vdd.n3239 gnd 0.006957f
C3881 vdd.n3240 gnd 0.006957f
C3882 vdd.n3241 gnd 0.006957f
C3883 vdd.n3242 gnd 0.006957f
C3884 vdd.n3243 gnd 0.006957f
C3885 vdd.n3245 gnd 0.006957f
C3886 vdd.n3246 gnd 0.015797f
C3887 vdd.n3247 gnd 0.015797f
C3888 vdd.n3248 gnd 0.014897f
C3889 vdd.n3249 gnd 0.006957f
C3890 vdd.n3250 gnd 0.006957f
C3891 vdd.n3251 gnd 0.006957f
C3892 vdd.n3252 gnd 0.006957f
C3893 vdd.n3253 gnd 0.006957f
C3894 vdd.n3254 gnd 0.006957f
C3895 vdd.n3255 gnd 0.711008f
C3896 vdd.n3256 gnd 0.006957f
C3897 vdd.n3257 gnd 0.006957f
C3898 vdd.n3258 gnd 0.006957f
C3899 vdd.n3259 gnd 0.006957f
C3900 vdd.n3260 gnd 0.006957f
C3901 vdd.n3261 gnd 0.507116f
C3902 vdd.n3262 gnd 0.006957f
C3903 vdd.n3263 gnd 0.006957f
C3904 vdd.n3264 gnd 0.006957f
C3905 vdd.n3265 gnd 0.015797f
C3906 vdd.n3266 gnd 0.014897f
C3907 vdd.n3267 gnd 0.015797f
C3908 vdd.n3269 gnd 0.006957f
C3909 vdd.n3270 gnd 0.006957f
C3910 vdd.n3271 gnd 0.005371f
C3911 vdd.n3272 gnd 0.009943f
C3912 vdd.n3273 gnd 0.005065f
C3913 vdd.n3274 gnd 0.006957f
C3914 vdd.n3275 gnd 0.006957f
C3915 vdd.n3277 gnd 0.006957f
C3916 vdd.n3278 gnd 0.006957f
C3917 vdd.n3279 gnd 0.006957f
C3918 vdd.n3280 gnd 0.006957f
C3919 vdd.n3281 gnd 0.006957f
C3920 vdd.n3282 gnd 0.006957f
C3921 vdd.n3284 gnd 0.006957f
C3922 vdd.n3285 gnd 0.006957f
C3923 vdd.n3286 gnd 0.006957f
C3924 vdd.n3287 gnd 0.006957f
C3925 vdd.n3288 gnd 0.006957f
C3926 vdd.n3289 gnd 0.006957f
C3927 vdd.n3291 gnd 0.006957f
C3928 vdd.n3292 gnd 0.006957f
C3929 vdd.n3293 gnd 0.006957f
C3930 vdd.n3294 gnd 0.006957f
C3931 vdd.n3295 gnd 0.006957f
C3932 vdd.n3296 gnd 0.006957f
C3933 vdd.n3298 gnd 0.006957f
C3934 vdd.n3299 gnd 0.006957f
C3935 vdd.n3300 gnd 0.006957f
C3936 vdd.n3302 gnd 0.006957f
C3937 vdd.n3303 gnd 0.006957f
C3938 vdd.n3304 gnd 0.006957f
C3939 vdd.n3305 gnd 0.006957f
C3940 vdd.n3306 gnd 0.006957f
C3941 vdd.n3307 gnd 0.006957f
C3942 vdd.n3309 gnd 0.006957f
C3943 vdd.n3310 gnd 0.006957f
C3944 vdd.n3311 gnd 0.006957f
C3945 vdd.n3312 gnd 0.006957f
C3946 vdd.n3313 gnd 0.006957f
C3947 vdd.n3314 gnd 0.006957f
C3948 vdd.n3316 gnd 0.006957f
C3949 vdd.n3317 gnd 0.006957f
C3950 vdd.n3318 gnd 0.006957f
C3951 vdd.n3319 gnd 0.006957f
C3952 vdd.n3320 gnd 0.006957f
C3953 vdd.n3321 gnd 0.006957f
C3954 vdd.n3323 gnd 0.006957f
C3955 vdd.n3324 gnd 0.006957f
C3956 vdd.n3326 gnd 0.006957f
C3957 vdd.n3327 gnd 0.006957f
C3958 vdd.n3328 gnd 0.015797f
C3959 vdd.n3329 gnd 0.014897f
C3960 vdd.n3330 gnd 0.014897f
C3961 vdd.n3331 gnd 0.961951f
C3962 vdd.n3332 gnd 0.014897f
C3963 vdd.n3333 gnd 0.015797f
C3964 vdd.n3334 gnd 0.014897f
C3965 vdd.n3335 gnd 0.006957f
C3966 vdd.n3336 gnd 0.005371f
C3967 vdd.n3337 gnd 0.006957f
C3968 vdd.n3339 gnd 0.006957f
C3969 vdd.n3340 gnd 0.006957f
C3970 vdd.n3341 gnd 0.006957f
C3971 vdd.n3342 gnd 0.006957f
C3972 vdd.n3343 gnd 0.006957f
C3973 vdd.n3344 gnd 0.006957f
C3974 vdd.n3346 gnd 0.006957f
C3975 vdd.n3347 gnd 0.006957f
C3976 vdd.n3348 gnd 0.006957f
C3977 vdd.n3349 gnd 0.006957f
C3978 vdd.n3350 gnd 0.006957f
C3979 vdd.n3351 gnd 0.006957f
C3980 vdd.n3353 gnd 0.006957f
C3981 vdd.n3354 gnd 0.006957f
C3982 vdd.n3355 gnd 0.006957f
C3983 vdd.n3356 gnd 0.006957f
C3984 vdd.n3357 gnd 0.006957f
C3985 vdd.n3358 gnd 0.006957f
C3986 vdd.n3360 gnd 0.006957f
C3987 vdd.n3361 gnd 0.006957f
C3988 vdd.n3363 gnd 0.006957f
C3989 vdd.n3364 gnd 0.042961f
C3990 vdd.n3365 gnd 1.09007f
C3991 vdd.n3367 gnd 0.004323f
C3992 vdd.n3368 gnd 0.008235f
C3993 vdd.n3369 gnd 0.010231f
C3994 vdd.n3370 gnd 0.010231f
C3995 vdd.n3371 gnd 0.008235f
C3996 vdd.n3372 gnd 0.008235f
C3997 vdd.n3373 gnd 0.010231f
C3998 vdd.n3374 gnd 0.010231f
C3999 vdd.n3375 gnd 0.008235f
C4000 vdd.n3376 gnd 0.008235f
C4001 vdd.n3377 gnd 0.010231f
C4002 vdd.n3378 gnd 0.010231f
C4003 vdd.n3379 gnd 0.008235f
C4004 vdd.n3380 gnd 0.008235f
C4005 vdd.n3381 gnd 0.010231f
C4006 vdd.n3382 gnd 0.010231f
C4007 vdd.n3383 gnd 0.008235f
C4008 vdd.n3384 gnd 0.008235f
C4009 vdd.n3385 gnd 0.010231f
C4010 vdd.n3386 gnd 0.010231f
C4011 vdd.n3387 gnd 0.008235f
C4012 vdd.n3388 gnd 0.008235f
C4013 vdd.n3389 gnd 0.010231f
C4014 vdd.n3390 gnd 0.010231f
C4015 vdd.n3391 gnd 0.008235f
C4016 vdd.n3392 gnd 0.008235f
C4017 vdd.n3393 gnd 0.010231f
C4018 vdd.n3394 gnd 0.010231f
C4019 vdd.n3395 gnd 0.008235f
C4020 vdd.n3396 gnd 0.008235f
C4021 vdd.n3397 gnd 0.010231f
C4022 vdd.n3398 gnd 0.010231f
C4023 vdd.n3399 gnd 0.008235f
C4024 vdd.n3400 gnd 0.008235f
C4025 vdd.n3401 gnd 0.010231f
C4026 vdd.n3402 gnd 0.010231f
C4027 vdd.n3403 gnd 0.008235f
C4028 vdd.n3404 gnd 0.010231f
C4029 vdd.n3405 gnd 0.010231f
C4030 vdd.n3406 gnd 0.008235f
C4031 vdd.n3407 gnd 0.010231f
C4032 vdd.n3408 gnd 0.010231f
C4033 vdd.n3409 gnd 0.010231f
C4034 vdd.n3410 gnd 0.016799f
C4035 vdd.n3411 gnd 0.010231f
C4036 vdd.n3412 gnd 0.010231f
C4037 vdd.n3413 gnd 0.0056f
C4038 vdd.n3414 gnd 0.008235f
C4039 vdd.n3415 gnd 0.010231f
C4040 vdd.n3416 gnd 0.010231f
C4041 vdd.n3417 gnd 0.008235f
C4042 vdd.n3418 gnd 0.008235f
C4043 vdd.n3419 gnd 0.010231f
C4044 vdd.n3420 gnd 0.010231f
C4045 vdd.n3421 gnd 0.008235f
C4046 vdd.n3422 gnd 0.008235f
C4047 vdd.n3423 gnd 0.010231f
C4048 vdd.n3424 gnd 0.010231f
C4049 vdd.n3425 gnd 0.008235f
C4050 vdd.n3426 gnd 0.008235f
C4051 vdd.n3427 gnd 0.010231f
C4052 vdd.n3428 gnd 0.010231f
C4053 vdd.n3429 gnd 0.008235f
C4054 vdd.n3430 gnd 0.008235f
C4055 vdd.n3431 gnd 0.010231f
C4056 vdd.n3432 gnd 0.010231f
C4057 vdd.n3433 gnd 0.008235f
C4058 vdd.n3434 gnd 0.008235f
C4059 vdd.n3435 gnd 0.010231f
C4060 vdd.n3436 gnd 0.010231f
C4061 vdd.n3437 gnd 0.008235f
C4062 vdd.n3438 gnd 0.008235f
C4063 vdd.n3439 gnd 0.010231f
C4064 vdd.n3440 gnd 0.010231f
C4065 vdd.n3441 gnd 0.008235f
C4066 vdd.n3442 gnd 0.008235f
C4067 vdd.n3443 gnd 0.010231f
C4068 vdd.n3444 gnd 0.010231f
C4069 vdd.n3445 gnd 0.008235f
C4070 vdd.n3446 gnd 0.008235f
C4071 vdd.n3447 gnd 0.010231f
C4072 vdd.n3448 gnd 0.010231f
C4073 vdd.n3449 gnd 0.008235f
C4074 vdd.n3450 gnd 0.010231f
C4075 vdd.n3451 gnd 0.010231f
C4076 vdd.n3452 gnd 0.008235f
C4077 vdd.n3453 gnd 0.010231f
C4078 vdd.n3454 gnd 0.010231f
C4079 vdd.n3455 gnd 0.010231f
C4080 vdd.t210 gnd 0.125873f
C4081 vdd.t211 gnd 0.134524f
C4082 vdd.t209 gnd 0.164388f
C4083 vdd.n3456 gnd 0.210723f
C4084 vdd.n3457 gnd 0.177045f
C4085 vdd.n3458 gnd 0.016799f
C4086 vdd.n3459 gnd 0.010231f
C4087 vdd.n3460 gnd 0.010231f
C4088 vdd.n3461 gnd 0.006876f
C4089 vdd.n3462 gnd 0.008235f
C4090 vdd.n3463 gnd 0.010231f
C4091 vdd.n3464 gnd 0.010231f
C4092 vdd.n3465 gnd 0.008235f
C4093 vdd.n3466 gnd 0.008235f
C4094 vdd.n3467 gnd 0.010231f
C4095 vdd.n3468 gnd 0.010231f
C4096 vdd.n3469 gnd 0.008235f
C4097 vdd.n3470 gnd 0.008235f
C4098 vdd.n3471 gnd 0.010231f
C4099 vdd.n3472 gnd 0.010231f
C4100 vdd.n3473 gnd 0.008235f
C4101 vdd.n3474 gnd 0.008235f
C4102 vdd.n3475 gnd 0.010231f
C4103 vdd.n3476 gnd 0.010231f
C4104 vdd.n3477 gnd 0.008235f
C4105 vdd.n3478 gnd 0.008235f
C4106 vdd.n3479 gnd 0.010231f
C4107 vdd.n3480 gnd 0.010231f
C4108 vdd.n3481 gnd 0.008235f
C4109 vdd.n3482 gnd 0.008235f
C4110 vdd.n3483 gnd 0.010231f
C4111 vdd.n3484 gnd 0.010231f
C4112 vdd.n3485 gnd 0.008235f
C4113 vdd.n3486 gnd 0.008235f
C4114 vdd.n3488 gnd 1.09007f
C4115 vdd.n3490 gnd 0.008235f
C4116 vdd.n3491 gnd 0.008235f
C4117 vdd.n3492 gnd 0.006835f
C4118 vdd.n3493 gnd 0.025281f
C4119 vdd.n3495 gnd 12.7668f
C4120 vdd.n3496 gnd 0.025281f
C4121 vdd.n3497 gnd 0.003912f
C4122 vdd.n3498 gnd 0.025281f
C4123 vdd.n3499 gnd 0.024751f
C4124 vdd.n3500 gnd 0.010231f
C4125 vdd.n3501 gnd 0.008235f
C4126 vdd.n3502 gnd 0.010231f
C4127 vdd.n3503 gnd 0.632588f
C4128 vdd.n3504 gnd 0.010231f
C4129 vdd.n3505 gnd 0.008235f
C4130 vdd.n3506 gnd 0.010231f
C4131 vdd.n3507 gnd 0.010231f
C4132 vdd.n3508 gnd 0.010231f
C4133 vdd.n3509 gnd 0.008235f
C4134 vdd.n3510 gnd 0.010231f
C4135 vdd.n3511 gnd 1.0456f
C4136 vdd.n3512 gnd 0.010231f
C4137 vdd.n3513 gnd 0.008235f
C4138 vdd.n3514 gnd 0.010231f
C4139 vdd.n3515 gnd 0.010231f
C4140 vdd.n3516 gnd 0.010231f
C4141 vdd.n3517 gnd 0.008235f
C4142 vdd.n3518 gnd 0.010231f
C4143 vdd.n3519 gnd 0.674412f
C4144 vdd.n3520 gnd 0.716236f
C4145 vdd.n3521 gnd 0.010231f
C4146 vdd.n3522 gnd 0.008235f
C4147 vdd.n3523 gnd 0.010231f
C4148 vdd.n3524 gnd 0.010231f
C4149 vdd.n3525 gnd 0.010231f
C4150 vdd.n3526 gnd 0.008235f
C4151 vdd.n3527 gnd 0.010231f
C4152 vdd.n3528 gnd 0.867847f
C4153 vdd.n3529 gnd 0.010231f
C4154 vdd.n3530 gnd 0.008235f
C4155 vdd.n3531 gnd 0.010231f
C4156 vdd.n3532 gnd 0.010231f
C4157 vdd.n3533 gnd 0.010231f
C4158 vdd.n3534 gnd 0.008235f
C4159 vdd.n3535 gnd 0.010231f
C4160 vdd.t25 gnd 0.5228f
C4161 vdd.n3536 gnd 0.841707f
C4162 vdd.n3537 gnd 0.010231f
C4163 vdd.n3538 gnd 0.008235f
C4164 vdd.n3539 gnd 0.010231f
C4165 vdd.n3540 gnd 0.010231f
C4166 vdd.n3541 gnd 0.010231f
C4167 vdd.n3542 gnd 0.008235f
C4168 vdd.n3543 gnd 0.010231f
C4169 vdd.n3544 gnd 0.663956f
C4170 vdd.n3545 gnd 0.010231f
C4171 vdd.n3546 gnd 0.008235f
C4172 vdd.n3547 gnd 0.010231f
C4173 vdd.n3548 gnd 0.010231f
C4174 vdd.n3549 gnd 0.010231f
C4175 vdd.n3550 gnd 0.008235f
C4176 vdd.n3551 gnd 0.010231f
C4177 vdd.n3552 gnd 0.831251f
C4178 vdd.n3553 gnd 0.559396f
C4179 vdd.n3554 gnd 0.010231f
C4180 vdd.n3555 gnd 0.008235f
C4181 vdd.n3556 gnd 0.010231f
C4182 vdd.n3557 gnd 0.010231f
C4183 vdd.n3558 gnd 0.010231f
C4184 vdd.n3559 gnd 0.008235f
C4185 vdd.n3560 gnd 0.010231f
C4186 vdd.n3561 gnd 0.737148f
C4187 vdd.n3562 gnd 0.010231f
C4188 vdd.n3563 gnd 0.008235f
C4189 vdd.n3564 gnd 0.010231f
C4190 vdd.n3565 gnd 0.010231f
C4191 vdd.n3566 gnd 0.010231f
C4192 vdd.n3567 gnd 0.010231f
C4193 vdd.n3568 gnd 0.010231f
C4194 vdd.n3569 gnd 0.008235f
C4195 vdd.n3570 gnd 0.008235f
C4196 vdd.n3571 gnd 0.010231f
C4197 vdd.t6 gnd 0.5228f
C4198 vdd.n3572 gnd 0.867847f
C4199 vdd.n3573 gnd 0.010231f
C4200 vdd.n3574 gnd 0.008235f
C4201 vdd.n3575 gnd 0.010231f
C4202 vdd.n3576 gnd 0.010231f
C4203 vdd.n3577 gnd 0.010231f
C4204 vdd.n3578 gnd 0.008235f
C4205 vdd.n3579 gnd 0.010231f
C4206 vdd.n3580 gnd 0.820795f
C4207 vdd.n3581 gnd 0.010231f
C4208 vdd.n3582 gnd 0.010231f
C4209 vdd.n3583 gnd 0.008235f
C4210 vdd.n3584 gnd 0.008235f
C4211 vdd.n3585 gnd 0.010231f
C4212 vdd.n3586 gnd 0.010231f
C4213 vdd.n3587 gnd 0.010231f
C4214 vdd.n3588 gnd 0.008235f
C4215 vdd.n3589 gnd 0.010231f
C4216 vdd.n3590 gnd 0.008235f
C4217 vdd.n3591 gnd 0.008235f
C4218 vdd.n3592 gnd 0.010231f
C4219 vdd.n3593 gnd 0.010231f
C4220 vdd.n3594 gnd 0.010231f
C4221 vdd.n3595 gnd 0.008235f
C4222 vdd.n3596 gnd 0.010231f
C4223 vdd.n3597 gnd 0.008235f
C4224 vdd.n3598 gnd 0.008235f
C4225 vdd.n3599 gnd 0.010231f
C4226 vdd.n3600 gnd 0.010231f
C4227 vdd.n3601 gnd 0.010231f
C4228 vdd.n3602 gnd 0.008235f
C4229 vdd.n3603 gnd 0.867847f
C4230 vdd.n3604 gnd 0.010231f
C4231 vdd.n3605 gnd 0.008235f
C4232 vdd.n3606 gnd 0.008235f
C4233 vdd.n3607 gnd 0.010231f
C4234 vdd.n3608 gnd 0.010231f
C4235 vdd.n3609 gnd 0.010231f
C4236 vdd.n3610 gnd 0.008235f
C4237 vdd.n3611 gnd 0.010231f
C4238 vdd.n3612 gnd 0.008235f
C4239 vdd.n3613 gnd 0.008235f
C4240 vdd.n3614 gnd 0.010231f
C4241 vdd.n3615 gnd 0.010231f
C4242 vdd.n3616 gnd 0.010231f
C4243 vdd.n3617 gnd 0.008235f
C4244 vdd.n3618 gnd 0.010231f
C4245 vdd.n3619 gnd 0.008235f
C4246 vdd.n3620 gnd 0.006835f
C4247 vdd.n3621 gnd 0.024751f
C4248 vdd.n3622 gnd 0.025281f
C4249 vdd.n3623 gnd 0.003912f
C4250 vdd.n3624 gnd 0.025281f
C4251 vdd.n3626 gnd 2.47807f
C4252 vdd.n3627 gnd 1.54226f
C4253 vdd.n3628 gnd 0.024751f
C4254 vdd.n3629 gnd 0.006835f
C4255 vdd.n3630 gnd 0.008235f
C4256 vdd.n3631 gnd 0.008235f
C4257 vdd.n3632 gnd 0.010231f
C4258 vdd.n3633 gnd 1.0456f
C4259 vdd.n3634 gnd 1.0456f
C4260 vdd.n3635 gnd 0.956723f
C4261 vdd.n3636 gnd 0.010231f
C4262 vdd.n3637 gnd 0.008235f
C4263 vdd.n3638 gnd 0.008235f
C4264 vdd.n3639 gnd 0.008235f
C4265 vdd.n3640 gnd 0.010231f
C4266 vdd.n3641 gnd 0.778971f
C4267 vdd.t12 gnd 0.5228f
C4268 vdd.n3642 gnd 0.789427f
C4269 vdd.n3643 gnd 0.60122f
C4270 vdd.n3644 gnd 0.010231f
C4271 vdd.n3645 gnd 0.008235f
C4272 vdd.n3646 gnd 0.008235f
C4273 vdd.n3647 gnd 0.008235f
C4274 vdd.n3648 gnd 0.010231f
C4275 vdd.n3649 gnd 0.622132f
C4276 vdd.n3650 gnd 0.768516f
C4277 vdd.t20 gnd 0.5228f
C4278 vdd.n3651 gnd 0.799883f
C4279 vdd.n3652 gnd 0.010231f
C4280 vdd.n3653 gnd 0.008235f
C4281 vdd.n3654 gnd 0.008235f
C4282 vdd.n3655 gnd 0.008235f
C4283 vdd.n3656 gnd 0.010231f
C4284 vdd.n3657 gnd 0.867847f
C4285 vdd.t74 gnd 0.5228f
C4286 vdd.n3658 gnd 0.632588f
C4287 vdd.n3659 gnd 0.75806f
C4288 vdd.n3660 gnd 0.010231f
C4289 vdd.n3661 gnd 0.008235f
C4290 vdd.n3662 gnd 0.008235f
C4291 vdd.n3663 gnd 0.008235f
C4292 vdd.n3664 gnd 0.010231f
C4293 vdd.n3665 gnd 0.580308f
C4294 vdd.t18 gnd 0.5228f
C4295 vdd.n3666 gnd 0.867847f
C4296 vdd.t116 gnd 0.5228f
C4297 vdd.n3667 gnd 0.643044f
C4298 vdd.n3668 gnd 0.010231f
C4299 vdd.n3669 gnd 0.008235f
C4300 vdd.n3670 gnd 0.007863f
C4301 vdd.n3671 gnd 0.603486f
C4302 vdd.n3672 gnd 2.98812f
C4303 a_n2982_13878.n0 gnd 2.53375f
C4304 a_n2982_13878.n1 gnd 3.78544f
C4305 a_n2982_13878.n2 gnd 3.42814f
C4306 a_n2982_13878.n3 gnd 0.971817f
C4307 a_n2982_13878.n4 gnd 0.20945f
C4308 a_n2982_13878.n5 gnd 0.20945f
C4309 a_n2982_13878.n6 gnd 0.458034f
C4310 a_n2982_13878.n7 gnd 0.20945f
C4311 a_n2982_13878.n8 gnd 0.27462f
C4312 a_n2982_13878.n9 gnd 0.20945f
C4313 a_n2982_13878.n10 gnd 0.20945f
C4314 a_n2982_13878.n11 gnd 0.791576f
C4315 a_n2982_13878.n12 gnd 0.20945f
C4316 a_n2982_13878.n13 gnd 0.904041f
C4317 a_n2982_13878.n14 gnd 0.198733f
C4318 a_n2982_13878.n15 gnd 0.146371f
C4319 a_n2982_13878.n16 gnd 0.230048f
C4320 a_n2982_13878.n17 gnd 0.177686f
C4321 a_n2982_13878.n18 gnd 0.198733f
C4322 a_n2982_13878.n19 gnd 0.146371f
C4323 a_n2982_13878.n20 gnd 0.956403f
C4324 a_n2982_13878.n21 gnd 0.20945f
C4325 a_n2982_13878.n22 gnd 0.73719f
C4326 a_n2982_13878.n23 gnd 0.20945f
C4327 a_n2982_13878.n24 gnd 0.20945f
C4328 a_n2982_13878.n25 gnd 0.477018f
C4329 a_n2982_13878.n26 gnd 0.27462f
C4330 a_n2982_13878.n27 gnd 0.20945f
C4331 a_n2982_13878.n28 gnd 0.529381f
C4332 a_n2982_13878.n29 gnd 0.20945f
C4333 a_n2982_13878.n30 gnd 0.20945f
C4334 a_n2982_13878.n31 gnd 0.931898f
C4335 a_n2982_13878.n32 gnd 0.27462f
C4336 a_n2982_13878.n33 gnd 3.08362f
C4337 a_n2982_13878.n34 gnd 0.27462f
C4338 a_n2982_13878.n35 gnd 1.16191f
C4339 a_n2982_13878.n36 gnd 2.12168f
C4340 a_n2982_13878.n37 gnd 1.72437f
C4341 a_n2982_13878.n38 gnd 1.16191f
C4342 a_n2982_13878.n39 gnd 1.72437f
C4343 a_n2982_13878.n40 gnd 2.32061f
C4344 a_n2982_13878.n41 gnd 0.008404f
C4345 a_n2982_13878.n42 gnd 4.05e-19
C4346 a_n2982_13878.n44 gnd 0.008109f
C4347 a_n2982_13878.n45 gnd 0.011792f
C4348 a_n2982_13878.n46 gnd 0.007801f
C4349 a_n2982_13878.n48 gnd 0.277816f
C4350 a_n2982_13878.n49 gnd 0.008404f
C4351 a_n2982_13878.n50 gnd 4.05e-19
C4352 a_n2982_13878.n52 gnd 0.008109f
C4353 a_n2982_13878.n53 gnd 0.011792f
C4354 a_n2982_13878.n54 gnd 0.007801f
C4355 a_n2982_13878.n56 gnd 0.277816f
C4356 a_n2982_13878.n57 gnd 0.008109f
C4357 a_n2982_13878.n58 gnd 0.276683f
C4358 a_n2982_13878.n59 gnd 0.008109f
C4359 a_n2982_13878.n60 gnd 0.276683f
C4360 a_n2982_13878.n61 gnd 0.008109f
C4361 a_n2982_13878.n62 gnd 0.276683f
C4362 a_n2982_13878.n63 gnd 0.008109f
C4363 a_n2982_13878.n64 gnd 1.64574f
C4364 a_n2982_13878.n65 gnd 0.276683f
C4365 a_n2982_13878.n66 gnd 0.277816f
C4366 a_n2982_13878.n68 gnd 0.007801f
C4367 a_n2982_13878.n69 gnd 0.011792f
C4368 a_n2982_13878.n70 gnd 0.008109f
C4369 a_n2982_13878.n72 gnd 4.05e-19
C4370 a_n2982_13878.n73 gnd 0.008404f
C4371 a_n2982_13878.n74 gnd 0.104725f
C4372 a_n2982_13878.n75 gnd 0.008404f
C4373 a_n2982_13878.n76 gnd 4.05e-19
C4374 a_n2982_13878.n78 gnd 0.008109f
C4375 a_n2982_13878.n79 gnd 0.011792f
C4376 a_n2982_13878.n80 gnd 0.007801f
C4377 a_n2982_13878.n82 gnd 0.277816f
C4378 a_n2982_13878.t36 gnd 0.145277f
C4379 a_n2982_13878.t42 gnd 1.3603f
C4380 a_n2982_13878.t18 gnd 0.145277f
C4381 a_n2982_13878.t40 gnd 0.145277f
C4382 a_n2982_13878.n83 gnd 1.02333f
C4383 a_n2982_13878.t23 gnd 0.675756f
C4384 a_n2982_13878.n84 gnd 0.29709f
C4385 a_n2982_13878.t37 gnd 0.675756f
C4386 a_n2982_13878.t51 gnd 0.675756f
C4387 a_n2982_13878.n85 gnd 0.288167f
C4388 a_n2982_13878.t35 gnd 0.675756f
C4389 a_n2982_13878.n86 gnd 0.299644f
C4390 a_n2982_13878.t45 gnd 0.675756f
C4391 a_n2982_13878.t39 gnd 0.675756f
C4392 a_n2982_13878.n87 gnd 0.293009f
C4393 a_n2982_13878.t41 gnd 0.689824f
C4394 a_n2982_13878.t78 gnd 0.675756f
C4395 a_n2982_13878.n88 gnd 0.29709f
C4396 a_n2982_13878.t88 gnd 0.675756f
C4397 a_n2982_13878.t93 gnd 0.675756f
C4398 a_n2982_13878.n89 gnd 0.288167f
C4399 a_n2982_13878.t97 gnd 0.675756f
C4400 a_n2982_13878.n90 gnd 0.299644f
C4401 a_n2982_13878.t68 gnd 0.675756f
C4402 a_n2982_13878.t71 gnd 0.675756f
C4403 a_n2982_13878.n91 gnd 0.293009f
C4404 a_n2982_13878.t101 gnd 0.689824f
C4405 a_n2982_13878.t29 gnd 0.686627f
C4406 a_n2982_13878.t47 gnd 0.675756f
C4407 a_n2982_13878.t49 gnd 0.675756f
C4408 a_n2982_13878.t25 gnd 0.675756f
C4409 a_n2982_13878.n92 gnd 0.293584f
C4410 a_n2982_13878.t53 gnd 0.675756f
C4411 a_n2982_13878.t13 gnd 0.675756f
C4412 a_n2982_13878.t19 gnd 0.675756f
C4413 a_n2982_13878.n93 gnd 0.297105f
C4414 a_n2982_13878.t27 gnd 0.675756f
C4415 a_n2982_13878.t55 gnd 0.675756f
C4416 a_n2982_13878.t21 gnd 0.675756f
C4417 a_n2982_13878.n94 gnd 0.293009f
C4418 a_n2982_13878.t31 gnd 0.675756f
C4419 a_n2982_13878.t33 gnd 0.689824f
C4420 a_n2982_13878.t102 gnd 0.689824f
C4421 a_n2982_13878.t79 gnd 0.675756f
C4422 a_n2982_13878.t84 gnd 0.675756f
C4423 a_n2982_13878.t72 gnd 0.675756f
C4424 a_n2982_13878.n95 gnd 0.296972f
C4425 a_n2982_13878.t89 gnd 0.675756f
C4426 a_n2982_13878.t98 gnd 0.675756f
C4427 a_n2982_13878.t99 gnd 0.675756f
C4428 a_n2982_13878.n96 gnd 0.293332f
C4429 a_n2982_13878.t66 gnd 0.675756f
C4430 a_n2982_13878.t81 gnd 0.675756f
C4431 a_n2982_13878.t69 gnd 0.675756f
C4432 a_n2982_13878.n97 gnd 0.29709f
C4433 a_n2982_13878.t76 gnd 0.675756f
C4434 a_n2982_13878.t95 gnd 0.686627f
C4435 a_n2982_13878.n98 gnd 0.299206f
C4436 a_n2982_13878.n99 gnd 0.293584f
C4437 a_n2982_13878.n100 gnd 0.288167f
C4438 a_n2982_13878.n101 gnd 0.297105f
C4439 a_n2982_13878.n102 gnd 0.299644f
C4440 a_n2982_13878.n103 gnd 0.293009f
C4441 a_n2982_13878.n104 gnd 0.299205f
C4442 a_n2982_13878.t2 gnd 0.112993f
C4443 a_n2982_13878.t6 gnd 0.112993f
C4444 a_n2982_13878.n105 gnd 1.00066f
C4445 a_n2982_13878.t9 gnd 0.112993f
C4446 a_n2982_13878.t4 gnd 0.112993f
C4447 a_n2982_13878.n106 gnd 0.998444f
C4448 a_n2982_13878.t10 gnd 0.112993f
C4449 a_n2982_13878.t1 gnd 0.112993f
C4450 a_n2982_13878.n107 gnd 1.00066f
C4451 a_n2982_13878.t8 gnd 0.112993f
C4452 a_n2982_13878.t0 gnd 0.112993f
C4453 a_n2982_13878.n108 gnd 0.998444f
C4454 a_n2982_13878.t7 gnd 0.112993f
C4455 a_n2982_13878.t59 gnd 0.112993f
C4456 a_n2982_13878.n109 gnd 0.998444f
C4457 a_n2982_13878.t60 gnd 0.112993f
C4458 a_n2982_13878.t63 gnd 0.112993f
C4459 a_n2982_13878.n110 gnd 0.998444f
C4460 a_n2982_13878.t62 gnd 0.112993f
C4461 a_n2982_13878.t3 gnd 0.112993f
C4462 a_n2982_13878.n111 gnd 1.00066f
C4463 a_n2982_13878.t5 gnd 0.112993f
C4464 a_n2982_13878.t61 gnd 0.112993f
C4465 a_n2982_13878.n112 gnd 0.998444f
C4466 a_n2982_13878.n113 gnd 0.299205f
C4467 a_n2982_13878.n114 gnd 0.296972f
C4468 a_n2982_13878.n115 gnd 0.299644f
C4469 a_n2982_13878.n116 gnd 0.293332f
C4470 a_n2982_13878.n117 gnd 0.288167f
C4471 a_n2982_13878.n118 gnd 0.29709f
C4472 a_n2982_13878.n119 gnd 0.299206f
C4473 a_n2982_13878.t34 gnd 1.3603f
C4474 a_n2982_13878.t22 gnd 0.145277f
C4475 a_n2982_13878.t32 gnd 0.145277f
C4476 a_n2982_13878.n120 gnd 1.02333f
C4477 a_n2982_13878.t28 gnd 0.145277f
C4478 a_n2982_13878.t56 gnd 0.145277f
C4479 a_n2982_13878.n121 gnd 1.02333f
C4480 a_n2982_13878.t14 gnd 0.145277f
C4481 a_n2982_13878.t20 gnd 0.145277f
C4482 a_n2982_13878.n122 gnd 1.02333f
C4483 a_n2982_13878.t26 gnd 0.145277f
C4484 a_n2982_13878.t54 gnd 0.145277f
C4485 a_n2982_13878.n123 gnd 1.02333f
C4486 a_n2982_13878.t48 gnd 0.145277f
C4487 a_n2982_13878.t50 gnd 0.145277f
C4488 a_n2982_13878.n124 gnd 1.02333f
C4489 a_n2982_13878.t30 gnd 1.35759f
C4490 a_n2982_13878.n125 gnd 0.994805f
C4491 a_n2982_13878.t77 gnd 0.675756f
C4492 a_n2982_13878.t87 gnd 0.675756f
C4493 a_n2982_13878.t103 gnd 0.675756f
C4494 a_n2982_13878.n126 gnd 0.297105f
C4495 a_n2982_13878.t90 gnd 0.675756f
C4496 a_n2982_13878.t73 gnd 0.675756f
C4497 a_n2982_13878.t74 gnd 0.675756f
C4498 a_n2982_13878.n127 gnd 0.297105f
C4499 a_n2982_13878.t94 gnd 0.675756f
C4500 a_n2982_13878.t83 gnd 0.675756f
C4501 a_n2982_13878.t82 gnd 0.675756f
C4502 a_n2982_13878.n128 gnd 0.297105f
C4503 a_n2982_13878.t86 gnd 0.675756f
C4504 a_n2982_13878.t75 gnd 0.675756f
C4505 a_n2982_13878.t64 gnd 0.675756f
C4506 a_n2982_13878.n129 gnd 0.297105f
C4507 a_n2982_13878.t91 gnd 0.687079f
C4508 a_n2982_13878.n130 gnd 0.293332f
C4509 a_n2982_13878.n131 gnd 0.288005f
C4510 a_n2982_13878.t100 gnd 0.687079f
C4511 a_n2982_13878.n132 gnd 0.293332f
C4512 a_n2982_13878.n133 gnd 0.288005f
C4513 a_n2982_13878.t85 gnd 0.687079f
C4514 a_n2982_13878.n134 gnd 0.293332f
C4515 a_n2982_13878.n135 gnd 0.288005f
C4516 a_n2982_13878.t80 gnd 0.687079f
C4517 a_n2982_13878.n136 gnd 0.293332f
C4518 a_n2982_13878.n137 gnd 0.288005f
C4519 a_n2982_13878.n138 gnd 1.32386f
C4520 a_n2982_13878.t70 gnd 0.675756f
C4521 a_n2982_13878.n139 gnd 0.299205f
C4522 a_n2982_13878.t96 gnd 0.675756f
C4523 a_n2982_13878.n140 gnd 0.296972f
C4524 a_n2982_13878.n141 gnd 0.297105f
C4525 a_n2982_13878.t92 gnd 0.675756f
C4526 a_n2982_13878.n142 gnd 0.293332f
C4527 a_n2982_13878.t65 gnd 0.675756f
C4528 a_n2982_13878.n143 gnd 0.293584f
C4529 a_n2982_13878.n144 gnd 0.299206f
C4530 a_n2982_13878.t67 gnd 0.686627f
C4531 a_n2982_13878.t17 gnd 0.675756f
C4532 a_n2982_13878.n145 gnd 0.299205f
C4533 a_n2982_13878.t11 gnd 0.675756f
C4534 a_n2982_13878.n146 gnd 0.296972f
C4535 a_n2982_13878.n147 gnd 0.297105f
C4536 a_n2982_13878.t15 gnd 0.675756f
C4537 a_n2982_13878.n148 gnd 0.293332f
C4538 a_n2982_13878.t43 gnd 0.675756f
C4539 a_n2982_13878.n149 gnd 0.293584f
C4540 a_n2982_13878.n150 gnd 0.299206f
C4541 a_n2982_13878.t57 gnd 0.686627f
C4542 a_n2982_13878.n151 gnd 1.30834f
C4543 a_n2982_13878.t58 gnd 1.35758f
C4544 a_n2982_13878.t24 gnd 0.145277f
C4545 a_n2982_13878.t38 gnd 0.145277f
C4546 a_n2982_13878.n152 gnd 1.02333f
C4547 a_n2982_13878.t52 gnd 0.145277f
C4548 a_n2982_13878.t44 gnd 0.145277f
C4549 a_n2982_13878.n153 gnd 1.02333f
C4550 a_n2982_13878.t46 gnd 0.145277f
C4551 a_n2982_13878.t16 gnd 0.145277f
C4552 a_n2982_13878.n154 gnd 1.02333f
C4553 a_n2982_13878.n155 gnd 1.02333f
C4554 a_n2982_13878.t12 gnd 0.145277f
C4555 CSoutput.n0 gnd 0.048956f
C4556 CSoutput.t202 gnd 0.323832f
C4557 CSoutput.n1 gnd 0.146226f
C4558 CSoutput.n2 gnd 0.048956f
C4559 CSoutput.t200 gnd 0.323832f
C4560 CSoutput.n3 gnd 0.038801f
C4561 CSoutput.n4 gnd 0.048956f
C4562 CSoutput.t212 gnd 0.323832f
C4563 CSoutput.n5 gnd 0.033459f
C4564 CSoutput.n6 gnd 0.048956f
C4565 CSoutput.t197 gnd 0.323832f
C4566 CSoutput.t207 gnd 0.323832f
C4567 CSoutput.n7 gnd 0.144632f
C4568 CSoutput.n8 gnd 0.048956f
C4569 CSoutput.t210 gnd 0.323832f
C4570 CSoutput.n9 gnd 0.031901f
C4571 CSoutput.n10 gnd 0.048956f
C4572 CSoutput.t193 gnd 0.323832f
C4573 CSoutput.t199 gnd 0.323832f
C4574 CSoutput.n11 gnd 0.144632f
C4575 CSoutput.n12 gnd 0.048956f
C4576 CSoutput.t204 gnd 0.323832f
C4577 CSoutput.n13 gnd 0.033459f
C4578 CSoutput.n14 gnd 0.048956f
C4579 CSoutput.t213 gnd 0.323832f
C4580 CSoutput.t196 gnd 0.323832f
C4581 CSoutput.n15 gnd 0.144632f
C4582 CSoutput.n16 gnd 0.048956f
C4583 CSoutput.t203 gnd 0.323832f
C4584 CSoutput.n17 gnd 0.035736f
C4585 CSoutput.t192 gnd 0.386987f
C4586 CSoutput.t201 gnd 0.323832f
C4587 CSoutput.n18 gnd 0.184639f
C4588 CSoutput.n19 gnd 0.179164f
C4589 CSoutput.n20 gnd 0.207852f
C4590 CSoutput.n21 gnd 0.048956f
C4591 CSoutput.n22 gnd 0.040859f
C4592 CSoutput.n23 gnd 0.144632f
C4593 CSoutput.n24 gnd 0.039387f
C4594 CSoutput.n25 gnd 0.038801f
C4595 CSoutput.n26 gnd 0.048956f
C4596 CSoutput.n27 gnd 0.048956f
C4597 CSoutput.n28 gnd 0.040545f
C4598 CSoutput.n29 gnd 0.034424f
C4599 CSoutput.n30 gnd 0.147852f
C4600 CSoutput.n31 gnd 0.034898f
C4601 CSoutput.n32 gnd 0.048956f
C4602 CSoutput.n33 gnd 0.048956f
C4603 CSoutput.n34 gnd 0.048956f
C4604 CSoutput.n35 gnd 0.040113f
C4605 CSoutput.n36 gnd 0.144632f
C4606 CSoutput.n37 gnd 0.038362f
C4607 CSoutput.n38 gnd 0.039826f
C4608 CSoutput.n39 gnd 0.048956f
C4609 CSoutput.n40 gnd 0.048956f
C4610 CSoutput.n41 gnd 0.040851f
C4611 CSoutput.n42 gnd 0.037338f
C4612 CSoutput.n43 gnd 0.144632f
C4613 CSoutput.n44 gnd 0.038284f
C4614 CSoutput.n45 gnd 0.048956f
C4615 CSoutput.n46 gnd 0.048956f
C4616 CSoutput.n47 gnd 0.048956f
C4617 CSoutput.n48 gnd 0.038284f
C4618 CSoutput.n49 gnd 0.144632f
C4619 CSoutput.n50 gnd 0.037338f
C4620 CSoutput.n51 gnd 0.040851f
C4621 CSoutput.n52 gnd 0.048956f
C4622 CSoutput.n53 gnd 0.048956f
C4623 CSoutput.n54 gnd 0.039826f
C4624 CSoutput.n55 gnd 0.038362f
C4625 CSoutput.n56 gnd 0.144632f
C4626 CSoutput.n57 gnd 0.040113f
C4627 CSoutput.n58 gnd 0.048956f
C4628 CSoutput.n59 gnd 0.048956f
C4629 CSoutput.n60 gnd 0.048956f
C4630 CSoutput.n61 gnd 0.034898f
C4631 CSoutput.n62 gnd 0.147852f
C4632 CSoutput.n63 gnd 0.034424f
C4633 CSoutput.t208 gnd 0.323832f
C4634 CSoutput.n64 gnd 0.144632f
C4635 CSoutput.n65 gnd 0.040545f
C4636 CSoutput.n66 gnd 0.048956f
C4637 CSoutput.n67 gnd 0.048956f
C4638 CSoutput.n68 gnd 0.048956f
C4639 CSoutput.n69 gnd 0.039387f
C4640 CSoutput.n70 gnd 0.144632f
C4641 CSoutput.n71 gnd 0.040859f
C4642 CSoutput.n72 gnd 0.035736f
C4643 CSoutput.n73 gnd 0.048956f
C4644 CSoutput.n74 gnd 0.048956f
C4645 CSoutput.n75 gnd 0.03706f
C4646 CSoutput.n76 gnd 0.02201f
C4647 CSoutput.t194 gnd 0.363848f
C4648 CSoutput.n77 gnd 0.180745f
C4649 CSoutput.n78 gnd 0.739309f
C4650 CSoutput.t181 gnd 0.061065f
C4651 CSoutput.t124 gnd 0.061065f
C4652 CSoutput.n79 gnd 0.472789f
C4653 CSoutput.t102 gnd 0.061065f
C4654 CSoutput.t77 gnd 0.061065f
C4655 CSoutput.n80 gnd 0.471946f
C4656 CSoutput.n81 gnd 0.479024f
C4657 CSoutput.t186 gnd 0.061065f
C4658 CSoutput.t129 gnd 0.061065f
C4659 CSoutput.n82 gnd 0.471946f
C4660 CSoutput.n83 gnd 0.236043f
C4661 CSoutput.t110 gnd 0.061065f
C4662 CSoutput.t112 gnd 0.061065f
C4663 CSoutput.n84 gnd 0.471946f
C4664 CSoutput.n85 gnd 0.236043f
C4665 CSoutput.t172 gnd 0.061065f
C4666 CSoutput.t72 gnd 0.061065f
C4667 CSoutput.n86 gnd 0.471946f
C4668 CSoutput.n87 gnd 0.236043f
C4669 CSoutput.t136 gnd 0.061065f
C4670 CSoutput.t170 gnd 0.061065f
C4671 CSoutput.n88 gnd 0.471946f
C4672 CSoutput.n89 gnd 0.236043f
C4673 CSoutput.t185 gnd 0.061065f
C4674 CSoutput.t79 gnd 0.061065f
C4675 CSoutput.n90 gnd 0.471946f
C4676 CSoutput.n91 gnd 0.236043f
C4677 CSoutput.t159 gnd 0.061065f
C4678 CSoutput.t139 gnd 0.061065f
C4679 CSoutput.n92 gnd 0.471946f
C4680 CSoutput.n93 gnd 0.236043f
C4681 CSoutput.t154 gnd 0.061065f
C4682 CSoutput.t93 gnd 0.061065f
C4683 CSoutput.n94 gnd 0.471946f
C4684 CSoutput.n95 gnd 0.236043f
C4685 CSoutput.t86 gnd 0.061065f
C4686 CSoutput.t73 gnd 0.061065f
C4687 CSoutput.n96 gnd 0.471946f
C4688 CSoutput.n97 gnd 0.432848f
C4689 CSoutput.t173 gnd 0.061065f
C4690 CSoutput.t103 gnd 0.061065f
C4691 CSoutput.n98 gnd 0.472789f
C4692 CSoutput.t145 gnd 0.061065f
C4693 CSoutput.t117 gnd 0.061065f
C4694 CSoutput.n99 gnd 0.471946f
C4695 CSoutput.n100 gnd 0.479024f
C4696 CSoutput.t132 gnd 0.061065f
C4697 CSoutput.t178 gnd 0.061065f
C4698 CSoutput.n101 gnd 0.471946f
C4699 CSoutput.n102 gnd 0.236043f
C4700 CSoutput.t167 gnd 0.061065f
C4701 CSoutput.t191 gnd 0.061065f
C4702 CSoutput.n103 gnd 0.471946f
C4703 CSoutput.n104 gnd 0.236043f
C4704 CSoutput.t130 gnd 0.061065f
C4705 CSoutput.t90 gnd 0.061065f
C4706 CSoutput.n105 gnd 0.471946f
C4707 CSoutput.n106 gnd 0.236043f
C4708 CSoutput.t175 gnd 0.061065f
C4709 CSoutput.t98 gnd 0.061065f
C4710 CSoutput.n107 gnd 0.471946f
C4711 CSoutput.n108 gnd 0.236043f
C4712 CSoutput.t81 gnd 0.061065f
C4713 CSoutput.t182 gnd 0.061065f
C4714 CSoutput.n109 gnd 0.471946f
C4715 CSoutput.n110 gnd 0.236043f
C4716 CSoutput.t116 gnd 0.061065f
C4717 CSoutput.t104 gnd 0.061065f
C4718 CSoutput.n111 gnd 0.471946f
C4719 CSoutput.n112 gnd 0.236043f
C4720 CSoutput.t100 gnd 0.061065f
C4721 CSoutput.t151 gnd 0.061065f
C4722 CSoutput.n113 gnd 0.471946f
C4723 CSoutput.n114 gnd 0.236043f
C4724 CSoutput.t133 gnd 0.061065f
C4725 CSoutput.t125 gnd 0.061065f
C4726 CSoutput.n115 gnd 0.471946f
C4727 CSoutput.n116 gnd 0.351999f
C4728 CSoutput.n117 gnd 0.443869f
C4729 CSoutput.t141 gnd 0.061065f
C4730 CSoutput.t94 gnd 0.061065f
C4731 CSoutput.n118 gnd 0.472789f
C4732 CSoutput.t97 gnd 0.061065f
C4733 CSoutput.t143 gnd 0.061065f
C4734 CSoutput.n119 gnd 0.471946f
C4735 CSoutput.n120 gnd 0.479024f
C4736 CSoutput.t161 gnd 0.061065f
C4737 CSoutput.t89 gnd 0.061065f
C4738 CSoutput.n121 gnd 0.471946f
C4739 CSoutput.n122 gnd 0.236043f
C4740 CSoutput.t120 gnd 0.061065f
C4741 CSoutput.t165 gnd 0.061065f
C4742 CSoutput.n123 gnd 0.471946f
C4743 CSoutput.n124 gnd 0.236043f
C4744 CSoutput.t87 gnd 0.061065f
C4745 CSoutput.t118 gnd 0.061065f
C4746 CSoutput.n125 gnd 0.471946f
C4747 CSoutput.n126 gnd 0.236043f
C4748 CSoutput.t156 gnd 0.061065f
C4749 CSoutput.t101 gnd 0.061065f
C4750 CSoutput.n127 gnd 0.471946f
C4751 CSoutput.n128 gnd 0.236043f
C4752 CSoutput.t140 gnd 0.061065f
C4753 CSoutput.t85 gnd 0.061065f
C4754 CSoutput.n129 gnd 0.471946f
C4755 CSoutput.n130 gnd 0.236043f
C4756 CSoutput.t142 gnd 0.061065f
C4757 CSoutput.t95 gnd 0.061065f
C4758 CSoutput.n131 gnd 0.471946f
C4759 CSoutput.n132 gnd 0.236043f
C4760 CSoutput.t88 gnd 0.061065f
C4761 CSoutput.t148 gnd 0.061065f
C4762 CSoutput.n133 gnd 0.471946f
C4763 CSoutput.n134 gnd 0.236043f
C4764 CSoutput.t162 gnd 0.061065f
C4765 CSoutput.t160 gnd 0.061065f
C4766 CSoutput.n135 gnd 0.471946f
C4767 CSoutput.n136 gnd 0.351999f
C4768 CSoutput.n137 gnd 0.496132f
C4769 CSoutput.n138 gnd 9.50409f
C4770 CSoutput.n140 gnd 0.866018f
C4771 CSoutput.n141 gnd 0.649514f
C4772 CSoutput.n142 gnd 0.866018f
C4773 CSoutput.n143 gnd 0.866018f
C4774 CSoutput.n144 gnd 2.33159f
C4775 CSoutput.n145 gnd 0.866018f
C4776 CSoutput.n146 gnd 0.866018f
C4777 CSoutput.t209 gnd 1.08252f
C4778 CSoutput.n147 gnd 0.866018f
C4779 CSoutput.n148 gnd 0.866018f
C4780 CSoutput.n152 gnd 0.866018f
C4781 CSoutput.n156 gnd 0.866018f
C4782 CSoutput.n157 gnd 0.866018f
C4783 CSoutput.n159 gnd 0.866018f
C4784 CSoutput.n164 gnd 0.866018f
C4785 CSoutput.n166 gnd 0.866018f
C4786 CSoutput.n167 gnd 0.866018f
C4787 CSoutput.n169 gnd 0.866018f
C4788 CSoutput.n170 gnd 0.866018f
C4789 CSoutput.n172 gnd 0.866018f
C4790 CSoutput.t195 gnd 14.471099f
C4791 CSoutput.n174 gnd 0.866018f
C4792 CSoutput.n175 gnd 0.649514f
C4793 CSoutput.n176 gnd 0.866018f
C4794 CSoutput.n177 gnd 0.866018f
C4795 CSoutput.n178 gnd 2.33159f
C4796 CSoutput.n179 gnd 0.866018f
C4797 CSoutput.n180 gnd 0.866018f
C4798 CSoutput.t198 gnd 1.08252f
C4799 CSoutput.n181 gnd 0.866018f
C4800 CSoutput.n182 gnd 0.866018f
C4801 CSoutput.n186 gnd 0.866018f
C4802 CSoutput.n190 gnd 0.866018f
C4803 CSoutput.n191 gnd 0.866018f
C4804 CSoutput.n193 gnd 0.866018f
C4805 CSoutput.n198 gnd 0.866018f
C4806 CSoutput.n200 gnd 0.866018f
C4807 CSoutput.n201 gnd 0.866018f
C4808 CSoutput.n203 gnd 0.866018f
C4809 CSoutput.n204 gnd 0.866018f
C4810 CSoutput.n206 gnd 0.866018f
C4811 CSoutput.n207 gnd 0.649514f
C4812 CSoutput.n209 gnd 0.866018f
C4813 CSoutput.n210 gnd 0.649514f
C4814 CSoutput.n211 gnd 0.866018f
C4815 CSoutput.n212 gnd 0.866018f
C4816 CSoutput.n213 gnd 2.33159f
C4817 CSoutput.n214 gnd 0.866018f
C4818 CSoutput.n215 gnd 0.866018f
C4819 CSoutput.t206 gnd 1.08252f
C4820 CSoutput.n216 gnd 0.866018f
C4821 CSoutput.n217 gnd 2.33159f
C4822 CSoutput.n219 gnd 0.866018f
C4823 CSoutput.n220 gnd 0.866018f
C4824 CSoutput.n222 gnd 0.866018f
C4825 CSoutput.n223 gnd 0.866018f
C4826 CSoutput.t211 gnd 14.2352f
C4827 CSoutput.t205 gnd 14.471099f
C4828 CSoutput.n229 gnd 2.71683f
C4829 CSoutput.n230 gnd 11.0674f
C4830 CSoutput.n231 gnd 11.5305f
C4831 CSoutput.n236 gnd 2.94305f
C4832 CSoutput.n242 gnd 0.866018f
C4833 CSoutput.n244 gnd 0.866018f
C4834 CSoutput.n246 gnd 0.866018f
C4835 CSoutput.n248 gnd 0.866018f
C4836 CSoutput.n250 gnd 0.866018f
C4837 CSoutput.n256 gnd 0.866018f
C4838 CSoutput.n263 gnd 1.58881f
C4839 CSoutput.n264 gnd 1.58881f
C4840 CSoutput.n265 gnd 0.866018f
C4841 CSoutput.n266 gnd 0.866018f
C4842 CSoutput.n268 gnd 0.649514f
C4843 CSoutput.n269 gnd 0.55625f
C4844 CSoutput.n271 gnd 0.649514f
C4845 CSoutput.n272 gnd 0.55625f
C4846 CSoutput.n273 gnd 0.649514f
C4847 CSoutput.n275 gnd 0.866018f
C4848 CSoutput.n277 gnd 2.33159f
C4849 CSoutput.n278 gnd 2.71683f
C4850 CSoutput.n279 gnd 10.1791f
C4851 CSoutput.n281 gnd 0.649514f
C4852 CSoutput.n282 gnd 1.67124f
C4853 CSoutput.n283 gnd 0.649514f
C4854 CSoutput.n285 gnd 0.866018f
C4855 CSoutput.n287 gnd 2.33159f
C4856 CSoutput.n288 gnd 5.07803f
C4857 CSoutput.t123 gnd 0.061065f
C4858 CSoutput.t135 gnd 0.061065f
C4859 CSoutput.n289 gnd 0.472789f
C4860 CSoutput.t76 gnd 0.061065f
C4861 CSoutput.t189 gnd 0.061065f
C4862 CSoutput.n290 gnd 0.471946f
C4863 CSoutput.n291 gnd 0.479024f
C4864 CSoutput.t183 gnd 0.061065f
C4865 CSoutput.t163 gnd 0.061065f
C4866 CSoutput.n292 gnd 0.471946f
C4867 CSoutput.n293 gnd 0.236043f
C4868 CSoutput.t92 gnd 0.061065f
C4869 CSoutput.t96 gnd 0.061065f
C4870 CSoutput.n294 gnd 0.471946f
C4871 CSoutput.n295 gnd 0.236043f
C4872 CSoutput.t82 gnd 0.061065f
C4873 CSoutput.t134 gnd 0.061065f
C4874 CSoutput.n296 gnd 0.471946f
C4875 CSoutput.n297 gnd 0.236043f
C4876 CSoutput.t169 gnd 0.061065f
C4877 CSoutput.t174 gnd 0.061065f
C4878 CSoutput.n298 gnd 0.471946f
C4879 CSoutput.n299 gnd 0.236043f
C4880 CSoutput.t78 gnd 0.061065f
C4881 CSoutput.t184 gnd 0.061065f
C4882 CSoutput.n300 gnd 0.471946f
C4883 CSoutput.n301 gnd 0.236043f
C4884 CSoutput.t138 gnd 0.061065f
C4885 CSoutput.t114 gnd 0.061065f
C4886 CSoutput.n302 gnd 0.471946f
C4887 CSoutput.n303 gnd 0.236043f
C4888 CSoutput.t99 gnd 0.061065f
C4889 CSoutput.t109 gnd 0.061065f
C4890 CSoutput.n304 gnd 0.471946f
C4891 CSoutput.n305 gnd 0.236043f
C4892 CSoutput.t83 gnd 0.061065f
C4893 CSoutput.t84 gnd 0.061065f
C4894 CSoutput.n306 gnd 0.471946f
C4895 CSoutput.n307 gnd 0.432848f
C4896 CSoutput.t153 gnd 0.061065f
C4897 CSoutput.t80 gnd 0.061065f
C4898 CSoutput.n308 gnd 0.472789f
C4899 CSoutput.t179 gnd 0.061065f
C4900 CSoutput.t171 gnd 0.061065f
C4901 CSoutput.n309 gnd 0.471946f
C4902 CSoutput.n310 gnd 0.479024f
C4903 CSoutput.t108 gnd 0.061065f
C4904 CSoutput.t166 gnd 0.061065f
C4905 CSoutput.n311 gnd 0.471946f
C4906 CSoutput.n312 gnd 0.236043f
C4907 CSoutput.t119 gnd 0.061065f
C4908 CSoutput.t168 gnd 0.061065f
C4909 CSoutput.n313 gnd 0.471946f
C4910 CSoutput.n314 gnd 0.236043f
C4911 CSoutput.t147 gnd 0.061065f
C4912 CSoutput.t176 gnd 0.061065f
C4913 CSoutput.n315 gnd 0.471946f
C4914 CSoutput.n316 gnd 0.236043f
C4915 CSoutput.t131 gnd 0.061065f
C4916 CSoutput.t180 gnd 0.061065f
C4917 CSoutput.n317 gnd 0.471946f
C4918 CSoutput.n318 gnd 0.236043f
C4919 CSoutput.t128 gnd 0.061065f
C4920 CSoutput.t113 gnd 0.061065f
C4921 CSoutput.n319 gnd 0.471946f
C4922 CSoutput.n320 gnd 0.236043f
C4923 CSoutput.t152 gnd 0.061065f
C4924 CSoutput.t190 gnd 0.061065f
C4925 CSoutput.n321 gnd 0.471946f
C4926 CSoutput.n322 gnd 0.236043f
C4927 CSoutput.t127 gnd 0.061065f
C4928 CSoutput.t107 gnd 0.061065f
C4929 CSoutput.n323 gnd 0.471946f
C4930 CSoutput.n324 gnd 0.236043f
C4931 CSoutput.t158 gnd 0.061065f
C4932 CSoutput.t122 gnd 0.061065f
C4933 CSoutput.n325 gnd 0.471946f
C4934 CSoutput.n326 gnd 0.351999f
C4935 CSoutput.n327 gnd 0.443869f
C4936 CSoutput.t149 gnd 0.061065f
C4937 CSoutput.t137 gnd 0.061065f
C4938 CSoutput.n328 gnd 0.472789f
C4939 CSoutput.t126 gnd 0.061065f
C4940 CSoutput.t106 gnd 0.061065f
C4941 CSoutput.n329 gnd 0.471946f
C4942 CSoutput.n330 gnd 0.479024f
C4943 CSoutput.t75 gnd 0.061065f
C4944 CSoutput.t164 gnd 0.061065f
C4945 CSoutput.n331 gnd 0.471946f
C4946 CSoutput.n332 gnd 0.236043f
C4947 CSoutput.t115 gnd 0.061065f
C4948 CSoutput.t105 gnd 0.061065f
C4949 CSoutput.n333 gnd 0.471946f
C4950 CSoutput.n334 gnd 0.236043f
C4951 CSoutput.t146 gnd 0.061065f
C4952 CSoutput.t157 gnd 0.061065f
C4953 CSoutput.n335 gnd 0.471946f
C4954 CSoutput.n336 gnd 0.236043f
C4955 CSoutput.t91 gnd 0.061065f
C4956 CSoutput.t188 gnd 0.061065f
C4957 CSoutput.n337 gnd 0.471946f
C4958 CSoutput.n338 gnd 0.236043f
C4959 CSoutput.t155 gnd 0.061065f
C4960 CSoutput.t144 gnd 0.061065f
C4961 CSoutput.n339 gnd 0.471946f
C4962 CSoutput.n340 gnd 0.236043f
C4963 CSoutput.t150 gnd 0.061065f
C4964 CSoutput.t187 gnd 0.061065f
C4965 CSoutput.n341 gnd 0.471946f
C4966 CSoutput.n342 gnd 0.236043f
C4967 CSoutput.t111 gnd 0.061065f
C4968 CSoutput.t74 gnd 0.061065f
C4969 CSoutput.n343 gnd 0.471946f
C4970 CSoutput.n344 gnd 0.236043f
C4971 CSoutput.t121 gnd 0.061065f
C4972 CSoutput.t177 gnd 0.061065f
C4973 CSoutput.n345 gnd 0.471944f
C4974 CSoutput.n346 gnd 0.352001f
C4975 CSoutput.n347 gnd 0.496132f
C4976 CSoutput.n348 gnd 13.661f
C4977 CSoutput.t30 gnd 0.053432f
C4978 CSoutput.t68 gnd 0.053432f
C4979 CSoutput.n349 gnd 0.473726f
C4980 CSoutput.t24 gnd 0.053432f
C4981 CSoutput.t29 gnd 0.053432f
C4982 CSoutput.n350 gnd 0.472146f
C4983 CSoutput.n351 gnd 0.439952f
C4984 CSoutput.t18 gnd 0.053432f
C4985 CSoutput.t33 gnd 0.053432f
C4986 CSoutput.n352 gnd 0.472146f
C4987 CSoutput.n353 gnd 0.216875f
C4988 CSoutput.t42 gnd 0.053432f
C4989 CSoutput.t25 gnd 0.053432f
C4990 CSoutput.n354 gnd 0.472146f
C4991 CSoutput.n355 gnd 0.216875f
C4992 CSoutput.t32 gnd 0.053432f
C4993 CSoutput.t61 gnd 0.053432f
C4994 CSoutput.n356 gnd 0.472146f
C4995 CSoutput.n357 gnd 0.216875f
C4996 CSoutput.t39 gnd 0.053432f
C4997 CSoutput.t46 gnd 0.053432f
C4998 CSoutput.n358 gnd 0.472146f
C4999 CSoutput.n359 gnd 0.400015f
C5000 CSoutput.t65 gnd 0.053432f
C5001 CSoutput.t0 gnd 0.053432f
C5002 CSoutput.n360 gnd 0.473726f
C5003 CSoutput.t9 gnd 0.053432f
C5004 CSoutput.t59 gnd 0.053432f
C5005 CSoutput.n361 gnd 0.472146f
C5006 CSoutput.n362 gnd 0.439952f
C5007 CSoutput.t2 gnd 0.053432f
C5008 CSoutput.t54 gnd 0.053432f
C5009 CSoutput.n363 gnd 0.472146f
C5010 CSoutput.n364 gnd 0.216875f
C5011 CSoutput.t60 gnd 0.053432f
C5012 CSoutput.t1 gnd 0.053432f
C5013 CSoutput.n365 gnd 0.472146f
C5014 CSoutput.n366 gnd 0.216875f
C5015 CSoutput.t48 gnd 0.053432f
C5016 CSoutput.t36 gnd 0.053432f
C5017 CSoutput.n367 gnd 0.472146f
C5018 CSoutput.n368 gnd 0.216875f
C5019 CSoutput.t3 gnd 0.053432f
C5020 CSoutput.t49 gnd 0.053432f
C5021 CSoutput.n369 gnd 0.472146f
C5022 CSoutput.n370 gnd 0.329263f
C5023 CSoutput.n371 gnd 0.415304f
C5024 CSoutput.t10 gnd 0.053432f
C5025 CSoutput.t62 gnd 0.053432f
C5026 CSoutput.n372 gnd 0.473726f
C5027 CSoutput.t23 gnd 0.053432f
C5028 CSoutput.t26 gnd 0.053432f
C5029 CSoutput.n373 gnd 0.472146f
C5030 CSoutput.n374 gnd 0.439952f
C5031 CSoutput.t4 gnd 0.053432f
C5032 CSoutput.t51 gnd 0.053432f
C5033 CSoutput.n375 gnd 0.472146f
C5034 CSoutput.n376 gnd 0.216875f
C5035 CSoutput.t31 gnd 0.053432f
C5036 CSoutput.t11 gnd 0.053432f
C5037 CSoutput.n377 gnd 0.472146f
C5038 CSoutput.n378 gnd 0.216875f
C5039 CSoutput.t16 gnd 0.053432f
C5040 CSoutput.t71 gnd 0.053432f
C5041 CSoutput.n379 gnd 0.472146f
C5042 CSoutput.n380 gnd 0.216875f
C5043 CSoutput.t17 gnd 0.053432f
C5044 CSoutput.t21 gnd 0.053432f
C5045 CSoutput.n381 gnd 0.472146f
C5046 CSoutput.n382 gnd 0.329263f
C5047 CSoutput.n383 gnd 0.445971f
C5048 CSoutput.n384 gnd 13.269501f
C5049 CSoutput.t20 gnd 0.053432f
C5050 CSoutput.t50 gnd 0.053432f
C5051 CSoutput.n385 gnd 0.473726f
C5052 CSoutput.t47 gnd 0.053432f
C5053 CSoutput.t35 gnd 0.053432f
C5054 CSoutput.n386 gnd 0.472146f
C5055 CSoutput.n387 gnd 0.439952f
C5056 CSoutput.t53 gnd 0.053432f
C5057 CSoutput.t27 gnd 0.053432f
C5058 CSoutput.n388 gnd 0.472146f
C5059 CSoutput.n389 gnd 0.216875f
C5060 CSoutput.t40 gnd 0.053432f
C5061 CSoutput.t63 gnd 0.053432f
C5062 CSoutput.n390 gnd 0.472146f
C5063 CSoutput.n391 gnd 0.216875f
C5064 CSoutput.t15 gnd 0.053432f
C5065 CSoutput.t52 gnd 0.053432f
C5066 CSoutput.n392 gnd 0.472146f
C5067 CSoutput.n393 gnd 0.216875f
C5068 CSoutput.t8 gnd 0.053432f
C5069 CSoutput.t55 gnd 0.053432f
C5070 CSoutput.n394 gnd 0.472146f
C5071 CSoutput.n395 gnd 0.400015f
C5072 CSoutput.t12 gnd 0.053432f
C5073 CSoutput.t7 gnd 0.053432f
C5074 CSoutput.n396 gnd 0.473726f
C5075 CSoutput.t5 gnd 0.053432f
C5076 CSoutput.t69 gnd 0.053432f
C5077 CSoutput.n397 gnd 0.472146f
C5078 CSoutput.n398 gnd 0.439952f
C5079 CSoutput.t70 gnd 0.053432f
C5080 CSoutput.t13 gnd 0.053432f
C5081 CSoutput.n399 gnd 0.472146f
C5082 CSoutput.n400 gnd 0.216875f
C5083 CSoutput.t14 gnd 0.053432f
C5084 CSoutput.t45 gnd 0.053432f
C5085 CSoutput.n401 gnd 0.472146f
C5086 CSoutput.n402 gnd 0.216875f
C5087 CSoutput.t44 gnd 0.053432f
C5088 CSoutput.t64 gnd 0.053432f
C5089 CSoutput.n403 gnd 0.472146f
C5090 CSoutput.n404 gnd 0.216875f
C5091 CSoutput.t67 gnd 0.053432f
C5092 CSoutput.t58 gnd 0.053432f
C5093 CSoutput.n405 gnd 0.472146f
C5094 CSoutput.n406 gnd 0.329263f
C5095 CSoutput.n407 gnd 0.415304f
C5096 CSoutput.t38 gnd 0.053432f
C5097 CSoutput.t56 gnd 0.053432f
C5098 CSoutput.n408 gnd 0.473726f
C5099 CSoutput.t19 gnd 0.053432f
C5100 CSoutput.t28 gnd 0.053432f
C5101 CSoutput.n409 gnd 0.472146f
C5102 CSoutput.n410 gnd 0.439952f
C5103 CSoutput.t34 gnd 0.053432f
C5104 CSoutput.t43 gnd 0.053432f
C5105 CSoutput.n411 gnd 0.472146f
C5106 CSoutput.n412 gnd 0.216875f
C5107 CSoutput.t57 gnd 0.053432f
C5108 CSoutput.t37 gnd 0.053432f
C5109 CSoutput.n413 gnd 0.472146f
C5110 CSoutput.n414 gnd 0.216875f
C5111 CSoutput.t41 gnd 0.053432f
C5112 CSoutput.t66 gnd 0.053432f
C5113 CSoutput.n415 gnd 0.472146f
C5114 CSoutput.n416 gnd 0.216875f
C5115 CSoutput.t6 gnd 0.053432f
C5116 CSoutput.t22 gnd 0.053432f
C5117 CSoutput.n417 gnd 0.472146f
C5118 CSoutput.n418 gnd 0.329263f
C5119 CSoutput.n419 gnd 0.445971f
C5120 CSoutput.n420 gnd 7.88743f
C5121 CSoutput.n421 gnd 14.775301f
C5122 commonsourceibias.n0 gnd 0.01231f
C5123 commonsourceibias.t89 gnd 0.186396f
C5124 commonsourceibias.t51 gnd 0.17235f
C5125 commonsourceibias.n1 gnd 0.068768f
C5126 commonsourceibias.n2 gnd 0.009225f
C5127 commonsourceibias.t95 gnd 0.17235f
C5128 commonsourceibias.n3 gnd 0.007462f
C5129 commonsourceibias.n4 gnd 0.009225f
C5130 commonsourceibias.t90 gnd 0.17235f
C5131 commonsourceibias.n5 gnd 0.008906f
C5132 commonsourceibias.n6 gnd 0.009225f
C5133 commonsourceibias.t101 gnd 0.17235f
C5134 commonsourceibias.n7 gnd 0.068768f
C5135 commonsourceibias.t86 gnd 0.17235f
C5136 commonsourceibias.n8 gnd 0.007451f
C5137 commonsourceibias.n9 gnd 0.01231f
C5138 commonsourceibias.t8 gnd 0.186396f
C5139 commonsourceibias.t38 gnd 0.17235f
C5140 commonsourceibias.n10 gnd 0.068768f
C5141 commonsourceibias.n11 gnd 0.009225f
C5142 commonsourceibias.t0 gnd 0.17235f
C5143 commonsourceibias.n12 gnd 0.007462f
C5144 commonsourceibias.n13 gnd 0.009225f
C5145 commonsourceibias.t6 gnd 0.17235f
C5146 commonsourceibias.n14 gnd 0.008906f
C5147 commonsourceibias.n15 gnd 0.009225f
C5148 commonsourceibias.t44 gnd 0.17235f
C5149 commonsourceibias.n16 gnd 0.068768f
C5150 commonsourceibias.t12 gnd 0.17235f
C5151 commonsourceibias.n17 gnd 0.007451f
C5152 commonsourceibias.n18 gnd 0.009225f
C5153 commonsourceibias.t20 gnd 0.17235f
C5154 commonsourceibias.t2 gnd 0.17235f
C5155 commonsourceibias.n19 gnd 0.068768f
C5156 commonsourceibias.n20 gnd 0.009225f
C5157 commonsourceibias.t10 gnd 0.17235f
C5158 commonsourceibias.n21 gnd 0.068768f
C5159 commonsourceibias.n22 gnd 0.009225f
C5160 commonsourceibias.t34 gnd 0.17235f
C5161 commonsourceibias.n23 gnd 0.068768f
C5162 commonsourceibias.n24 gnd 0.046441f
C5163 commonsourceibias.t16 gnd 0.17235f
C5164 commonsourceibias.t22 gnd 0.194477f
C5165 commonsourceibias.n25 gnd 0.079804f
C5166 commonsourceibias.n26 gnd 0.082619f
C5167 commonsourceibias.n27 gnd 0.01137f
C5168 commonsourceibias.n28 gnd 0.012578f
C5169 commonsourceibias.n29 gnd 0.009225f
C5170 commonsourceibias.n30 gnd 0.009225f
C5171 commonsourceibias.n31 gnd 0.012496f
C5172 commonsourceibias.n32 gnd 0.007462f
C5173 commonsourceibias.n33 gnd 0.012651f
C5174 commonsourceibias.n34 gnd 0.009225f
C5175 commonsourceibias.n35 gnd 0.009225f
C5176 commonsourceibias.n36 gnd 0.012728f
C5177 commonsourceibias.n37 gnd 0.010975f
C5178 commonsourceibias.n38 gnd 0.008906f
C5179 commonsourceibias.n39 gnd 0.009225f
C5180 commonsourceibias.n40 gnd 0.009225f
C5181 commonsourceibias.n41 gnd 0.011283f
C5182 commonsourceibias.n42 gnd 0.012665f
C5183 commonsourceibias.n43 gnd 0.068768f
C5184 commonsourceibias.n44 gnd 0.01258f
C5185 commonsourceibias.n45 gnd 0.009225f
C5186 commonsourceibias.n46 gnd 0.009225f
C5187 commonsourceibias.n47 gnd 0.009225f
C5188 commonsourceibias.n48 gnd 0.01258f
C5189 commonsourceibias.n49 gnd 0.068768f
C5190 commonsourceibias.n50 gnd 0.012665f
C5191 commonsourceibias.n51 gnd 0.011283f
C5192 commonsourceibias.n52 gnd 0.009225f
C5193 commonsourceibias.n53 gnd 0.009225f
C5194 commonsourceibias.n54 gnd 0.009225f
C5195 commonsourceibias.n55 gnd 0.010975f
C5196 commonsourceibias.n56 gnd 0.012728f
C5197 commonsourceibias.n57 gnd 0.068768f
C5198 commonsourceibias.n58 gnd 0.012651f
C5199 commonsourceibias.n59 gnd 0.009225f
C5200 commonsourceibias.n60 gnd 0.009225f
C5201 commonsourceibias.n61 gnd 0.009225f
C5202 commonsourceibias.n62 gnd 0.012496f
C5203 commonsourceibias.n63 gnd 0.068768f
C5204 commonsourceibias.n64 gnd 0.012578f
C5205 commonsourceibias.n65 gnd 0.01137f
C5206 commonsourceibias.n66 gnd 0.009225f
C5207 commonsourceibias.n67 gnd 0.009225f
C5208 commonsourceibias.n68 gnd 0.009358f
C5209 commonsourceibias.n69 gnd 0.009674f
C5210 commonsourceibias.n70 gnd 0.082281f
C5211 commonsourceibias.n71 gnd 0.091278f
C5212 commonsourceibias.t9 gnd 0.019906f
C5213 commonsourceibias.t39 gnd 0.019906f
C5214 commonsourceibias.n72 gnd 0.1759f
C5215 commonsourceibias.n73 gnd 0.151991f
C5216 commonsourceibias.t1 gnd 0.019906f
C5217 commonsourceibias.t7 gnd 0.019906f
C5218 commonsourceibias.n74 gnd 0.1759f
C5219 commonsourceibias.n75 gnd 0.080798f
C5220 commonsourceibias.t45 gnd 0.019906f
C5221 commonsourceibias.t13 gnd 0.019906f
C5222 commonsourceibias.n76 gnd 0.1759f
C5223 commonsourceibias.n77 gnd 0.067503f
C5224 commonsourceibias.t17 gnd 0.019906f
C5225 commonsourceibias.t23 gnd 0.019906f
C5226 commonsourceibias.n78 gnd 0.176489f
C5227 commonsourceibias.t11 gnd 0.019906f
C5228 commonsourceibias.t35 gnd 0.019906f
C5229 commonsourceibias.n79 gnd 0.1759f
C5230 commonsourceibias.n80 gnd 0.163906f
C5231 commonsourceibias.t21 gnd 0.019906f
C5232 commonsourceibias.t3 gnd 0.019906f
C5233 commonsourceibias.n81 gnd 0.1759f
C5234 commonsourceibias.n82 gnd 0.067503f
C5235 commonsourceibias.n83 gnd 0.081739f
C5236 commonsourceibias.n84 gnd 0.009225f
C5237 commonsourceibias.t77 gnd 0.17235f
C5238 commonsourceibias.t94 gnd 0.17235f
C5239 commonsourceibias.n85 gnd 0.068768f
C5240 commonsourceibias.n86 gnd 0.009225f
C5241 commonsourceibias.t87 gnd 0.17235f
C5242 commonsourceibias.n87 gnd 0.068768f
C5243 commonsourceibias.n88 gnd 0.009225f
C5244 commonsourceibias.t58 gnd 0.17235f
C5245 commonsourceibias.n89 gnd 0.068768f
C5246 commonsourceibias.n90 gnd 0.046441f
C5247 commonsourceibias.t80 gnd 0.17235f
C5248 commonsourceibias.t73 gnd 0.194477f
C5249 commonsourceibias.n91 gnd 0.079804f
C5250 commonsourceibias.n92 gnd 0.082619f
C5251 commonsourceibias.n93 gnd 0.01137f
C5252 commonsourceibias.n94 gnd 0.012578f
C5253 commonsourceibias.n95 gnd 0.009225f
C5254 commonsourceibias.n96 gnd 0.009225f
C5255 commonsourceibias.n97 gnd 0.012496f
C5256 commonsourceibias.n98 gnd 0.007462f
C5257 commonsourceibias.n99 gnd 0.012651f
C5258 commonsourceibias.n100 gnd 0.009225f
C5259 commonsourceibias.n101 gnd 0.009225f
C5260 commonsourceibias.n102 gnd 0.012728f
C5261 commonsourceibias.n103 gnd 0.010975f
C5262 commonsourceibias.n104 gnd 0.008906f
C5263 commonsourceibias.n105 gnd 0.009225f
C5264 commonsourceibias.n106 gnd 0.009225f
C5265 commonsourceibias.n107 gnd 0.011283f
C5266 commonsourceibias.n108 gnd 0.012665f
C5267 commonsourceibias.n109 gnd 0.068768f
C5268 commonsourceibias.n110 gnd 0.01258f
C5269 commonsourceibias.n111 gnd 0.009181f
C5270 commonsourceibias.n112 gnd 0.066685f
C5271 commonsourceibias.n113 gnd 0.009181f
C5272 commonsourceibias.n114 gnd 0.01258f
C5273 commonsourceibias.n115 gnd 0.068768f
C5274 commonsourceibias.n116 gnd 0.012665f
C5275 commonsourceibias.n117 gnd 0.011283f
C5276 commonsourceibias.n118 gnd 0.009225f
C5277 commonsourceibias.n119 gnd 0.009225f
C5278 commonsourceibias.n120 gnd 0.009225f
C5279 commonsourceibias.n121 gnd 0.010975f
C5280 commonsourceibias.n122 gnd 0.012728f
C5281 commonsourceibias.n123 gnd 0.068768f
C5282 commonsourceibias.n124 gnd 0.012651f
C5283 commonsourceibias.n125 gnd 0.009225f
C5284 commonsourceibias.n126 gnd 0.009225f
C5285 commonsourceibias.n127 gnd 0.009225f
C5286 commonsourceibias.n128 gnd 0.012496f
C5287 commonsourceibias.n129 gnd 0.068768f
C5288 commonsourceibias.n130 gnd 0.012578f
C5289 commonsourceibias.n131 gnd 0.01137f
C5290 commonsourceibias.n132 gnd 0.009225f
C5291 commonsourceibias.n133 gnd 0.009225f
C5292 commonsourceibias.n134 gnd 0.009358f
C5293 commonsourceibias.n135 gnd 0.009674f
C5294 commonsourceibias.n136 gnd 0.082281f
C5295 commonsourceibias.n137 gnd 0.053268f
C5296 commonsourceibias.n138 gnd 0.01231f
C5297 commonsourceibias.t54 gnd 0.186396f
C5298 commonsourceibias.t119 gnd 0.17235f
C5299 commonsourceibias.n139 gnd 0.068768f
C5300 commonsourceibias.n140 gnd 0.009225f
C5301 commonsourceibias.t110 gnd 0.17235f
C5302 commonsourceibias.n141 gnd 0.007462f
C5303 commonsourceibias.n142 gnd 0.009225f
C5304 commonsourceibias.t60 gnd 0.17235f
C5305 commonsourceibias.n143 gnd 0.008906f
C5306 commonsourceibias.n144 gnd 0.009225f
C5307 commonsourceibias.t117 gnd 0.17235f
C5308 commonsourceibias.n145 gnd 0.068768f
C5309 commonsourceibias.t65 gnd 0.17235f
C5310 commonsourceibias.n146 gnd 0.007451f
C5311 commonsourceibias.n147 gnd 0.009225f
C5312 commonsourceibias.t59 gnd 0.17235f
C5313 commonsourceibias.t118 gnd 0.17235f
C5314 commonsourceibias.n148 gnd 0.068768f
C5315 commonsourceibias.n149 gnd 0.009225f
C5316 commonsourceibias.t71 gnd 0.17235f
C5317 commonsourceibias.n150 gnd 0.068768f
C5318 commonsourceibias.n151 gnd 0.009225f
C5319 commonsourceibias.t83 gnd 0.17235f
C5320 commonsourceibias.n152 gnd 0.068768f
C5321 commonsourceibias.n153 gnd 0.046441f
C5322 commonsourceibias.t116 gnd 0.17235f
C5323 commonsourceibias.t70 gnd 0.194477f
C5324 commonsourceibias.n154 gnd 0.079804f
C5325 commonsourceibias.n155 gnd 0.082619f
C5326 commonsourceibias.n156 gnd 0.01137f
C5327 commonsourceibias.n157 gnd 0.012578f
C5328 commonsourceibias.n158 gnd 0.009225f
C5329 commonsourceibias.n159 gnd 0.009225f
C5330 commonsourceibias.n160 gnd 0.012496f
C5331 commonsourceibias.n161 gnd 0.007462f
C5332 commonsourceibias.n162 gnd 0.012651f
C5333 commonsourceibias.n163 gnd 0.009225f
C5334 commonsourceibias.n164 gnd 0.009225f
C5335 commonsourceibias.n165 gnd 0.012728f
C5336 commonsourceibias.n166 gnd 0.010975f
C5337 commonsourceibias.n167 gnd 0.008906f
C5338 commonsourceibias.n168 gnd 0.009225f
C5339 commonsourceibias.n169 gnd 0.009225f
C5340 commonsourceibias.n170 gnd 0.011283f
C5341 commonsourceibias.n171 gnd 0.012665f
C5342 commonsourceibias.n172 gnd 0.068768f
C5343 commonsourceibias.n173 gnd 0.01258f
C5344 commonsourceibias.n174 gnd 0.009225f
C5345 commonsourceibias.n175 gnd 0.009225f
C5346 commonsourceibias.n176 gnd 0.009225f
C5347 commonsourceibias.n177 gnd 0.01258f
C5348 commonsourceibias.n178 gnd 0.068768f
C5349 commonsourceibias.n179 gnd 0.012665f
C5350 commonsourceibias.n180 gnd 0.011283f
C5351 commonsourceibias.n181 gnd 0.009225f
C5352 commonsourceibias.n182 gnd 0.009225f
C5353 commonsourceibias.n183 gnd 0.009225f
C5354 commonsourceibias.n184 gnd 0.010975f
C5355 commonsourceibias.n185 gnd 0.012728f
C5356 commonsourceibias.n186 gnd 0.068768f
C5357 commonsourceibias.n187 gnd 0.012651f
C5358 commonsourceibias.n188 gnd 0.009225f
C5359 commonsourceibias.n189 gnd 0.009225f
C5360 commonsourceibias.n190 gnd 0.009225f
C5361 commonsourceibias.n191 gnd 0.012496f
C5362 commonsourceibias.n192 gnd 0.068768f
C5363 commonsourceibias.n193 gnd 0.012578f
C5364 commonsourceibias.n194 gnd 0.01137f
C5365 commonsourceibias.n195 gnd 0.009225f
C5366 commonsourceibias.n196 gnd 0.009225f
C5367 commonsourceibias.n197 gnd 0.009358f
C5368 commonsourceibias.n198 gnd 0.009674f
C5369 commonsourceibias.n199 gnd 0.082281f
C5370 commonsourceibias.n200 gnd 0.028001f
C5371 commonsourceibias.n201 gnd 0.147196f
C5372 commonsourceibias.n202 gnd 0.01231f
C5373 commonsourceibias.t57 gnd 0.17235f
C5374 commonsourceibias.n203 gnd 0.068768f
C5375 commonsourceibias.n204 gnd 0.009225f
C5376 commonsourceibias.t96 gnd 0.17235f
C5377 commonsourceibias.n205 gnd 0.007462f
C5378 commonsourceibias.n206 gnd 0.009225f
C5379 commonsourceibias.t93 gnd 0.17235f
C5380 commonsourceibias.n207 gnd 0.008906f
C5381 commonsourceibias.n208 gnd 0.009225f
C5382 commonsourceibias.t115 gnd 0.17235f
C5383 commonsourceibias.n209 gnd 0.068768f
C5384 commonsourceibias.t68 gnd 0.17235f
C5385 commonsourceibias.n210 gnd 0.007451f
C5386 commonsourceibias.n211 gnd 0.009225f
C5387 commonsourceibias.t88 gnd 0.17235f
C5388 commonsourceibias.t108 gnd 0.17235f
C5389 commonsourceibias.n212 gnd 0.068768f
C5390 commonsourceibias.n213 gnd 0.009225f
C5391 commonsourceibias.t103 gnd 0.17235f
C5392 commonsourceibias.n214 gnd 0.068768f
C5393 commonsourceibias.n215 gnd 0.009225f
C5394 commonsourceibias.t48 gnd 0.17235f
C5395 commonsourceibias.n216 gnd 0.068768f
C5396 commonsourceibias.n217 gnd 0.046441f
C5397 commonsourceibias.t102 gnd 0.17235f
C5398 commonsourceibias.t98 gnd 0.194477f
C5399 commonsourceibias.n218 gnd 0.079804f
C5400 commonsourceibias.n219 gnd 0.082619f
C5401 commonsourceibias.n220 gnd 0.01137f
C5402 commonsourceibias.n221 gnd 0.012578f
C5403 commonsourceibias.n222 gnd 0.009225f
C5404 commonsourceibias.n223 gnd 0.009225f
C5405 commonsourceibias.n224 gnd 0.012496f
C5406 commonsourceibias.n225 gnd 0.007462f
C5407 commonsourceibias.n226 gnd 0.012651f
C5408 commonsourceibias.n227 gnd 0.009225f
C5409 commonsourceibias.n228 gnd 0.009225f
C5410 commonsourceibias.n229 gnd 0.012728f
C5411 commonsourceibias.n230 gnd 0.010975f
C5412 commonsourceibias.n231 gnd 0.008906f
C5413 commonsourceibias.n232 gnd 0.009225f
C5414 commonsourceibias.n233 gnd 0.009225f
C5415 commonsourceibias.n234 gnd 0.011283f
C5416 commonsourceibias.n235 gnd 0.012665f
C5417 commonsourceibias.n236 gnd 0.068768f
C5418 commonsourceibias.n237 gnd 0.01258f
C5419 commonsourceibias.n238 gnd 0.009225f
C5420 commonsourceibias.n239 gnd 0.009225f
C5421 commonsourceibias.n240 gnd 0.009225f
C5422 commonsourceibias.n241 gnd 0.01258f
C5423 commonsourceibias.n242 gnd 0.068768f
C5424 commonsourceibias.n243 gnd 0.012665f
C5425 commonsourceibias.n244 gnd 0.011283f
C5426 commonsourceibias.n245 gnd 0.009225f
C5427 commonsourceibias.n246 gnd 0.009225f
C5428 commonsourceibias.n247 gnd 0.009225f
C5429 commonsourceibias.n248 gnd 0.010975f
C5430 commonsourceibias.n249 gnd 0.012728f
C5431 commonsourceibias.n250 gnd 0.068768f
C5432 commonsourceibias.n251 gnd 0.012651f
C5433 commonsourceibias.n252 gnd 0.009225f
C5434 commonsourceibias.n253 gnd 0.009225f
C5435 commonsourceibias.n254 gnd 0.009225f
C5436 commonsourceibias.n255 gnd 0.012496f
C5437 commonsourceibias.n256 gnd 0.068768f
C5438 commonsourceibias.n257 gnd 0.012578f
C5439 commonsourceibias.n258 gnd 0.01137f
C5440 commonsourceibias.n259 gnd 0.009225f
C5441 commonsourceibias.n260 gnd 0.009225f
C5442 commonsourceibias.n261 gnd 0.009358f
C5443 commonsourceibias.n262 gnd 0.009674f
C5444 commonsourceibias.t109 gnd 0.186396f
C5445 commonsourceibias.n263 gnd 0.082281f
C5446 commonsourceibias.n264 gnd 0.028001f
C5447 commonsourceibias.n265 gnd 0.438243f
C5448 commonsourceibias.n266 gnd 0.01231f
C5449 commonsourceibias.t69 gnd 0.186396f
C5450 commonsourceibias.t99 gnd 0.17235f
C5451 commonsourceibias.n267 gnd 0.068768f
C5452 commonsourceibias.n268 gnd 0.009225f
C5453 commonsourceibias.t84 gnd 0.17235f
C5454 commonsourceibias.n269 gnd 0.007462f
C5455 commonsourceibias.n270 gnd 0.009225f
C5456 commonsourceibias.t72 gnd 0.17235f
C5457 commonsourceibias.n271 gnd 0.008906f
C5458 commonsourceibias.n272 gnd 0.009225f
C5459 commonsourceibias.t66 gnd 0.17235f
C5460 commonsourceibias.n273 gnd 0.007451f
C5461 commonsourceibias.n274 gnd 0.009225f
C5462 commonsourceibias.t56 gnd 0.17235f
C5463 commonsourceibias.t79 gnd 0.17235f
C5464 commonsourceibias.n275 gnd 0.068768f
C5465 commonsourceibias.n276 gnd 0.009225f
C5466 commonsourceibias.t67 gnd 0.17235f
C5467 commonsourceibias.n277 gnd 0.068768f
C5468 commonsourceibias.n278 gnd 0.009225f
C5469 commonsourceibias.t104 gnd 0.17235f
C5470 commonsourceibias.n279 gnd 0.068768f
C5471 commonsourceibias.n280 gnd 0.046441f
C5472 commonsourceibias.t64 gnd 0.17235f
C5473 commonsourceibias.t111 gnd 0.194477f
C5474 commonsourceibias.n281 gnd 0.079804f
C5475 commonsourceibias.n282 gnd 0.082619f
C5476 commonsourceibias.n283 gnd 0.01137f
C5477 commonsourceibias.n284 gnd 0.012578f
C5478 commonsourceibias.n285 gnd 0.009225f
C5479 commonsourceibias.n286 gnd 0.009225f
C5480 commonsourceibias.n287 gnd 0.012496f
C5481 commonsourceibias.n288 gnd 0.007462f
C5482 commonsourceibias.n289 gnd 0.012651f
C5483 commonsourceibias.n290 gnd 0.009225f
C5484 commonsourceibias.n291 gnd 0.009225f
C5485 commonsourceibias.n292 gnd 0.012728f
C5486 commonsourceibias.n293 gnd 0.010975f
C5487 commonsourceibias.n294 gnd 0.008906f
C5488 commonsourceibias.n295 gnd 0.009225f
C5489 commonsourceibias.n296 gnd 0.009225f
C5490 commonsourceibias.n297 gnd 0.011283f
C5491 commonsourceibias.n298 gnd 0.012665f
C5492 commonsourceibias.n299 gnd 0.068768f
C5493 commonsourceibias.n300 gnd 0.01258f
C5494 commonsourceibias.n301 gnd 0.009181f
C5495 commonsourceibias.t41 gnd 0.019906f
C5496 commonsourceibias.t33 gnd 0.019906f
C5497 commonsourceibias.n302 gnd 0.176489f
C5498 commonsourceibias.t43 gnd 0.019906f
C5499 commonsourceibias.t29 gnd 0.019906f
C5500 commonsourceibias.n303 gnd 0.1759f
C5501 commonsourceibias.n304 gnd 0.163906f
C5502 commonsourceibias.t19 gnd 0.019906f
C5503 commonsourceibias.t37 gnd 0.019906f
C5504 commonsourceibias.n305 gnd 0.1759f
C5505 commonsourceibias.n306 gnd 0.067503f
C5506 commonsourceibias.n307 gnd 0.01231f
C5507 commonsourceibias.t46 gnd 0.17235f
C5508 commonsourceibias.n308 gnd 0.068768f
C5509 commonsourceibias.n309 gnd 0.009225f
C5510 commonsourceibias.t14 gnd 0.17235f
C5511 commonsourceibias.n310 gnd 0.007462f
C5512 commonsourceibias.n311 gnd 0.009225f
C5513 commonsourceibias.t24 gnd 0.17235f
C5514 commonsourceibias.n312 gnd 0.008906f
C5515 commonsourceibias.n313 gnd 0.009225f
C5516 commonsourceibias.t30 gnd 0.17235f
C5517 commonsourceibias.n314 gnd 0.007451f
C5518 commonsourceibias.n315 gnd 0.009225f
C5519 commonsourceibias.t36 gnd 0.17235f
C5520 commonsourceibias.t18 gnd 0.17235f
C5521 commonsourceibias.n316 gnd 0.068768f
C5522 commonsourceibias.n317 gnd 0.009225f
C5523 commonsourceibias.t28 gnd 0.17235f
C5524 commonsourceibias.n318 gnd 0.068768f
C5525 commonsourceibias.n319 gnd 0.009225f
C5526 commonsourceibias.t42 gnd 0.17235f
C5527 commonsourceibias.n320 gnd 0.068768f
C5528 commonsourceibias.n321 gnd 0.046441f
C5529 commonsourceibias.t32 gnd 0.17235f
C5530 commonsourceibias.t40 gnd 0.194477f
C5531 commonsourceibias.n322 gnd 0.079804f
C5532 commonsourceibias.n323 gnd 0.082619f
C5533 commonsourceibias.n324 gnd 0.01137f
C5534 commonsourceibias.n325 gnd 0.012578f
C5535 commonsourceibias.n326 gnd 0.009225f
C5536 commonsourceibias.n327 gnd 0.009225f
C5537 commonsourceibias.n328 gnd 0.012496f
C5538 commonsourceibias.n329 gnd 0.007462f
C5539 commonsourceibias.n330 gnd 0.012651f
C5540 commonsourceibias.n331 gnd 0.009225f
C5541 commonsourceibias.n332 gnd 0.009225f
C5542 commonsourceibias.n333 gnd 0.012728f
C5543 commonsourceibias.n334 gnd 0.010975f
C5544 commonsourceibias.n335 gnd 0.008906f
C5545 commonsourceibias.n336 gnd 0.009225f
C5546 commonsourceibias.n337 gnd 0.009225f
C5547 commonsourceibias.n338 gnd 0.011283f
C5548 commonsourceibias.n339 gnd 0.012665f
C5549 commonsourceibias.n340 gnd 0.068768f
C5550 commonsourceibias.n341 gnd 0.01258f
C5551 commonsourceibias.n342 gnd 0.009225f
C5552 commonsourceibias.n343 gnd 0.009225f
C5553 commonsourceibias.n344 gnd 0.009225f
C5554 commonsourceibias.n345 gnd 0.01258f
C5555 commonsourceibias.n346 gnd 0.068768f
C5556 commonsourceibias.n347 gnd 0.012665f
C5557 commonsourceibias.t4 gnd 0.17235f
C5558 commonsourceibias.n348 gnd 0.068768f
C5559 commonsourceibias.n349 gnd 0.011283f
C5560 commonsourceibias.n350 gnd 0.009225f
C5561 commonsourceibias.n351 gnd 0.009225f
C5562 commonsourceibias.n352 gnd 0.009225f
C5563 commonsourceibias.n353 gnd 0.010975f
C5564 commonsourceibias.n354 gnd 0.012728f
C5565 commonsourceibias.n355 gnd 0.068768f
C5566 commonsourceibias.n356 gnd 0.012651f
C5567 commonsourceibias.n357 gnd 0.009225f
C5568 commonsourceibias.n358 gnd 0.009225f
C5569 commonsourceibias.n359 gnd 0.009225f
C5570 commonsourceibias.n360 gnd 0.012496f
C5571 commonsourceibias.n361 gnd 0.068768f
C5572 commonsourceibias.n362 gnd 0.012578f
C5573 commonsourceibias.n363 gnd 0.01137f
C5574 commonsourceibias.n364 gnd 0.009225f
C5575 commonsourceibias.n365 gnd 0.009225f
C5576 commonsourceibias.n366 gnd 0.009358f
C5577 commonsourceibias.n367 gnd 0.009674f
C5578 commonsourceibias.t26 gnd 0.186396f
C5579 commonsourceibias.n368 gnd 0.082281f
C5580 commonsourceibias.n369 gnd 0.091278f
C5581 commonsourceibias.t47 gnd 0.019906f
C5582 commonsourceibias.t27 gnd 0.019906f
C5583 commonsourceibias.n370 gnd 0.1759f
C5584 commonsourceibias.n371 gnd 0.151991f
C5585 commonsourceibias.t25 gnd 0.019906f
C5586 commonsourceibias.t15 gnd 0.019906f
C5587 commonsourceibias.n372 gnd 0.1759f
C5588 commonsourceibias.n373 gnd 0.080798f
C5589 commonsourceibias.t31 gnd 0.019906f
C5590 commonsourceibias.t5 gnd 0.019906f
C5591 commonsourceibias.n374 gnd 0.1759f
C5592 commonsourceibias.n375 gnd 0.067503f
C5593 commonsourceibias.n376 gnd 0.081739f
C5594 commonsourceibias.n377 gnd 0.066685f
C5595 commonsourceibias.n378 gnd 0.009181f
C5596 commonsourceibias.n379 gnd 0.01258f
C5597 commonsourceibias.n380 gnd 0.068768f
C5598 commonsourceibias.n381 gnd 0.012665f
C5599 commonsourceibias.t92 gnd 0.17235f
C5600 commonsourceibias.n382 gnd 0.068768f
C5601 commonsourceibias.n383 gnd 0.011283f
C5602 commonsourceibias.n384 gnd 0.009225f
C5603 commonsourceibias.n385 gnd 0.009225f
C5604 commonsourceibias.n386 gnd 0.009225f
C5605 commonsourceibias.n387 gnd 0.010975f
C5606 commonsourceibias.n388 gnd 0.012728f
C5607 commonsourceibias.n389 gnd 0.068768f
C5608 commonsourceibias.n390 gnd 0.012651f
C5609 commonsourceibias.n391 gnd 0.009225f
C5610 commonsourceibias.n392 gnd 0.009225f
C5611 commonsourceibias.n393 gnd 0.009225f
C5612 commonsourceibias.n394 gnd 0.012496f
C5613 commonsourceibias.n395 gnd 0.068768f
C5614 commonsourceibias.n396 gnd 0.012578f
C5615 commonsourceibias.n397 gnd 0.01137f
C5616 commonsourceibias.n398 gnd 0.009225f
C5617 commonsourceibias.n399 gnd 0.009225f
C5618 commonsourceibias.n400 gnd 0.009358f
C5619 commonsourceibias.n401 gnd 0.009674f
C5620 commonsourceibias.n402 gnd 0.082281f
C5621 commonsourceibias.n403 gnd 0.053268f
C5622 commonsourceibias.n404 gnd 0.01231f
C5623 commonsourceibias.t107 gnd 0.17235f
C5624 commonsourceibias.n405 gnd 0.068768f
C5625 commonsourceibias.n406 gnd 0.009225f
C5626 commonsourceibias.t50 gnd 0.17235f
C5627 commonsourceibias.n407 gnd 0.007462f
C5628 commonsourceibias.n408 gnd 0.009225f
C5629 commonsourceibias.t114 gnd 0.17235f
C5630 commonsourceibias.n409 gnd 0.008906f
C5631 commonsourceibias.n410 gnd 0.009225f
C5632 commonsourceibias.t49 gnd 0.17235f
C5633 commonsourceibias.n411 gnd 0.007451f
C5634 commonsourceibias.n412 gnd 0.009225f
C5635 commonsourceibias.t74 gnd 0.17235f
C5636 commonsourceibias.t105 gnd 0.17235f
C5637 commonsourceibias.n413 gnd 0.068768f
C5638 commonsourceibias.n414 gnd 0.009225f
C5639 commonsourceibias.t55 gnd 0.17235f
C5640 commonsourceibias.n415 gnd 0.068768f
C5641 commonsourceibias.n416 gnd 0.009225f
C5642 commonsourceibias.t75 gnd 0.17235f
C5643 commonsourceibias.n417 gnd 0.068768f
C5644 commonsourceibias.n418 gnd 0.046441f
C5645 commonsourceibias.t61 gnd 0.17235f
C5646 commonsourceibias.t52 gnd 0.194477f
C5647 commonsourceibias.n419 gnd 0.079804f
C5648 commonsourceibias.n420 gnd 0.082619f
C5649 commonsourceibias.n421 gnd 0.01137f
C5650 commonsourceibias.n422 gnd 0.012578f
C5651 commonsourceibias.n423 gnd 0.009225f
C5652 commonsourceibias.n424 gnd 0.009225f
C5653 commonsourceibias.n425 gnd 0.012496f
C5654 commonsourceibias.n426 gnd 0.007462f
C5655 commonsourceibias.n427 gnd 0.012651f
C5656 commonsourceibias.n428 gnd 0.009225f
C5657 commonsourceibias.n429 gnd 0.009225f
C5658 commonsourceibias.n430 gnd 0.012728f
C5659 commonsourceibias.n431 gnd 0.010975f
C5660 commonsourceibias.n432 gnd 0.008906f
C5661 commonsourceibias.n433 gnd 0.009225f
C5662 commonsourceibias.n434 gnd 0.009225f
C5663 commonsourceibias.n435 gnd 0.011283f
C5664 commonsourceibias.n436 gnd 0.012665f
C5665 commonsourceibias.n437 gnd 0.068768f
C5666 commonsourceibias.n438 gnd 0.01258f
C5667 commonsourceibias.n439 gnd 0.009225f
C5668 commonsourceibias.n440 gnd 0.009225f
C5669 commonsourceibias.n441 gnd 0.009225f
C5670 commonsourceibias.n442 gnd 0.01258f
C5671 commonsourceibias.n443 gnd 0.068768f
C5672 commonsourceibias.n444 gnd 0.012665f
C5673 commonsourceibias.t106 gnd 0.17235f
C5674 commonsourceibias.n445 gnd 0.068768f
C5675 commonsourceibias.n446 gnd 0.011283f
C5676 commonsourceibias.n447 gnd 0.009225f
C5677 commonsourceibias.n448 gnd 0.009225f
C5678 commonsourceibias.n449 gnd 0.009225f
C5679 commonsourceibias.n450 gnd 0.010975f
C5680 commonsourceibias.n451 gnd 0.012728f
C5681 commonsourceibias.n452 gnd 0.068768f
C5682 commonsourceibias.n453 gnd 0.012651f
C5683 commonsourceibias.n454 gnd 0.009225f
C5684 commonsourceibias.n455 gnd 0.009225f
C5685 commonsourceibias.n456 gnd 0.009225f
C5686 commonsourceibias.n457 gnd 0.012496f
C5687 commonsourceibias.n458 gnd 0.068768f
C5688 commonsourceibias.n459 gnd 0.012578f
C5689 commonsourceibias.n460 gnd 0.01137f
C5690 commonsourceibias.n461 gnd 0.009225f
C5691 commonsourceibias.n462 gnd 0.009225f
C5692 commonsourceibias.n463 gnd 0.009358f
C5693 commonsourceibias.n464 gnd 0.009674f
C5694 commonsourceibias.t112 gnd 0.186396f
C5695 commonsourceibias.n465 gnd 0.082281f
C5696 commonsourceibias.n466 gnd 0.028001f
C5697 commonsourceibias.n467 gnd 0.147196f
C5698 commonsourceibias.n468 gnd 0.01231f
C5699 commonsourceibias.t81 gnd 0.17235f
C5700 commonsourceibias.n469 gnd 0.068768f
C5701 commonsourceibias.n470 gnd 0.009225f
C5702 commonsourceibias.t91 gnd 0.17235f
C5703 commonsourceibias.n471 gnd 0.007462f
C5704 commonsourceibias.n472 gnd 0.009225f
C5705 commonsourceibias.t100 gnd 0.17235f
C5706 commonsourceibias.n473 gnd 0.008906f
C5707 commonsourceibias.n474 gnd 0.009225f
C5708 commonsourceibias.t85 gnd 0.17235f
C5709 commonsourceibias.n475 gnd 0.007451f
C5710 commonsourceibias.n476 gnd 0.009225f
C5711 commonsourceibias.t82 gnd 0.17235f
C5712 commonsourceibias.t62 gnd 0.17235f
C5713 commonsourceibias.n477 gnd 0.068768f
C5714 commonsourceibias.n478 gnd 0.009225f
C5715 commonsourceibias.t53 gnd 0.17235f
C5716 commonsourceibias.n479 gnd 0.068768f
C5717 commonsourceibias.n480 gnd 0.009225f
C5718 commonsourceibias.t78 gnd 0.17235f
C5719 commonsourceibias.n481 gnd 0.068768f
C5720 commonsourceibias.n482 gnd 0.046441f
C5721 commonsourceibias.t97 gnd 0.17235f
C5722 commonsourceibias.t113 gnd 0.194477f
C5723 commonsourceibias.n483 gnd 0.079804f
C5724 commonsourceibias.n484 gnd 0.082619f
C5725 commonsourceibias.n485 gnd 0.01137f
C5726 commonsourceibias.n486 gnd 0.012578f
C5727 commonsourceibias.n487 gnd 0.009225f
C5728 commonsourceibias.n488 gnd 0.009225f
C5729 commonsourceibias.n489 gnd 0.012496f
C5730 commonsourceibias.n490 gnd 0.007462f
C5731 commonsourceibias.n491 gnd 0.012651f
C5732 commonsourceibias.n492 gnd 0.009225f
C5733 commonsourceibias.n493 gnd 0.009225f
C5734 commonsourceibias.n494 gnd 0.012728f
C5735 commonsourceibias.n495 gnd 0.010975f
C5736 commonsourceibias.n496 gnd 0.008906f
C5737 commonsourceibias.n497 gnd 0.009225f
C5738 commonsourceibias.n498 gnd 0.009225f
C5739 commonsourceibias.n499 gnd 0.011283f
C5740 commonsourceibias.n500 gnd 0.012665f
C5741 commonsourceibias.n501 gnd 0.068768f
C5742 commonsourceibias.n502 gnd 0.01258f
C5743 commonsourceibias.n503 gnd 0.009225f
C5744 commonsourceibias.n504 gnd 0.009225f
C5745 commonsourceibias.n505 gnd 0.009225f
C5746 commonsourceibias.n506 gnd 0.01258f
C5747 commonsourceibias.n507 gnd 0.068768f
C5748 commonsourceibias.n508 gnd 0.012665f
C5749 commonsourceibias.t76 gnd 0.17235f
C5750 commonsourceibias.n509 gnd 0.068768f
C5751 commonsourceibias.n510 gnd 0.011283f
C5752 commonsourceibias.n511 gnd 0.009225f
C5753 commonsourceibias.n512 gnd 0.009225f
C5754 commonsourceibias.n513 gnd 0.009225f
C5755 commonsourceibias.n514 gnd 0.010975f
C5756 commonsourceibias.n515 gnd 0.012728f
C5757 commonsourceibias.n516 gnd 0.068768f
C5758 commonsourceibias.n517 gnd 0.012651f
C5759 commonsourceibias.n518 gnd 0.009225f
C5760 commonsourceibias.n519 gnd 0.009225f
C5761 commonsourceibias.n520 gnd 0.009225f
C5762 commonsourceibias.n521 gnd 0.012496f
C5763 commonsourceibias.n522 gnd 0.068768f
C5764 commonsourceibias.n523 gnd 0.012578f
C5765 commonsourceibias.n524 gnd 0.01137f
C5766 commonsourceibias.n525 gnd 0.009225f
C5767 commonsourceibias.n526 gnd 0.009225f
C5768 commonsourceibias.n527 gnd 0.009358f
C5769 commonsourceibias.n528 gnd 0.009674f
C5770 commonsourceibias.t63 gnd 0.186396f
C5771 commonsourceibias.n529 gnd 0.082281f
C5772 commonsourceibias.n530 gnd 0.028001f
C5773 commonsourceibias.n531 gnd 0.194447f
C5774 commonsourceibias.n532 gnd 4.93338f
C5775 a_n9628_8799.t30 gnd 0.112861f
C5776 a_n9628_8799.t13 gnd 0.145107f
C5777 a_n9628_8799.t12 gnd 0.145107f
C5778 a_n9628_8799.n0 gnd 1.14448f
C5779 a_n9628_8799.t38 gnd 0.145107f
C5780 a_n9628_8799.t18 gnd 0.145107f
C5781 a_n9628_8799.n1 gnd 1.14259f
C5782 a_n9628_8799.n2 gnd 1.02705f
C5783 a_n9628_8799.t0 gnd 0.145107f
C5784 a_n9628_8799.t15 gnd 0.145107f
C5785 a_n9628_8799.n3 gnd 1.14259f
C5786 a_n9628_8799.n4 gnd 0.506252f
C5787 a_n9628_8799.t11 gnd 0.145107f
C5788 a_n9628_8799.t14 gnd 0.145107f
C5789 a_n9628_8799.n5 gnd 1.14259f
C5790 a_n9628_8799.n6 gnd 0.506252f
C5791 a_n9628_8799.t8 gnd 0.145107f
C5792 a_n9628_8799.t36 gnd 0.145107f
C5793 a_n9628_8799.n7 gnd 1.14259f
C5794 a_n9628_8799.n8 gnd 0.506252f
C5795 a_n9628_8799.t3 gnd 0.145107f
C5796 a_n9628_8799.t9 gnd 0.145107f
C5797 a_n9628_8799.n9 gnd 1.14259f
C5798 a_n9628_8799.n10 gnd 3.67858f
C5799 a_n9628_8799.t17 gnd 0.145107f
C5800 a_n9628_8799.t39 gnd 0.145107f
C5801 a_n9628_8799.n11 gnd 1.14448f
C5802 a_n9628_8799.t5 gnd 0.145107f
C5803 a_n9628_8799.t4 gnd 0.145107f
C5804 a_n9628_8799.n12 gnd 1.14259f
C5805 a_n9628_8799.n13 gnd 1.02705f
C5806 a_n9628_8799.t2 gnd 0.145107f
C5807 a_n9628_8799.t16 gnd 0.145107f
C5808 a_n9628_8799.n14 gnd 1.14259f
C5809 a_n9628_8799.n15 gnd 0.506252f
C5810 a_n9628_8799.t35 gnd 0.145107f
C5811 a_n9628_8799.t10 gnd 0.145107f
C5812 a_n9628_8799.n16 gnd 1.14259f
C5813 a_n9628_8799.n17 gnd 0.506252f
C5814 a_n9628_8799.t6 gnd 0.145107f
C5815 a_n9628_8799.t37 gnd 0.145107f
C5816 a_n9628_8799.n18 gnd 1.14259f
C5817 a_n9628_8799.n19 gnd 0.506252f
C5818 a_n9628_8799.t7 gnd 0.145107f
C5819 a_n9628_8799.t1 gnd 0.145107f
C5820 a_n9628_8799.n20 gnd 1.14259f
C5821 a_n9628_8799.n21 gnd 2.55397f
C5822 a_n9628_8799.n22 gnd 7.67998f
C5823 a_n9628_8799.n23 gnd 0.052301f
C5824 a_n9628_8799.t86 gnd 0.60168f
C5825 a_n9628_8799.n24 gnd 0.268722f
C5826 a_n9628_8799.n25 gnd 0.052301f
C5827 a_n9628_8799.n26 gnd 0.011868f
C5828 a_n9628_8799.t122 gnd 0.60168f
C5829 a_n9628_8799.n27 gnd 0.052301f
C5830 a_n9628_8799.t143 gnd 0.60168f
C5831 a_n9628_8799.n28 gnd 0.265659f
C5832 a_n9628_8799.t144 gnd 0.60168f
C5833 a_n9628_8799.n29 gnd 0.052301f
C5834 a_n9628_8799.t72 gnd 0.60168f
C5835 a_n9628_8799.n30 gnd 0.265981f
C5836 a_n9628_8799.n31 gnd 0.052301f
C5837 a_n9628_8799.n32 gnd 0.011868f
C5838 a_n9628_8799.t112 gnd 0.60168f
C5839 a_n9628_8799.n33 gnd 0.052301f
C5840 a_n9628_8799.t119 gnd 0.60168f
C5841 a_n9628_8799.n34 gnd 0.268722f
C5842 a_n9628_8799.n35 gnd 0.052301f
C5843 a_n9628_8799.n36 gnd 0.011868f
C5844 a_n9628_8799.t48 gnd 0.60168f
C5845 a_n9628_8799.n37 gnd 0.165234f
C5846 a_n9628_8799.t91 gnd 0.60168f
C5847 a_n9628_8799.t89 gnd 0.613068f
C5848 a_n9628_8799.n38 gnd 0.252229f
C5849 a_n9628_8799.n39 gnd 0.265014f
C5850 a_n9628_8799.n40 gnd 0.011868f
C5851 a_n9628_8799.t123 gnd 0.60168f
C5852 a_n9628_8799.n41 gnd 0.268722f
C5853 a_n9628_8799.n42 gnd 0.052301f
C5854 a_n9628_8799.n43 gnd 0.052301f
C5855 a_n9628_8799.n44 gnd 0.052301f
C5856 a_n9628_8799.n45 gnd 0.266626f
C5857 a_n9628_8799.t87 gnd 0.60168f
C5858 a_n9628_8799.n46 gnd 0.265336f
C5859 a_n9628_8799.n47 gnd 0.011868f
C5860 a_n9628_8799.n48 gnd 0.052301f
C5861 a_n9628_8799.n49 gnd 0.052301f
C5862 a_n9628_8799.n50 gnd 0.052301f
C5863 a_n9628_8799.n51 gnd 0.011868f
C5864 a_n9628_8799.t42 gnd 0.60168f
C5865 a_n9628_8799.n52 gnd 0.266303f
C5866 a_n9628_8799.t74 gnd 0.60168f
C5867 a_n9628_8799.n53 gnd 0.265659f
C5868 a_n9628_8799.n54 gnd 0.052301f
C5869 a_n9628_8799.n55 gnd 0.052301f
C5870 a_n9628_8799.n56 gnd 0.052301f
C5871 a_n9628_8799.n57 gnd 0.268722f
C5872 a_n9628_8799.n58 gnd 0.011868f
C5873 a_n9628_8799.t147 gnd 0.60168f
C5874 a_n9628_8799.n59 gnd 0.265981f
C5875 a_n9628_8799.n60 gnd 0.052301f
C5876 a_n9628_8799.n61 gnd 0.052301f
C5877 a_n9628_8799.n62 gnd 0.052301f
C5878 a_n9628_8799.n63 gnd 0.011868f
C5879 a_n9628_8799.t108 gnd 0.60168f
C5880 a_n9628_8799.n64 gnd 0.268722f
C5881 a_n9628_8799.n65 gnd 0.011868f
C5882 a_n9628_8799.n66 gnd 0.052301f
C5883 a_n9628_8799.n67 gnd 0.052301f
C5884 a_n9628_8799.n68 gnd 0.052301f
C5885 a_n9628_8799.n69 gnd 0.266303f
C5886 a_n9628_8799.n70 gnd 0.011868f
C5887 a_n9628_8799.t90 gnd 0.60168f
C5888 a_n9628_8799.n71 gnd 0.268722f
C5889 a_n9628_8799.n72 gnd 0.052301f
C5890 a_n9628_8799.n73 gnd 0.052301f
C5891 a_n9628_8799.n74 gnd 0.052301f
C5892 a_n9628_8799.n75 gnd 0.265336f
C5893 a_n9628_8799.t142 gnd 0.60168f
C5894 a_n9628_8799.n76 gnd 0.266626f
C5895 a_n9628_8799.n77 gnd 0.011868f
C5896 a_n9628_8799.n78 gnd 0.052301f
C5897 a_n9628_8799.n79 gnd 0.052301f
C5898 a_n9628_8799.n80 gnd 0.052301f
C5899 a_n9628_8799.n81 gnd 0.011868f
C5900 a_n9628_8799.t88 gnd 0.60168f
C5901 a_n9628_8799.n82 gnd 0.265014f
C5902 a_n9628_8799.t120 gnd 0.60168f
C5903 a_n9628_8799.n83 gnd 0.26324f
C5904 a_n9628_8799.n84 gnd 0.296534f
C5905 a_n9628_8799.n85 gnd 0.052301f
C5906 a_n9628_8799.t97 gnd 0.60168f
C5907 a_n9628_8799.n86 gnd 0.268722f
C5908 a_n9628_8799.n87 gnd 0.052301f
C5909 a_n9628_8799.n88 gnd 0.011868f
C5910 a_n9628_8799.t136 gnd 0.60168f
C5911 a_n9628_8799.n89 gnd 0.052301f
C5912 a_n9628_8799.t155 gnd 0.60168f
C5913 a_n9628_8799.n90 gnd 0.265659f
C5914 a_n9628_8799.t157 gnd 0.60168f
C5915 a_n9628_8799.n91 gnd 0.052301f
C5916 a_n9628_8799.t81 gnd 0.60168f
C5917 a_n9628_8799.n92 gnd 0.265981f
C5918 a_n9628_8799.n93 gnd 0.052301f
C5919 a_n9628_8799.n94 gnd 0.011868f
C5920 a_n9628_8799.t125 gnd 0.60168f
C5921 a_n9628_8799.n95 gnd 0.052301f
C5922 a_n9628_8799.t132 gnd 0.60168f
C5923 a_n9628_8799.n96 gnd 0.268722f
C5924 a_n9628_8799.n97 gnd 0.052301f
C5925 a_n9628_8799.n98 gnd 0.011868f
C5926 a_n9628_8799.t60 gnd 0.60168f
C5927 a_n9628_8799.n99 gnd 0.165234f
C5928 a_n9628_8799.t104 gnd 0.60168f
C5929 a_n9628_8799.t102 gnd 0.613068f
C5930 a_n9628_8799.n100 gnd 0.252229f
C5931 a_n9628_8799.n101 gnd 0.265014f
C5932 a_n9628_8799.n102 gnd 0.011868f
C5933 a_n9628_8799.t140 gnd 0.60168f
C5934 a_n9628_8799.n103 gnd 0.268722f
C5935 a_n9628_8799.n104 gnd 0.052301f
C5936 a_n9628_8799.n105 gnd 0.052301f
C5937 a_n9628_8799.n106 gnd 0.052301f
C5938 a_n9628_8799.n107 gnd 0.266626f
C5939 a_n9628_8799.t98 gnd 0.60168f
C5940 a_n9628_8799.n108 gnd 0.265336f
C5941 a_n9628_8799.n109 gnd 0.011868f
C5942 a_n9628_8799.n110 gnd 0.052301f
C5943 a_n9628_8799.n111 gnd 0.052301f
C5944 a_n9628_8799.n112 gnd 0.052301f
C5945 a_n9628_8799.n113 gnd 0.011868f
C5946 a_n9628_8799.t56 gnd 0.60168f
C5947 a_n9628_8799.n114 gnd 0.266303f
C5948 a_n9628_8799.t84 gnd 0.60168f
C5949 a_n9628_8799.n115 gnd 0.265659f
C5950 a_n9628_8799.n116 gnd 0.052301f
C5951 a_n9628_8799.n117 gnd 0.052301f
C5952 a_n9628_8799.n118 gnd 0.052301f
C5953 a_n9628_8799.n119 gnd 0.268722f
C5954 a_n9628_8799.n120 gnd 0.011868f
C5955 a_n9628_8799.t159 gnd 0.60168f
C5956 a_n9628_8799.n121 gnd 0.265981f
C5957 a_n9628_8799.n122 gnd 0.052301f
C5958 a_n9628_8799.n123 gnd 0.052301f
C5959 a_n9628_8799.n124 gnd 0.052301f
C5960 a_n9628_8799.n125 gnd 0.011868f
C5961 a_n9628_8799.t121 gnd 0.60168f
C5962 a_n9628_8799.n126 gnd 0.268722f
C5963 a_n9628_8799.n127 gnd 0.011868f
C5964 a_n9628_8799.n128 gnd 0.052301f
C5965 a_n9628_8799.n129 gnd 0.052301f
C5966 a_n9628_8799.n130 gnd 0.052301f
C5967 a_n9628_8799.n131 gnd 0.266303f
C5968 a_n9628_8799.n132 gnd 0.011868f
C5969 a_n9628_8799.t103 gnd 0.60168f
C5970 a_n9628_8799.n133 gnd 0.268722f
C5971 a_n9628_8799.n134 gnd 0.052301f
C5972 a_n9628_8799.n135 gnd 0.052301f
C5973 a_n9628_8799.n136 gnd 0.052301f
C5974 a_n9628_8799.n137 gnd 0.265336f
C5975 a_n9628_8799.t154 gnd 0.60168f
C5976 a_n9628_8799.n138 gnd 0.266626f
C5977 a_n9628_8799.n139 gnd 0.011868f
C5978 a_n9628_8799.n140 gnd 0.052301f
C5979 a_n9628_8799.n141 gnd 0.052301f
C5980 a_n9628_8799.n142 gnd 0.052301f
C5981 a_n9628_8799.n143 gnd 0.011868f
C5982 a_n9628_8799.t99 gnd 0.60168f
C5983 a_n9628_8799.n144 gnd 0.265014f
C5984 a_n9628_8799.t133 gnd 0.60168f
C5985 a_n9628_8799.n145 gnd 0.26324f
C5986 a_n9628_8799.n146 gnd 0.130362f
C5987 a_n9628_8799.n147 gnd 0.904543f
C5988 a_n9628_8799.n148 gnd 0.052301f
C5989 a_n9628_8799.t63 gnd 0.60168f
C5990 a_n9628_8799.n149 gnd 0.268722f
C5991 a_n9628_8799.n150 gnd 0.052301f
C5992 a_n9628_8799.n151 gnd 0.011868f
C5993 a_n9628_8799.t82 gnd 0.60168f
C5994 a_n9628_8799.n152 gnd 0.052301f
C5995 a_n9628_8799.t116 gnd 0.60168f
C5996 a_n9628_8799.n153 gnd 0.265659f
C5997 a_n9628_8799.t96 gnd 0.60168f
C5998 a_n9628_8799.n154 gnd 0.052301f
C5999 a_n9628_8799.t100 gnd 0.60168f
C6000 a_n9628_8799.n155 gnd 0.265981f
C6001 a_n9628_8799.n156 gnd 0.052301f
C6002 a_n9628_8799.n157 gnd 0.011868f
C6003 a_n9628_8799.t127 gnd 0.60168f
C6004 a_n9628_8799.n158 gnd 0.052301f
C6005 a_n9628_8799.t43 gnd 0.60168f
C6006 a_n9628_8799.n159 gnd 0.268722f
C6007 a_n9628_8799.n160 gnd 0.052301f
C6008 a_n9628_8799.n161 gnd 0.011868f
C6009 a_n9628_8799.t69 gnd 0.60168f
C6010 a_n9628_8799.n162 gnd 0.165234f
C6011 a_n9628_8799.t52 gnd 0.60168f
C6012 a_n9628_8799.t73 gnd 0.613068f
C6013 a_n9628_8799.n163 gnd 0.252229f
C6014 a_n9628_8799.n164 gnd 0.265014f
C6015 a_n9628_8799.n165 gnd 0.011868f
C6016 a_n9628_8799.t114 gnd 0.60168f
C6017 a_n9628_8799.n166 gnd 0.268722f
C6018 a_n9628_8799.n167 gnd 0.052301f
C6019 a_n9628_8799.n168 gnd 0.052301f
C6020 a_n9628_8799.n169 gnd 0.052301f
C6021 a_n9628_8799.n170 gnd 0.266626f
C6022 a_n9628_8799.t92 gnd 0.60168f
C6023 a_n9628_8799.n171 gnd 0.265336f
C6024 a_n9628_8799.n172 gnd 0.011868f
C6025 a_n9628_8799.n173 gnd 0.052301f
C6026 a_n9628_8799.n174 gnd 0.052301f
C6027 a_n9628_8799.n175 gnd 0.052301f
C6028 a_n9628_8799.n176 gnd 0.011868f
C6029 a_n9628_8799.t109 gnd 0.60168f
C6030 a_n9628_8799.n177 gnd 0.266303f
C6031 a_n9628_8799.t61 gnd 0.60168f
C6032 a_n9628_8799.n178 gnd 0.265659f
C6033 a_n9628_8799.n179 gnd 0.052301f
C6034 a_n9628_8799.n180 gnd 0.052301f
C6035 a_n9628_8799.n181 gnd 0.052301f
C6036 a_n9628_8799.n182 gnd 0.268722f
C6037 a_n9628_8799.n183 gnd 0.011868f
C6038 a_n9628_8799.t77 gnd 0.60168f
C6039 a_n9628_8799.n184 gnd 0.265981f
C6040 a_n9628_8799.n185 gnd 0.052301f
C6041 a_n9628_8799.n186 gnd 0.052301f
C6042 a_n9628_8799.n187 gnd 0.052301f
C6043 a_n9628_8799.n188 gnd 0.011868f
C6044 a_n9628_8799.t53 gnd 0.60168f
C6045 a_n9628_8799.n189 gnd 0.268722f
C6046 a_n9628_8799.n190 gnd 0.011868f
C6047 a_n9628_8799.n191 gnd 0.052301f
C6048 a_n9628_8799.n192 gnd 0.052301f
C6049 a_n9628_8799.n193 gnd 0.052301f
C6050 a_n9628_8799.n194 gnd 0.266303f
C6051 a_n9628_8799.n195 gnd 0.011868f
C6052 a_n9628_8799.t135 gnd 0.60168f
C6053 a_n9628_8799.n196 gnd 0.268722f
C6054 a_n9628_8799.n197 gnd 0.052301f
C6055 a_n9628_8799.n198 gnd 0.052301f
C6056 a_n9628_8799.n199 gnd 0.052301f
C6057 a_n9628_8799.n200 gnd 0.265336f
C6058 a_n9628_8799.t145 gnd 0.60168f
C6059 a_n9628_8799.n201 gnd 0.266626f
C6060 a_n9628_8799.n202 gnd 0.011868f
C6061 a_n9628_8799.n203 gnd 0.052301f
C6062 a_n9628_8799.n204 gnd 0.052301f
C6063 a_n9628_8799.n205 gnd 0.052301f
C6064 a_n9628_8799.n206 gnd 0.011868f
C6065 a_n9628_8799.t40 gnd 0.60168f
C6066 a_n9628_8799.n207 gnd 0.265014f
C6067 a_n9628_8799.t105 gnd 0.60168f
C6068 a_n9628_8799.n208 gnd 0.26324f
C6069 a_n9628_8799.n209 gnd 0.130362f
C6070 a_n9628_8799.n210 gnd 1.82001f
C6071 a_n9628_8799.n211 gnd 0.052301f
C6072 a_n9628_8799.t47 gnd 0.60168f
C6073 a_n9628_8799.t45 gnd 0.60168f
C6074 a_n9628_8799.t131 gnd 0.60168f
C6075 a_n9628_8799.n212 gnd 0.268722f
C6076 a_n9628_8799.n213 gnd 0.052301f
C6077 a_n9628_8799.t67 gnd 0.60168f
C6078 a_n9628_8799.t50 gnd 0.60168f
C6079 a_n9628_8799.n214 gnd 0.052301f
C6080 a_n9628_8799.t138 gnd 0.60168f
C6081 a_n9628_8799.n215 gnd 0.268722f
C6082 a_n9628_8799.n216 gnd 0.052301f
C6083 a_n9628_8799.t93 gnd 0.60168f
C6084 a_n9628_8799.t68 gnd 0.60168f
C6085 a_n9628_8799.n217 gnd 0.052301f
C6086 a_n9628_8799.t156 gnd 0.60168f
C6087 a_n9628_8799.n218 gnd 0.268722f
C6088 a_n9628_8799.n219 gnd 0.052301f
C6089 a_n9628_8799.t111 gnd 0.60168f
C6090 a_n9628_8799.t71 gnd 0.60168f
C6091 a_n9628_8799.n220 gnd 0.052301f
C6092 a_n9628_8799.t150 gnd 0.60168f
C6093 a_n9628_8799.n221 gnd 0.268722f
C6094 a_n9628_8799.n222 gnd 0.052301f
C6095 a_n9628_8799.t113 gnd 0.60168f
C6096 a_n9628_8799.t85 gnd 0.60168f
C6097 a_n9628_8799.n223 gnd 0.052301f
C6098 a_n9628_8799.t46 gnd 0.60168f
C6099 a_n9628_8799.n224 gnd 0.268722f
C6100 a_n9628_8799.n225 gnd 0.052301f
C6101 a_n9628_8799.t134 gnd 0.60168f
C6102 a_n9628_8799.t115 gnd 0.60168f
C6103 a_n9628_8799.n226 gnd 0.052301f
C6104 a_n9628_8799.t51 gnd 0.60168f
C6105 a_n9628_8799.n227 gnd 0.268722f
C6106 a_n9628_8799.t137 gnd 0.613068f
C6107 a_n9628_8799.n228 gnd 0.252229f
C6108 a_n9628_8799.t141 gnd 0.60168f
C6109 a_n9628_8799.n229 gnd 0.265014f
C6110 a_n9628_8799.n230 gnd 0.011868f
C6111 a_n9628_8799.n231 gnd 0.165234f
C6112 a_n9628_8799.n232 gnd 0.052301f
C6113 a_n9628_8799.n233 gnd 0.052301f
C6114 a_n9628_8799.n234 gnd 0.011868f
C6115 a_n9628_8799.n235 gnd 0.266626f
C6116 a_n9628_8799.n236 gnd 0.265336f
C6117 a_n9628_8799.n237 gnd 0.011868f
C6118 a_n9628_8799.n238 gnd 0.052301f
C6119 a_n9628_8799.n239 gnd 0.052301f
C6120 a_n9628_8799.n240 gnd 0.052301f
C6121 a_n9628_8799.n241 gnd 0.011868f
C6122 a_n9628_8799.n242 gnd 0.266303f
C6123 a_n9628_8799.n243 gnd 0.265659f
C6124 a_n9628_8799.n244 gnd 0.011868f
C6125 a_n9628_8799.n245 gnd 0.052301f
C6126 a_n9628_8799.n246 gnd 0.052301f
C6127 a_n9628_8799.n247 gnd 0.052301f
C6128 a_n9628_8799.n248 gnd 0.011868f
C6129 a_n9628_8799.n249 gnd 0.265981f
C6130 a_n9628_8799.n250 gnd 0.265981f
C6131 a_n9628_8799.n251 gnd 0.011868f
C6132 a_n9628_8799.n252 gnd 0.052301f
C6133 a_n9628_8799.n253 gnd 0.052301f
C6134 a_n9628_8799.n254 gnd 0.052301f
C6135 a_n9628_8799.n255 gnd 0.011868f
C6136 a_n9628_8799.n256 gnd 0.265659f
C6137 a_n9628_8799.n257 gnd 0.266303f
C6138 a_n9628_8799.n258 gnd 0.011868f
C6139 a_n9628_8799.n259 gnd 0.052301f
C6140 a_n9628_8799.n260 gnd 0.052301f
C6141 a_n9628_8799.n261 gnd 0.052301f
C6142 a_n9628_8799.n262 gnd 0.011868f
C6143 a_n9628_8799.n263 gnd 0.265336f
C6144 a_n9628_8799.n264 gnd 0.266626f
C6145 a_n9628_8799.n265 gnd 0.011868f
C6146 a_n9628_8799.n266 gnd 0.052301f
C6147 a_n9628_8799.n267 gnd 0.052301f
C6148 a_n9628_8799.n268 gnd 0.052301f
C6149 a_n9628_8799.n269 gnd 0.011868f
C6150 a_n9628_8799.n270 gnd 0.265014f
C6151 a_n9628_8799.n271 gnd 0.26324f
C6152 a_n9628_8799.n272 gnd 0.296534f
C6153 a_n9628_8799.n273 gnd 0.052301f
C6154 a_n9628_8799.t58 gnd 0.60168f
C6155 a_n9628_8799.t57 gnd 0.60168f
C6156 a_n9628_8799.t148 gnd 0.60168f
C6157 a_n9628_8799.n274 gnd 0.268722f
C6158 a_n9628_8799.n275 gnd 0.052301f
C6159 a_n9628_8799.t76 gnd 0.60168f
C6160 a_n9628_8799.t65 gnd 0.60168f
C6161 a_n9628_8799.n276 gnd 0.052301f
C6162 a_n9628_8799.t151 gnd 0.60168f
C6163 a_n9628_8799.n277 gnd 0.268722f
C6164 a_n9628_8799.n278 gnd 0.052301f
C6165 a_n9628_8799.t107 gnd 0.60168f
C6166 a_n9628_8799.t79 gnd 0.60168f
C6167 a_n9628_8799.n279 gnd 0.052301f
C6168 a_n9628_8799.t49 gnd 0.60168f
C6169 a_n9628_8799.n280 gnd 0.268722f
C6170 a_n9628_8799.n281 gnd 0.052301f
C6171 a_n9628_8799.t124 gnd 0.60168f
C6172 a_n9628_8799.t80 gnd 0.60168f
C6173 a_n9628_8799.n282 gnd 0.052301f
C6174 a_n9628_8799.t41 gnd 0.60168f
C6175 a_n9628_8799.n283 gnd 0.268722f
C6176 a_n9628_8799.n284 gnd 0.052301f
C6177 a_n9628_8799.t129 gnd 0.60168f
C6178 a_n9628_8799.t95 gnd 0.60168f
C6179 a_n9628_8799.n285 gnd 0.052301f
C6180 a_n9628_8799.t59 gnd 0.60168f
C6181 a_n9628_8799.n286 gnd 0.268722f
C6182 a_n9628_8799.n287 gnd 0.052301f
C6183 a_n9628_8799.t149 gnd 0.60168f
C6184 a_n9628_8799.t130 gnd 0.60168f
C6185 a_n9628_8799.n288 gnd 0.052301f
C6186 a_n9628_8799.t66 gnd 0.60168f
C6187 a_n9628_8799.n289 gnd 0.268722f
C6188 a_n9628_8799.t152 gnd 0.613068f
C6189 a_n9628_8799.n290 gnd 0.252229f
C6190 a_n9628_8799.t153 gnd 0.60168f
C6191 a_n9628_8799.n291 gnd 0.265014f
C6192 a_n9628_8799.n292 gnd 0.011868f
C6193 a_n9628_8799.n293 gnd 0.165234f
C6194 a_n9628_8799.n294 gnd 0.052301f
C6195 a_n9628_8799.n295 gnd 0.052301f
C6196 a_n9628_8799.n296 gnd 0.011868f
C6197 a_n9628_8799.n297 gnd 0.266626f
C6198 a_n9628_8799.n298 gnd 0.265336f
C6199 a_n9628_8799.n299 gnd 0.011868f
C6200 a_n9628_8799.n300 gnd 0.052301f
C6201 a_n9628_8799.n301 gnd 0.052301f
C6202 a_n9628_8799.n302 gnd 0.052301f
C6203 a_n9628_8799.n303 gnd 0.011868f
C6204 a_n9628_8799.n304 gnd 0.266303f
C6205 a_n9628_8799.n305 gnd 0.265659f
C6206 a_n9628_8799.n306 gnd 0.011868f
C6207 a_n9628_8799.n307 gnd 0.052301f
C6208 a_n9628_8799.n308 gnd 0.052301f
C6209 a_n9628_8799.n309 gnd 0.052301f
C6210 a_n9628_8799.n310 gnd 0.011868f
C6211 a_n9628_8799.n311 gnd 0.265981f
C6212 a_n9628_8799.n312 gnd 0.265981f
C6213 a_n9628_8799.n313 gnd 0.011868f
C6214 a_n9628_8799.n314 gnd 0.052301f
C6215 a_n9628_8799.n315 gnd 0.052301f
C6216 a_n9628_8799.n316 gnd 0.052301f
C6217 a_n9628_8799.n317 gnd 0.011868f
C6218 a_n9628_8799.n318 gnd 0.265659f
C6219 a_n9628_8799.n319 gnd 0.266303f
C6220 a_n9628_8799.n320 gnd 0.011868f
C6221 a_n9628_8799.n321 gnd 0.052301f
C6222 a_n9628_8799.n322 gnd 0.052301f
C6223 a_n9628_8799.n323 gnd 0.052301f
C6224 a_n9628_8799.n324 gnd 0.011868f
C6225 a_n9628_8799.n325 gnd 0.265336f
C6226 a_n9628_8799.n326 gnd 0.266626f
C6227 a_n9628_8799.n327 gnd 0.011868f
C6228 a_n9628_8799.n328 gnd 0.052301f
C6229 a_n9628_8799.n329 gnd 0.052301f
C6230 a_n9628_8799.n330 gnd 0.052301f
C6231 a_n9628_8799.n331 gnd 0.011868f
C6232 a_n9628_8799.n332 gnd 0.265014f
C6233 a_n9628_8799.n333 gnd 0.26324f
C6234 a_n9628_8799.n334 gnd 0.130362f
C6235 a_n9628_8799.n335 gnd 0.904543f
C6236 a_n9628_8799.n336 gnd 0.052301f
C6237 a_n9628_8799.t106 gnd 0.60168f
C6238 a_n9628_8799.t128 gnd 0.60168f
C6239 a_n9628_8799.t64 gnd 0.60168f
C6240 a_n9628_8799.n337 gnd 0.268722f
C6241 a_n9628_8799.n338 gnd 0.052301f
C6242 a_n9628_8799.t146 gnd 0.60168f
C6243 a_n9628_8799.t83 gnd 0.60168f
C6244 a_n9628_8799.n339 gnd 0.052301f
C6245 a_n9628_8799.t139 gnd 0.60168f
C6246 a_n9628_8799.n340 gnd 0.268722f
C6247 a_n9628_8799.n341 gnd 0.052301f
C6248 a_n9628_8799.t70 gnd 0.60168f
C6249 a_n9628_8799.t118 gnd 0.60168f
C6250 a_n9628_8799.n342 gnd 0.052301f
C6251 a_n9628_8799.t55 gnd 0.60168f
C6252 a_n9628_8799.n343 gnd 0.268722f
C6253 a_n9628_8799.n344 gnd 0.052301f
C6254 a_n9628_8799.t101 gnd 0.60168f
C6255 a_n9628_8799.t78 gnd 0.60168f
C6256 a_n9628_8799.n345 gnd 0.052301f
C6257 a_n9628_8799.t126 gnd 0.60168f
C6258 a_n9628_8799.n346 gnd 0.268722f
C6259 a_n9628_8799.n347 gnd 0.052301f
C6260 a_n9628_8799.t62 gnd 0.60168f
C6261 a_n9628_8799.t110 gnd 0.60168f
C6262 a_n9628_8799.n348 gnd 0.052301f
C6263 a_n9628_8799.t44 gnd 0.60168f
C6264 a_n9628_8799.n349 gnd 0.268722f
C6265 a_n9628_8799.n350 gnd 0.052301f
C6266 a_n9628_8799.t94 gnd 0.60168f
C6267 a_n9628_8799.t158 gnd 0.60168f
C6268 a_n9628_8799.n351 gnd 0.052301f
C6269 a_n9628_8799.t117 gnd 0.60168f
C6270 a_n9628_8799.n352 gnd 0.268722f
C6271 a_n9628_8799.t75 gnd 0.613068f
C6272 a_n9628_8799.n353 gnd 0.252229f
C6273 a_n9628_8799.t54 gnd 0.60168f
C6274 a_n9628_8799.n354 gnd 0.265014f
C6275 a_n9628_8799.n355 gnd 0.011868f
C6276 a_n9628_8799.n356 gnd 0.165234f
C6277 a_n9628_8799.n357 gnd 0.052301f
C6278 a_n9628_8799.n358 gnd 0.052301f
C6279 a_n9628_8799.n359 gnd 0.011868f
C6280 a_n9628_8799.n360 gnd 0.266626f
C6281 a_n9628_8799.n361 gnd 0.265336f
C6282 a_n9628_8799.n362 gnd 0.011868f
C6283 a_n9628_8799.n363 gnd 0.052301f
C6284 a_n9628_8799.n364 gnd 0.052301f
C6285 a_n9628_8799.n365 gnd 0.052301f
C6286 a_n9628_8799.n366 gnd 0.011868f
C6287 a_n9628_8799.n367 gnd 0.266303f
C6288 a_n9628_8799.n368 gnd 0.265659f
C6289 a_n9628_8799.n369 gnd 0.011868f
C6290 a_n9628_8799.n370 gnd 0.052301f
C6291 a_n9628_8799.n371 gnd 0.052301f
C6292 a_n9628_8799.n372 gnd 0.052301f
C6293 a_n9628_8799.n373 gnd 0.011868f
C6294 a_n9628_8799.n374 gnd 0.265981f
C6295 a_n9628_8799.n375 gnd 0.265981f
C6296 a_n9628_8799.n376 gnd 0.011868f
C6297 a_n9628_8799.n377 gnd 0.052301f
C6298 a_n9628_8799.n378 gnd 0.052301f
C6299 a_n9628_8799.n379 gnd 0.052301f
C6300 a_n9628_8799.n380 gnd 0.011868f
C6301 a_n9628_8799.n381 gnd 0.265659f
C6302 a_n9628_8799.n382 gnd 0.266303f
C6303 a_n9628_8799.n383 gnd 0.011868f
C6304 a_n9628_8799.n384 gnd 0.052301f
C6305 a_n9628_8799.n385 gnd 0.052301f
C6306 a_n9628_8799.n386 gnd 0.052301f
C6307 a_n9628_8799.n387 gnd 0.011868f
C6308 a_n9628_8799.n388 gnd 0.265336f
C6309 a_n9628_8799.n389 gnd 0.266626f
C6310 a_n9628_8799.n390 gnd 0.011868f
C6311 a_n9628_8799.n391 gnd 0.052301f
C6312 a_n9628_8799.n392 gnd 0.052301f
C6313 a_n9628_8799.n393 gnd 0.052301f
C6314 a_n9628_8799.n394 gnd 0.011868f
C6315 a_n9628_8799.n395 gnd 0.265014f
C6316 a_n9628_8799.n396 gnd 0.26324f
C6317 a_n9628_8799.n397 gnd 0.130362f
C6318 a_n9628_8799.n398 gnd 1.45483f
C6319 a_n9628_8799.n399 gnd 17.495998f
C6320 a_n9628_8799.n400 gnd 4.40343f
C6321 a_n9628_8799.t24 gnd 0.112861f
C6322 a_n9628_8799.t25 gnd 0.112861f
C6323 a_n9628_8799.n401 gnd 0.999496f
C6324 a_n9628_8799.t20 gnd 0.112861f
C6325 a_n9628_8799.t21 gnd 0.112861f
C6326 a_n9628_8799.n402 gnd 0.997278f
C6327 a_n9628_8799.n403 gnd 0.736003f
C6328 a_n9628_8799.n404 gnd 0.473568f
C6329 a_n9628_8799.t19 gnd 0.112861f
C6330 a_n9628_8799.t31 gnd 0.112861f
C6331 a_n9628_8799.n405 gnd 0.997278f
C6332 a_n9628_8799.n406 gnd 0.331705f
C6333 a_n9628_8799.t32 gnd 0.112861f
C6334 a_n9628_8799.t28 gnd 0.112861f
C6335 a_n9628_8799.n407 gnd 0.997278f
C6336 a_n9628_8799.n408 gnd 2.58607f
C6337 a_n9628_8799.t29 gnd 0.112861f
C6338 a_n9628_8799.t27 gnd 0.112861f
C6339 a_n9628_8799.n409 gnd 0.999495f
C6340 a_n9628_8799.t22 gnd 0.112861f
C6341 a_n9628_8799.t26 gnd 0.112861f
C6342 a_n9628_8799.n410 gnd 0.997277f
C6343 a_n9628_8799.n411 gnd 0.736005f
C6344 a_n9628_8799.n412 gnd 2.0023f
C6345 a_n9628_8799.t33 gnd 0.112861f
C6346 a_n9628_8799.t23 gnd 0.112861f
C6347 a_n9628_8799.n413 gnd 0.997277f
C6348 a_n9628_8799.n414 gnd 0.736007f
C6349 a_n9628_8799.n415 gnd 0.999492f
C6350 a_n9628_8799.t34 gnd 0.112861f
C6351 a_n2903_n3924.n0 gnd 1.55666f
C6352 a_n2903_n3924.n1 gnd 1.85226f
C6353 a_n2903_n3924.n2 gnd 1.34545f
C6354 a_n2903_n3924.n3 gnd 1.34544f
C6355 a_n2903_n3924.n4 gnd 0.82212f
C6356 a_n2903_n3924.n5 gnd 1.64424f
C6357 a_n2903_n3924.n6 gnd 2.30935f
C6358 a_n2903_n3924.n7 gnd 1.18081f
C6359 a_n2903_n3924.n8 gnd 0.885216f
C6360 a_n2903_n3924.n9 gnd 1.97724f
C6361 a_n2903_n3924.t4 gnd 0.090392f
C6362 a_n2903_n3924.t10 gnd 0.090392f
C6363 a_n2903_n3924.n10 gnd 0.738246f
C6364 a_n2903_n3924.t23 gnd 0.939457f
C6365 a_n2903_n3924.t21 gnd 0.090392f
C6366 a_n2903_n3924.t33 gnd 0.090392f
C6367 a_n2903_n3924.n11 gnd 0.738247f
C6368 a_n2903_n3924.t26 gnd 0.090392f
C6369 a_n2903_n3924.t27 gnd 0.090392f
C6370 a_n2903_n3924.n12 gnd 0.738247f
C6371 a_n2903_n3924.t34 gnd 0.090392f
C6372 a_n2903_n3924.t24 gnd 0.090392f
C6373 a_n2903_n3924.n13 gnd 0.738247f
C6374 a_n2903_n3924.t29 gnd 0.939461f
C6375 a_n2903_n3924.t3 gnd 0.939461f
C6376 a_n2903_n3924.t17 gnd 0.090392f
C6377 a_n2903_n3924.t18 gnd 0.090392f
C6378 a_n2903_n3924.n14 gnd 0.738247f
C6379 a_n2903_n3924.t36 gnd 0.090392f
C6380 a_n2903_n3924.t5 gnd 0.090392f
C6381 a_n2903_n3924.n15 gnd 0.738247f
C6382 a_n2903_n3924.t15 gnd 0.090392f
C6383 a_n2903_n3924.t16 gnd 0.090392f
C6384 a_n2903_n3924.n16 gnd 0.738247f
C6385 a_n2903_n3924.t7 gnd 0.939461f
C6386 a_n2903_n3924.t6 gnd 0.090392f
C6387 a_n2903_n3924.t11 gnd 0.090392f
C6388 a_n2903_n3924.n17 gnd 0.738246f
C6389 a_n2903_n3924.t2 gnd 0.939457f
C6390 a_n2903_n3924.t25 gnd 0.939457f
C6391 a_n2903_n3924.t30 gnd 0.090392f
C6392 a_n2903_n3924.t19 gnd 0.090392f
C6393 a_n2903_n3924.n18 gnd 0.738246f
C6394 a_n2903_n3924.t28 gnd 0.090392f
C6395 a_n2903_n3924.t20 gnd 0.090392f
C6396 a_n2903_n3924.n19 gnd 0.738246f
C6397 a_n2903_n3924.t31 gnd 0.090392f
C6398 a_n2903_n3924.t32 gnd 0.090392f
C6399 a_n2903_n3924.n20 gnd 0.738246f
C6400 a_n2903_n3924.t22 gnd 0.939457f
C6401 a_n2903_n3924.n21 gnd 0.847907f
C6402 a_n2903_n3924.t35 gnd 1.16892f
C6403 a_n2903_n3924.t8 gnd 1.16726f
C6404 a_n2903_n3924.t9 gnd 1.16726f
C6405 a_n2903_n3924.t13 gnd 1.16726f
C6406 a_n2903_n3924.t38 gnd 1.16726f
C6407 a_n2903_n3924.t12 gnd 1.16726f
C6408 a_n2903_n3924.t37 gnd 1.16726f
C6409 a_n2903_n3924.t39 gnd 1.16889f
C6410 a_n2903_n3924.n22 gnd 0.847907f
C6411 a_n2903_n3924.t1 gnd 0.939457f
C6412 a_n2903_n3924.t14 gnd 0.090392f
C6413 a_n2903_n3924.n23 gnd 0.738243f
C6414 a_n2903_n3924.t0 gnd 0.090392f
C6415 plus.n0 gnd 0.022222f
C6416 plus.t9 gnd 0.314305f
C6417 plus.n1 gnd 0.022222f
C6418 plus.t5 gnd 0.314305f
C6419 plus.t6 gnd 0.314305f
C6420 plus.n2 gnd 0.139624f
C6421 plus.n3 gnd 0.022222f
C6422 plus.t16 gnd 0.314305f
C6423 plus.t17 gnd 0.314305f
C6424 plus.n4 gnd 0.139624f
C6425 plus.n5 gnd 0.022222f
C6426 plus.t13 gnd 0.314305f
C6427 plus.t10 gnd 0.314305f
C6428 plus.n6 gnd 0.142668f
C6429 plus.t12 gnd 0.324898f
C6430 plus.n7 gnd 0.130881f
C6431 plus.n8 gnd 0.094037f
C6432 plus.n9 gnd 0.005043f
C6433 plus.n10 gnd 0.139624f
C6434 plus.n11 gnd 0.005043f
C6435 plus.n12 gnd 0.022222f
C6436 plus.n13 gnd 0.022222f
C6437 plus.n14 gnd 0.022222f
C6438 plus.n15 gnd 0.005043f
C6439 plus.n16 gnd 0.139624f
C6440 plus.n17 gnd 0.005043f
C6441 plus.n18 gnd 0.022222f
C6442 plus.n19 gnd 0.022222f
C6443 plus.n20 gnd 0.022222f
C6444 plus.n21 gnd 0.005043f
C6445 plus.n22 gnd 0.139624f
C6446 plus.n23 gnd 0.005043f
C6447 plus.n24 gnd 0.139008f
C6448 plus.n25 gnd 0.250433f
C6449 plus.n26 gnd 0.022222f
C6450 plus.n27 gnd 0.005043f
C6451 plus.t7 gnd 0.314305f
C6452 plus.n28 gnd 0.022222f
C6453 plus.n29 gnd 0.005043f
C6454 plus.t20 gnd 0.314305f
C6455 plus.n30 gnd 0.022222f
C6456 plus.n31 gnd 0.005043f
C6457 plus.t19 gnd 0.314305f
C6458 plus.t15 gnd 0.324898f
C6459 plus.t14 gnd 0.314305f
C6460 plus.n32 gnd 0.142668f
C6461 plus.n33 gnd 0.130881f
C6462 plus.n34 gnd 0.094037f
C6463 plus.n35 gnd 0.022222f
C6464 plus.n36 gnd 0.139624f
C6465 plus.n37 gnd 0.005043f
C6466 plus.t18 gnd 0.314305f
C6467 plus.n38 gnd 0.139624f
C6468 plus.n39 gnd 0.022222f
C6469 plus.n40 gnd 0.022222f
C6470 plus.n41 gnd 0.022222f
C6471 plus.n42 gnd 0.139624f
C6472 plus.n43 gnd 0.005043f
C6473 plus.t8 gnd 0.314305f
C6474 plus.n44 gnd 0.139624f
C6475 plus.n45 gnd 0.022222f
C6476 plus.n46 gnd 0.022222f
C6477 plus.n47 gnd 0.022222f
C6478 plus.n48 gnd 0.139624f
C6479 plus.n49 gnd 0.005043f
C6480 plus.t11 gnd 0.314305f
C6481 plus.n50 gnd 0.139008f
C6482 plus.n51 gnd 0.636068f
C6483 plus.n52 gnd 0.972007f
C6484 plus.t3 gnd 0.038361f
C6485 plus.t2 gnd 0.00685f
C6486 plus.t0 gnd 0.00685f
C6487 plus.n53 gnd 0.022217f
C6488 plus.n54 gnd 0.17247f
C6489 plus.t4 gnd 0.00685f
C6490 plus.t1 gnd 0.00685f
C6491 plus.n55 gnd 0.022217f
C6492 plus.n56 gnd 0.12946f
C6493 plus.n57 gnd 2.47803f
.ends

