* NGSPICE file created from opamp506.ext - technology: sky130A

.subckt opamp506 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n2140_13878# a_n2318_13878# a_n2318_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n2140_13878# a_n2318_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=253.8 ps=1.42884k w=8 l=0.5
X4 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X5 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 gnd gnd plus gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X8 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=292.92 ps=1.65752k w=7 l=1
X9 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X10 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X12 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 a_n2318_8322# a_n2318_13878# a_n6308_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X15 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X17 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X18 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X19 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X20 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X22 a_n6308_8799# a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X23 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X25 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X26 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X28 a_n6308_8799# a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X29 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X30 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X31 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X32 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X33 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X35 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X36 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X39 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X40 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X42 a_n2140_13878# a_n2318_13878# a_n2318_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X43 a_n2318_13878# a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X44 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X46 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X47 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X49 outputibias outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X50 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X51 a_n6308_8799# a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X52 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 plus gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X54 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X56 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X57 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X58 CSoutput a_n2318_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X59 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X64 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X66 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X68 CSoutput a_n2318_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X69 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X71 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 a_n6308_8799# a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X74 a_n2318_13878# a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X75 a_n2318_13878# a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X76 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X77 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X80 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X81 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X82 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X83 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X84 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X85 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X86 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X89 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X90 a_n2318_8322# a_n2318_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X91 vdd a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X92 a_n2318_13878# a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X93 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X94 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X95 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X96 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X98 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X99 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X100 vdd a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X101 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X102 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X103 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X104 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X105 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X107 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X108 a_n6308_8799# a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X109 a_n2318_8322# a_n2318_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X110 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X111 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X112 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X113 a_n2318_13878# a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X114 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X115 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X116 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X117 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X118 a_n6308_8799# a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X119 a_n2140_13878# a_n2318_13878# a_n2318_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X120 gnd gnd minus gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X121 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X124 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X125 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X126 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X127 a_n2140_13878# a_n2318_13878# a_n2318_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X128 vdd a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X129 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 a_n2318_13878# a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X132 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 gnd gnd minus gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X134 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X135 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X137 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X140 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X141 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X142 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X144 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X147 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X149 a_n2140_13878# a_n2318_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X150 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X152 vdd a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X155 a_n2140_13878# a_n2318_13878# a_n2318_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 output outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X157 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X158 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X159 CSoutput a_n2318_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X160 a_n2318_8322# a_n2318_13878# a_n6308_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X161 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X162 output outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X163 output outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X164 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X166 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X167 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X168 vdd a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X169 plus gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X170 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X171 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X172 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X173 CSoutput a_n2318_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X174 output outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X175 gnd gnd minus gnd sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X176 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X178 a_n2140_13878# a_n2318_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X179 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X181 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X183 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 minus gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X186 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X187 a_n2318_8322# a_n2318_13878# a_n6308_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X188 vdd a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X189 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X191 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X192 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X193 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X195 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X197 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X198 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X200 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X201 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X202 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X203 a_n2140_13878# a_n2318_13878# a_n2318_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X204 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 a_n2318_8322# a_n2318_13878# a_n6308_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X206 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X208 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X214 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X216 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 a_n2318_8322# a_n2318_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X218 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X219 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X220 vdd a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X221 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X223 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X224 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X227 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X230 minus gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X231 a_n6308_8799# a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X232 a_n2318_8322# a_n2318_13878# a_n6308_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X233 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X234 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X236 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X237 a_n2140_13878# a_n2318_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X238 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X239 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X240 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X241 gnd commonsourceibias commonsourceibias gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X242 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X243 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X244 a_n2318_8322# a_n2318_13878# a_n6308_8799# vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X245 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X246 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X248 a_n2140_13878# a_n2318_13878# a_n2318_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X249 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X250 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X251 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X252 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X254 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X256 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X257 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X258 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X259 a_n6308_8799# a_n2318_13878# a_n2318_8322# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X260 a_n2318_13878# a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X261 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X262 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X263 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X265 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 gnd gnd plus gnd sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X267 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X270 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X271 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X272 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X273 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X274 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X275 a_n2318_8322# a_n2318_13878# a_n6308_8799# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 gnd gnd plus gnd sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X277 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X278 CSoutput a_n2318_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X279 diffpairibias diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X280 a_n3827_n3924# plus a_n6308_8799# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X281 vdd a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X282 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X283 a_n6308_8799# plus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X284 CSoutput a_n2318_8322# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X285 outputibias outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X286 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X289 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 a_n3827_n3924# minus a_n2318_13878# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X291 vdd CSoutput output gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X292 CSoutput a_n6308_8799# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 CSoutput commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 outputibias outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X295 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X296 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X297 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 a_n2318_8322# a_n2318_13878# a_n6308_8799# vdd sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X299 a_n2318_13878# minus a_n3827_n3924# gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X300 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 outputibias outputibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X302 output CSoutput vdd gnd sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X303 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X304 a_n2318_8322# a_n2318_13878# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X305 a_n2140_13878# a_n2318_13878# a_n2318_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X306 gnd commonsourceibias CSoutput gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 vdd a_n6308_8799# CSoutput vdd sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 commonsourceibias commonsourceibias gnd gnd sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 a_n2318_13878# a_n2318_13878# a_n2140_13878# vdd sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X310 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X311 a_n3827_n3924# diffpairibias gnd gnd sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
.ends

